
--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/ccs_in_v1.vhd 
--------------------------------------------------------------------------------
-- Catapult Synthesis - Sample I/O Port Library
--
-- Copyright (c) 2003-2017 Mentor Graphics Corp.
--       All Rights Reserved
--
-- This document may be used and distributed without restriction provided that
-- this copyright statement is not removed from the file and that any derivative
-- work contains this copyright notice.
--
-- The design information contained in this file is intended to be an example
-- of the functionality which the end user may study in preparation for creating
-- their own custom interfaces. This design does not necessarily present a 
-- complete implementation of the named protocol or standard.
--
--------------------------------------------------------------------------------

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;

PACKAGE ccs_in_pkg_v1 IS

COMPONENT ccs_in_v1
  GENERIC (
    rscid    : INTEGER;
    width    : INTEGER
  );
  PORT (
    idat   : OUT std_logic_vector(width-1 DOWNTO 0);
    dat    : IN  std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

END ccs_in_pkg_v1;

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all; -- Prevent STARC 2.1.1.2 violation

ENTITY ccs_in_v1 IS
  GENERIC (
    rscid : INTEGER;
    width : INTEGER
  );
  PORT (
    idat  : OUT std_logic_vector(width-1 DOWNTO 0);
    dat   : IN  std_logic_vector(width-1 DOWNTO 0)
  );
END ccs_in_v1;

ARCHITECTURE beh OF ccs_in_v1 IS
BEGIN

  idat <= dat;

END beh;


--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_io_sync_v2.vhd 
--------------------------------------------------------------------------------
-- Catapult Synthesis - Sample I/O Port Library
--
-- Copyright (c) 2003-2017 Mentor Graphics Corp.
--       All Rights Reserved
--
-- This document may be used and distributed without restriction provided that
-- this copyright statement is not removed from the file and that any derivative
-- work contains this copyright notice.
--
-- The design information contained in this file is intended to be an example
-- of the functionality which the end user may study in preparation for creating
-- their own custom interfaces. This design does not necessarily present a 
-- complete implementation of the named protocol or standard.
--
--------------------------------------------------------------------------------

LIBRARY ieee;

USE ieee.std_logic_1164.all;
PACKAGE mgc_io_sync_pkg_v2 IS

COMPONENT mgc_io_sync_v2
  GENERIC (
    valid    : INTEGER RANGE 0 TO 1
  );
  PORT (
    ld       : IN    std_logic;
    lz       : OUT   std_logic
  );
END COMPONENT;

END mgc_io_sync_pkg_v2;

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all; -- Prevent STARC 2.1.1.2 violation

ENTITY mgc_io_sync_v2 IS
  GENERIC (
    valid    : INTEGER RANGE 0 TO 1
  );
  PORT (
    ld       : IN    std_logic;
    lz       : OUT   std_logic
  );
END mgc_io_sync_v2;

ARCHITECTURE beh OF mgc_io_sync_v2 IS
BEGIN

  lz <= ld;

END beh;


--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/src/funcs.vhd 

-- a package of attributes that give verification tools a hint about
-- the function being implemented
PACKAGE attributes IS
  ATTRIBUTE CALYPTO_FUNC : string;
  ATTRIBUTE CALYPTO_DATA_ORDER : string;
end attributes;

-----------------------------------------------------------------------
-- Package that declares synthesizable functions needed for RTL output
-----------------------------------------------------------------------

LIBRARY ieee;

use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;

PACKAGE funcs IS

-----------------------------------------------------------------
-- utility functions
-----------------------------------------------------------------

   FUNCTION TO_STDLOGIC(arg1: BOOLEAN) RETURN STD_LOGIC;
--   FUNCTION TO_STDLOGIC(arg1: STD_ULOGIC_VECTOR(0 DOWNTO 0)) RETURN STD_LOGIC;
   FUNCTION TO_STDLOGIC(arg1: STD_LOGIC_VECTOR(0 DOWNTO 0)) RETURN STD_LOGIC;
   FUNCTION TO_STDLOGIC(arg1: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION TO_STDLOGIC(arg1: SIGNED(0 DOWNTO 0)) RETURN STD_LOGIC;
   FUNCTION TO_STDLOGICVECTOR(arg1: STD_LOGIC) RETURN STD_LOGIC_VECTOR;

   FUNCTION maximum(arg1, arg2 : INTEGER) RETURN INTEGER;
   FUNCTION minimum(arg1, arg2 : INTEGER) RETURN INTEGER;
   FUNCTION ifeqsel(arg1, arg2, seleq, selne : INTEGER) RETURN INTEGER;
   FUNCTION resolve_std_logic_vector(input1: STD_LOGIC_VECTOR; input2 : STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR;
   
-----------------------------------------------------------------
-- logic functions
-----------------------------------------------------------------

   FUNCTION and_s(inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC;
   FUNCTION or_s (inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC;
   FUNCTION xor_s(inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC;

   FUNCTION and_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR;
   FUNCTION or_v (inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR;
   FUNCTION xor_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR;

-----------------------------------------------------------------
-- mux functions
-----------------------------------------------------------------

   FUNCTION mux_s(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC       ) RETURN STD_LOGIC;
   FUNCTION mux_s(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR) RETURN STD_LOGIC;
   FUNCTION mux_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC       ) RETURN STD_LOGIC_VECTOR;
   FUNCTION mux_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR;

-----------------------------------------------------------------
-- latch functions
-----------------------------------------------------------------
   FUNCTION lat_s(dinput: STD_LOGIC       ; clk: STD_LOGIC; doutput: STD_LOGIC       ) RETURN STD_LOGIC;
   FUNCTION lat_v(dinput: STD_LOGIC_VECTOR; clk: STD_LOGIC; doutput: STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR;

-----------------------------------------------------------------
-- tristate functions
-----------------------------------------------------------------
--   FUNCTION tri_s(dinput: STD_LOGIC       ; control: STD_LOGIC) RETURN STD_LOGIC;
--   FUNCTION tri_v(dinput: STD_LOGIC_VECTOR; control: STD_LOGIC) RETURN STD_LOGIC_VECTOR;

-----------------------------------------------------------------
-- compare functions returning STD_LOGIC
-- in contrast to the functions returning boolean
-----------------------------------------------------------------

   FUNCTION "=" (l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION "=" (l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION "/="(l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION "/="(l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION "<="(l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION "<="(l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION "<" (l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION "<" (l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION ">="(l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION ">="(l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION ">" (l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION ">" (l, r: SIGNED  ) RETURN STD_LOGIC;

   -- RETURN 2 bits (left => lt, right => eq)
   FUNCTION cmp (l, r: STD_LOGIC_VECTOR) RETURN STD_LOGIC;

-----------------------------------------------------------------
-- Vectorized Overloaded Arithmetic Operators
-----------------------------------------------------------------

   FUNCTION faccu(arg: UNSIGNED; width: NATURAL) RETURN UNSIGNED;
 
   FUNCTION fabs(arg1: SIGNED  ) RETURN UNSIGNED;

   FUNCTION "/"  (l, r: UNSIGNED) RETURN UNSIGNED;
   FUNCTION "MOD"(l, r: UNSIGNED) RETURN UNSIGNED;
   FUNCTION "REM"(l, r: UNSIGNED) RETURN UNSIGNED;
   FUNCTION "**" (l, r: UNSIGNED) RETURN UNSIGNED;

   FUNCTION "/"  (l, r: SIGNED  ) RETURN SIGNED  ;
   FUNCTION "MOD"(l, r: SIGNED  ) RETURN SIGNED  ;
   FUNCTION "REM"(l, r: SIGNED  ) RETURN SIGNED  ;
   FUNCTION "**" (l, r: SIGNED  ) RETURN SIGNED  ;

-----------------------------------------------------------------
--               S H I F T   F U C T I O N S
-- negative shift shifts the opposite direction
-- *_stdar functions use shift functions from std_logic_arith
-----------------------------------------------------------------

   FUNCTION fshl(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshl(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED;

   FUNCTION fshl(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshr(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshl(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshr(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED  ;

   FUNCTION fshl(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshl(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;

   FUNCTION frot(arg1: STD_LOGIC_VECTOR; arg2: STD_LOGIC_VECTOR; signd2: BOOLEAN; sdir: INTEGER range -1 TO 1) RETURN STD_LOGIC_VECTOR;
   FUNCTION frol(arg1: STD_LOGIC_VECTOR; arg2: UNSIGNED) RETURN STD_LOGIC_VECTOR;
   FUNCTION fror(arg1: STD_LOGIC_VECTOR; arg2: UNSIGNED) RETURN STD_LOGIC_VECTOR;
   FUNCTION frol(arg1: STD_LOGIC_VECTOR; arg2: SIGNED  ) RETURN STD_LOGIC_VECTOR;
   FUNCTION fror(arg1: STD_LOGIC_VECTOR; arg2: SIGNED  ) RETURN STD_LOGIC_VECTOR;

   -----------------------------------------------------------------
   -- *_stdar functions use shift functions from std_logic_arith
   -----------------------------------------------------------------
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED;

   FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshr_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshr_stdar(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED  ;

   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;

-----------------------------------------------------------------
-- indexing functions: LSB always has index 0
-----------------------------------------------------------------

   FUNCTION readindex(vec: STD_LOGIC_VECTOR; index: INTEGER                 ) RETURN STD_LOGIC;
   FUNCTION readslice(vec: STD_LOGIC_VECTOR; index: INTEGER; width: POSITIVE) RETURN STD_LOGIC_VECTOR;

   FUNCTION writeindex(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC       ; index: INTEGER) RETURN STD_LOGIC_VECTOR;
   FUNCTION n_bits(p: NATURAL) RETURN POSITIVE;
   --FUNCTION writeslice(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC_VECTOR; index: INTEGER) RETURN STD_LOGIC_VECTOR;
   FUNCTION writeslice(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC_VECTOR; enable: STD_LOGIC_VECTOR; byte_width: INTEGER;  index: INTEGER) RETURN STD_LOGIC_VECTOR ;

   FUNCTION ceil_log2(size : NATURAL) return NATURAL;
   FUNCTION bits(size : NATURAL) return NATURAL;    

   PROCEDURE csa(a, b, c: IN INTEGER; s, cout: OUT STD_LOGIC_VECTOR);
   PROCEDURE csha(a, b: IN INTEGER; s, cout: OUT STD_LOGIC_VECTOR);
   
END funcs;


--------------------------- B O D Y ----------------------------


PACKAGE BODY funcs IS

-----------------------------------------------------------------
-- utility functions
-----------------------------------------------------------------

   FUNCTION TO_STDLOGIC(arg1: BOOLEAN) RETURN STD_LOGIC IS
     BEGIN IF arg1 THEN RETURN '1'; ELSE RETURN '0'; END IF; END;
--   FUNCTION TO_STDLOGIC(arg1: STD_ULOGIC_VECTOR(0 DOWNTO 0)) RETURN STD_LOGIC IS
--     BEGIN RETURN arg1(0); END;
   FUNCTION TO_STDLOGIC(arg1: STD_LOGIC_VECTOR(0 DOWNTO 0)) RETURN STD_LOGIC IS
     BEGIN RETURN arg1(0); END;
   FUNCTION TO_STDLOGIC(arg1: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN arg1(0); END;
   FUNCTION TO_STDLOGIC(arg1: SIGNED(0 DOWNTO 0)) RETURN STD_LOGIC IS
     BEGIN RETURN arg1(0); END;

   FUNCTION TO_STDLOGICVECTOR(arg1: STD_LOGIC) RETURN STD_LOGIC_VECTOR IS
     VARIABLE result: STD_LOGIC_VECTOR(0 DOWNTO 0);
   BEGIN
     result := (0 => arg1);
     RETURN result;
   END;

   FUNCTION maximum (arg1,arg2: INTEGER) RETURN INTEGER IS
   BEGIN
     IF(arg1 > arg2) THEN
       RETURN(arg1) ;
     ELSE
       RETURN(arg2) ;
     END IF;
   END;

   FUNCTION minimum (arg1,arg2: INTEGER) RETURN INTEGER IS
   BEGIN
     IF(arg1 < arg2) THEN
       RETURN(arg1) ;
     ELSE
       RETURN(arg2) ;
     END IF;
   END;

   FUNCTION ifeqsel(arg1, arg2, seleq, selne : INTEGER) RETURN INTEGER IS
   BEGIN
     IF(arg1 = arg2) THEN
       RETURN(seleq) ;
     ELSE
       RETURN(selne) ;
     END IF;
   END;

   FUNCTION resolve_std_logic_vector(input1: STD_LOGIC_VECTOR; input2: STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR IS
     CONSTANT len: INTEGER := input1'LENGTH;
     ALIAS input1a: STD_LOGIC_VECTOR(len-1 DOWNTO 0) IS input1;
     ALIAS input2a: STD_LOGIC_VECTOR(len-1 DOWNTO 0) IS input2;
     VARIABLE result: STD_LOGIC_VECTOR(len-1 DOWNTO 0);
   BEGIN
     result := (others => '0');
     --synopsys translate_off
     FOR i IN len-1 DOWNTO 0 LOOP
       result(i) := resolved(input1a(i) & input2a(i));
     END LOOP;
     --synopsys translate_on
     RETURN result;
   END;

   FUNCTION resolve_unsigned(input1: UNSIGNED; input2: UNSIGNED) RETURN UNSIGNED IS
   BEGIN RETURN UNSIGNED(resolve_std_logic_vector(STD_LOGIC_VECTOR(input1), STD_LOGIC_VECTOR(input2))); END;

   FUNCTION resolve_signed(input1: SIGNED; input2: SIGNED) RETURN SIGNED IS
   BEGIN RETURN SIGNED(resolve_std_logic_vector(STD_LOGIC_VECTOR(input1), STD_LOGIC_VECTOR(input2))); END;

-----------------------------------------------------------------
-- Logic Functions
-----------------------------------------------------------------

   FUNCTION "not"(arg1: UNSIGNED) RETURN UNSIGNED IS
     BEGIN RETURN UNSIGNED(not STD_LOGIC_VECTOR(arg1)); END;
   FUNCTION and_s(inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
     BEGIN RETURN TO_STDLOGIC(and_v(inputs, 1)); END;
   FUNCTION or_s (inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
     BEGIN RETURN TO_STDLOGIC(or_v(inputs, 1)); END;
   FUNCTION xor_s(inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
     BEGIN RETURN TO_STDLOGIC(xor_v(inputs, 1)); END;

   FUNCTION and_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR IS
     CONSTANT ilen: POSITIVE := inputs'LENGTH;
     CONSTANT ilenM1: POSITIVE := ilen-1; --2.1.6.3
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT ilenMolenM1: INTEGER := ilen-olen-1; --2.1.6.3
     VARIABLE inputsx: STD_LOGIC_VECTOR(ilen-1 DOWNTO 0);
     CONSTANT icnt2: POSITIVE:= inputs'LENGTH/olen;
     VARIABLE result: STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT ilen REM olen = 0 SEVERITY FAILURE;
     --synopsys translate_on
     inputsx := inputs;
     result := inputsx(olenM1 DOWNTO 0);
     FOR i IN icnt2-1 DOWNTO 1 LOOP
       inputsx(ilenMolenM1 DOWNTO 0) := inputsx(ilenM1 DOWNTO olen);
       result := result AND inputsx(olenM1 DOWNTO 0);
     END LOOP;
     RETURN result;
   END;

   FUNCTION or_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR IS
     CONSTANT ilen: POSITIVE := inputs'LENGTH;
     CONSTANT ilenM1: POSITIVE := ilen-1; --2.1.6.3
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT ilenMolenM1: INTEGER := ilen-olen-1; --2.1.6.3
     VARIABLE inputsx: STD_LOGIC_VECTOR(ilen-1 DOWNTO 0);
     CONSTANT icnt2: POSITIVE:= inputs'LENGTH/olen;
     VARIABLE result: STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT ilen REM olen = 0 SEVERITY FAILURE;
     --synopsys translate_on
     inputsx := inputs;
     result := inputsx(olenM1 DOWNTO 0);
     -- this if is added as a quick fix for a bug in catapult evaluating the loop even if inputs'LENGTH==1
     -- see dts0100971279
     IF icnt2 > 1 THEN
       FOR i IN icnt2-1 DOWNTO 1 LOOP
         inputsx(ilenMolenM1 DOWNTO 0) := inputsx(ilenM1 DOWNTO olen);
         result := result OR inputsx(olenM1 DOWNTO 0);
       END LOOP;
     END IF;
     RETURN result;
   END;

   FUNCTION xor_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR IS
     CONSTANT ilen: POSITIVE := inputs'LENGTH;
     CONSTANT ilenM1: POSITIVE := ilen-1; --2.1.6.3
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT ilenMolenM1: INTEGER := ilen-olen-1; --2.1.6.3
     VARIABLE inputsx: STD_LOGIC_VECTOR(ilen-1 DOWNTO 0);
     CONSTANT icnt2: POSITIVE:= inputs'LENGTH/olen;
     VARIABLE result: STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT ilen REM olen = 0 SEVERITY FAILURE;
     --synopsys translate_on
     inputsx := inputs;
     result := inputsx(olenM1 DOWNTO 0);
     FOR i IN icnt2-1 DOWNTO 1 LOOP
       inputsx(ilenMolenM1 DOWNTO 0) := inputsx(ilenM1 DOWNTO olen);
       result := result XOR inputsx(olenM1 DOWNTO 0);
     END LOOP;
     RETURN result;
   END;

-----------------------------------------------------------------
-- Muxes
-----------------------------------------------------------------
   
   FUNCTION mux_sel2_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(1 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 4;
     ALIAS    inputs0: STD_LOGIC_VECTOR( inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector( size-1 DOWNTO 0);
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "00" =>
       result := inputs0(1*size-1 DOWNTO 0*size);
     WHEN "01" =>
       result := inputs0(2*size-1 DOWNTO 1*size);
     WHEN "10" =>
       result := inputs0(3*size-1 DOWNTO 2*size);
     WHEN "11" =>
       result := inputs0(4*size-1 DOWNTO 3*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;
   
   FUNCTION mux_sel3_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(2 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 8;
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector(size-1 DOWNTO 0);
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "000" =>
       result := inputs0(1*size-1 DOWNTO 0*size);
     WHEN "001" =>
       result := inputs0(2*size-1 DOWNTO 1*size);
     WHEN "010" =>
       result := inputs0(3*size-1 DOWNTO 2*size);
     WHEN "011" =>
       result := inputs0(4*size-1 DOWNTO 3*size);
     WHEN "100" =>
       result := inputs0(5*size-1 DOWNTO 4*size);
     WHEN "101" =>
       result := inputs0(6*size-1 DOWNTO 5*size);
     WHEN "110" =>
       result := inputs0(7*size-1 DOWNTO 6*size);
     WHEN "111" =>
       result := inputs0(8*size-1 DOWNTO 7*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;
   
   FUNCTION mux_sel4_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(3 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 16;
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector(size-1 DOWNTO 0);
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "0000" =>
       result := inputs0( 1*size-1 DOWNTO 0*size);
     WHEN "0001" =>
       result := inputs0( 2*size-1 DOWNTO 1*size);
     WHEN "0010" =>
       result := inputs0( 3*size-1 DOWNTO 2*size);
     WHEN "0011" =>
       result := inputs0( 4*size-1 DOWNTO 3*size);
     WHEN "0100" =>
       result := inputs0( 5*size-1 DOWNTO 4*size);
     WHEN "0101" =>
       result := inputs0( 6*size-1 DOWNTO 5*size);
     WHEN "0110" =>
       result := inputs0( 7*size-1 DOWNTO 6*size);
     WHEN "0111" =>
       result := inputs0( 8*size-1 DOWNTO 7*size);
     WHEN "1000" =>
       result := inputs0( 9*size-1 DOWNTO 8*size);
     WHEN "1001" =>
       result := inputs0( 10*size-1 DOWNTO 9*size);
     WHEN "1010" =>
       result := inputs0( 11*size-1 DOWNTO 10*size);
     WHEN "1011" =>
       result := inputs0( 12*size-1 DOWNTO 11*size);
     WHEN "1100" =>
       result := inputs0( 13*size-1 DOWNTO 12*size);
     WHEN "1101" =>
       result := inputs0( 14*size-1 DOWNTO 13*size);
     WHEN "1110" =>
       result := inputs0( 15*size-1 DOWNTO 14*size);
     WHEN "1111" =>
       result := inputs0( 16*size-1 DOWNTO 15*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;
   
   FUNCTION mux_sel5_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(4 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 32;
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector(size-1 DOWNTO 0 );
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "00000" =>
       result := inputs0( 1*size-1 DOWNTO 0*size);
     WHEN "00001" =>
       result := inputs0( 2*size-1 DOWNTO 1*size);
     WHEN "00010" =>
       result := inputs0( 3*size-1 DOWNTO 2*size);
     WHEN "00011" =>
       result := inputs0( 4*size-1 DOWNTO 3*size);
     WHEN "00100" =>
       result := inputs0( 5*size-1 DOWNTO 4*size);
     WHEN "00101" =>
       result := inputs0( 6*size-1 DOWNTO 5*size);
     WHEN "00110" =>
       result := inputs0( 7*size-1 DOWNTO 6*size);
     WHEN "00111" =>
       result := inputs0( 8*size-1 DOWNTO 7*size);
     WHEN "01000" =>
       result := inputs0( 9*size-1 DOWNTO 8*size);
     WHEN "01001" =>
       result := inputs0( 10*size-1 DOWNTO 9*size);
     WHEN "01010" =>
       result := inputs0( 11*size-1 DOWNTO 10*size);
     WHEN "01011" =>
       result := inputs0( 12*size-1 DOWNTO 11*size);
     WHEN "01100" =>
       result := inputs0( 13*size-1 DOWNTO 12*size);
     WHEN "01101" =>
       result := inputs0( 14*size-1 DOWNTO 13*size);
     WHEN "01110" =>
       result := inputs0( 15*size-1 DOWNTO 14*size);
     WHEN "01111" =>
       result := inputs0( 16*size-1 DOWNTO 15*size);
     WHEN "10000" =>
       result := inputs0( 17*size-1 DOWNTO 16*size);
     WHEN "10001" =>
       result := inputs0( 18*size-1 DOWNTO 17*size);
     WHEN "10010" =>
       result := inputs0( 19*size-1 DOWNTO 18*size);
     WHEN "10011" =>
       result := inputs0( 20*size-1 DOWNTO 19*size);
     WHEN "10100" =>
       result := inputs0( 21*size-1 DOWNTO 20*size);
     WHEN "10101" =>
       result := inputs0( 22*size-1 DOWNTO 21*size);
     WHEN "10110" =>
       result := inputs0( 23*size-1 DOWNTO 22*size);
     WHEN "10111" =>
       result := inputs0( 24*size-1 DOWNTO 23*size);
     WHEN "11000" =>
       result := inputs0( 25*size-1 DOWNTO 24*size);
     WHEN "11001" =>
       result := inputs0( 26*size-1 DOWNTO 25*size);
     WHEN "11010" =>
       result := inputs0( 27*size-1 DOWNTO 26*size);
     WHEN "11011" =>
       result := inputs0( 28*size-1 DOWNTO 27*size);
     WHEN "11100" =>
       result := inputs0( 29*size-1 DOWNTO 28*size);
     WHEN "11101" =>
       result := inputs0( 30*size-1 DOWNTO 29*size);
     WHEN "11110" =>
       result := inputs0( 31*size-1 DOWNTO 30*size);
     WHEN "11111" =>
       result := inputs0( 32*size-1 DOWNTO 31*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;
   
   FUNCTION mux_sel6_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(5 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 64;
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector(size-1 DOWNTO 0);
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "000000" =>
       result := inputs0( 1*size-1 DOWNTO 0*size);
     WHEN "000001" =>
       result := inputs0( 2*size-1 DOWNTO 1*size);
     WHEN "000010" =>
       result := inputs0( 3*size-1 DOWNTO 2*size);
     WHEN "000011" =>
       result := inputs0( 4*size-1 DOWNTO 3*size);
     WHEN "000100" =>
       result := inputs0( 5*size-1 DOWNTO 4*size);
     WHEN "000101" =>
       result := inputs0( 6*size-1 DOWNTO 5*size);
     WHEN "000110" =>
       result := inputs0( 7*size-1 DOWNTO 6*size);
     WHEN "000111" =>
       result := inputs0( 8*size-1 DOWNTO 7*size);
     WHEN "001000" =>
       result := inputs0( 9*size-1 DOWNTO 8*size);
     WHEN "001001" =>
       result := inputs0( 10*size-1 DOWNTO 9*size);
     WHEN "001010" =>
       result := inputs0( 11*size-1 DOWNTO 10*size);
     WHEN "001011" =>
       result := inputs0( 12*size-1 DOWNTO 11*size);
     WHEN "001100" =>
       result := inputs0( 13*size-1 DOWNTO 12*size);
     WHEN "001101" =>
       result := inputs0( 14*size-1 DOWNTO 13*size);
     WHEN "001110" =>
       result := inputs0( 15*size-1 DOWNTO 14*size);
     WHEN "001111" =>
       result := inputs0( 16*size-1 DOWNTO 15*size);
     WHEN "010000" =>
       result := inputs0( 17*size-1 DOWNTO 16*size);
     WHEN "010001" =>
       result := inputs0( 18*size-1 DOWNTO 17*size);
     WHEN "010010" =>
       result := inputs0( 19*size-1 DOWNTO 18*size);
     WHEN "010011" =>
       result := inputs0( 20*size-1 DOWNTO 19*size);
     WHEN "010100" =>
       result := inputs0( 21*size-1 DOWNTO 20*size);
     WHEN "010101" =>
       result := inputs0( 22*size-1 DOWNTO 21*size);
     WHEN "010110" =>
       result := inputs0( 23*size-1 DOWNTO 22*size);
     WHEN "010111" =>
       result := inputs0( 24*size-1 DOWNTO 23*size);
     WHEN "011000" =>
       result := inputs0( 25*size-1 DOWNTO 24*size);
     WHEN "011001" =>
       result := inputs0( 26*size-1 DOWNTO 25*size);
     WHEN "011010" =>
       result := inputs0( 27*size-1 DOWNTO 26*size);
     WHEN "011011" =>
       result := inputs0( 28*size-1 DOWNTO 27*size);
     WHEN "011100" =>
       result := inputs0( 29*size-1 DOWNTO 28*size);
     WHEN "011101" =>
       result := inputs0( 30*size-1 DOWNTO 29*size);
     WHEN "011110" =>
       result := inputs0( 31*size-1 DOWNTO 30*size);
     WHEN "011111" =>
       result := inputs0( 32*size-1 DOWNTO 31*size);
     WHEN "100000" =>
       result := inputs0( 33*size-1 DOWNTO 32*size);
     WHEN "100001" =>
       result := inputs0( 34*size-1 DOWNTO 33*size);
     WHEN "100010" =>
       result := inputs0( 35*size-1 DOWNTO 34*size);
     WHEN "100011" =>
       result := inputs0( 36*size-1 DOWNTO 35*size);
     WHEN "100100" =>
       result := inputs0( 37*size-1 DOWNTO 36*size);
     WHEN "100101" =>
       result := inputs0( 38*size-1 DOWNTO 37*size);
     WHEN "100110" =>
       result := inputs0( 39*size-1 DOWNTO 38*size);
     WHEN "100111" =>
       result := inputs0( 40*size-1 DOWNTO 39*size);
     WHEN "101000" =>
       result := inputs0( 41*size-1 DOWNTO 40*size);
     WHEN "101001" =>
       result := inputs0( 42*size-1 DOWNTO 41*size);
     WHEN "101010" =>
       result := inputs0( 43*size-1 DOWNTO 42*size);
     WHEN "101011" =>
       result := inputs0( 44*size-1 DOWNTO 43*size);
     WHEN "101100" =>
       result := inputs0( 45*size-1 DOWNTO 44*size);
     WHEN "101101" =>
       result := inputs0( 46*size-1 DOWNTO 45*size);
     WHEN "101110" =>
       result := inputs0( 47*size-1 DOWNTO 46*size);
     WHEN "101111" =>
       result := inputs0( 48*size-1 DOWNTO 47*size);
     WHEN "110000" =>
       result := inputs0( 49*size-1 DOWNTO 48*size);
     WHEN "110001" =>
       result := inputs0( 50*size-1 DOWNTO 49*size);
     WHEN "110010" =>
       result := inputs0( 51*size-1 DOWNTO 50*size);
     WHEN "110011" =>
       result := inputs0( 52*size-1 DOWNTO 51*size);
     WHEN "110100" =>
       result := inputs0( 53*size-1 DOWNTO 52*size);
     WHEN "110101" =>
       result := inputs0( 54*size-1 DOWNTO 53*size);
     WHEN "110110" =>
       result := inputs0( 55*size-1 DOWNTO 54*size);
     WHEN "110111" =>
       result := inputs0( 56*size-1 DOWNTO 55*size);
     WHEN "111000" =>
       result := inputs0( 57*size-1 DOWNTO 56*size);
     WHEN "111001" =>
       result := inputs0( 58*size-1 DOWNTO 57*size);
     WHEN "111010" =>
       result := inputs0( 59*size-1 DOWNTO 58*size);
     WHEN "111011" =>
       result := inputs0( 60*size-1 DOWNTO 59*size);
     WHEN "111100" =>
       result := inputs0( 61*size-1 DOWNTO 60*size);
     WHEN "111101" =>
       result := inputs0( 62*size-1 DOWNTO 61*size);
     WHEN "111110" =>
       result := inputs0( 63*size-1 DOWNTO 62*size);
     WHEN "111111" =>
       result := inputs0( 64*size-1 DOWNTO 63*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;

   FUNCTION mux_s(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC) RETURN STD_LOGIC IS
   BEGIN RETURN TO_STDLOGIC(mux_v(inputs, sel)); END;

   FUNCTION mux_s(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
   BEGIN RETURN TO_STDLOGIC(mux_v(inputs, sel)); END;

   FUNCTION mux_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC) RETURN STD_LOGIC_VECTOR IS  --pragma hls_map_to_operator mux
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     CONSTANT size   : POSITIVE := inputs'LENGTH / 2;
     CONSTANT olen   : POSITIVE := inputs'LENGTH / 2;
     VARIABLE result : STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT inputs'LENGTH = olen * 2 SEVERITY FAILURE;
     --synopsys translate_on
       CASE sel IS
       WHEN '1'
     --synopsys translate_off
            | 'H'
     --synopsys translate_on
            =>
         result := inputs0( size-1 DOWNTO 0);
       WHEN '0' 
     --synopsys translate_off
            | 'L'
     --synopsys translate_on
            =>
         result := inputs0(2*size-1  DOWNTO size);
       WHEN others =>
         --synopsys translate_off
         result := resolve_std_logic_vector(inputs0(size-1 DOWNTO 0), inputs0( 2*size-1 DOWNTO size));
         --synopsys translate_on
       END CASE;
       RETURN result;
   END;
--   BEGIN RETURN mux_v(inputs, TO_STDLOGICVECTOR(sel)); END;

   FUNCTION mux_v(inputs: STD_LOGIC_VECTOR; sel : STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR IS --pragma hls_map_to_operator mux
     ALIAS    inputs0: STD_LOGIC_VECTOR( inputs'LENGTH-1 DOWNTO 0) IS inputs;
     ALIAS    sel0   : STD_LOGIC_VECTOR( sel'LENGTH-1 DOWNTO 0 ) IS sel;

     VARIABLE sellen : INTEGER RANGE 2-sel'LENGTH TO sel'LENGTH;
     CONSTANT size   : POSITIVE := inputs'LENGTH / 2;
     CONSTANT olen   : POSITIVE := inputs'LENGTH / 2**sel'LENGTH;
     VARIABLE result : STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
     TYPE inputs_array_type is array(natural range <>) of std_logic_vector( olen - 1 DOWNTO 0);
     VARIABLE inputs_array : inputs_array_type( 2**sel'LENGTH - 1 DOWNTO 0);
   BEGIN
     sellen := sel'LENGTH;
     --synopsys translate_off
     ASSERT inputs'LENGTH = olen * 2**sellen SEVERITY FAILURE;
     sellen := 2-sellen;
     --synopsys translate_on
     CASE sellen IS
     WHEN 1 =>
       CASE sel0(0) IS

       WHEN '1' 
     --synopsys translate_off
            | 'H'
     --synopsys translate_on
            =>
         result := inputs0(  size-1 DOWNTO 0);
       WHEN '0' 
     --synopsys translate_off
            | 'L'
     --synopsys translate_on
            =>
         result := inputs0(2*size-1 DOWNTO size);
       WHEN others =>
         --synopsys translate_off
         result := resolve_std_logic_vector(inputs0( size-1 DOWNTO 0), inputs0( 2*size-1 DOWNTO size));
         --synopsys translate_on
       END CASE;
     WHEN 2 =>
       result := mux_sel2_v(inputs, not sel);
     WHEN 3 =>
       result := mux_sel3_v(inputs, not sel);
     WHEN 4 =>
       result := mux_sel4_v(inputs, not sel);
     WHEN 5 =>
       result := mux_sel5_v(inputs, not sel);
     WHEN 6 =>
       result := mux_sel6_v(inputs, not sel);
     WHEN others =>
       -- synopsys translate_off
       IF(Is_X(sel0)) THEN
         result := (others => 'X');
       ELSE
       -- synopsys translate_on
         FOR i in 0 to 2**sel'LENGTH - 1 LOOP
           inputs_array(i) := inputs0( ((i + 1) * olen) - 1  DOWNTO i*olen);
         END LOOP;
         result := inputs_array(CONV_INTEGER( (UNSIGNED(NOT sel0)) ));
       -- synopsys translate_off
       END IF;
       -- synopsys translate_on
     END CASE;
     RETURN result;
   END;

 
-----------------------------------------------------------------
-- Latches
-----------------------------------------------------------------

   FUNCTION lat_s(dinput: STD_LOGIC; clk: STD_LOGIC; doutput: STD_LOGIC) RETURN STD_LOGIC IS
   BEGIN RETURN mux_s(STD_LOGIC_VECTOR'(doutput & dinput), clk); END;

   FUNCTION lat_v(dinput: STD_LOGIC_VECTOR ; clk: STD_LOGIC; doutput: STD_LOGIC_VECTOR ) RETURN STD_LOGIC_VECTOR IS
   BEGIN
     --synopsys translate_off
     ASSERT dinput'LENGTH = doutput'LENGTH SEVERITY FAILURE;
     --synopsys translate_on
     RETURN mux_v(doutput & dinput, clk);
   END;

-----------------------------------------------------------------
-- Tri-States
-----------------------------------------------------------------
--   FUNCTION tri_s(dinput: STD_LOGIC; control: STD_LOGIC) RETURN STD_LOGIC IS
--   BEGIN RETURN TO_STDLOGIC(tri_v(TO_STDLOGICVECTOR(dinput), control)); END;
--
--   FUNCTION tri_v(dinput: STD_LOGIC_VECTOR ; control: STD_LOGIC) RETURN STD_LOGIC_VECTOR IS
--     VARIABLE result: STD_LOGIC_VECTOR(dinput'range);
--   BEGIN
--     CASE control IS
--     WHEN '0' | 'L' =>
--       result := (others => 'Z');
--     WHEN '1' | 'H' =>
--       FOR i IN dinput'range LOOP
--         result(i) := to_UX01(dinput(i));
--       END LOOP;
--     WHEN others =>
--       -- synopsys translate_off
--       result := (others => 'X');
--       -- synopsys translate_on
--     END CASE;
--     RETURN result;
--   END;

-----------------------------------------------------------------
-- compare functions returning STD_LOGIC
-- in contrast to the functions returning boolean
-----------------------------------------------------------------

   FUNCTION "=" (l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN not or_s(STD_LOGIC_VECTOR(l) xor STD_LOGIC_VECTOR(r)); END;
   FUNCTION "=" (l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN not or_s(STD_LOGIC_VECTOR(l) xor STD_LOGIC_VECTOR(r)); END;
   FUNCTION "/="(l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN or_s(STD_LOGIC_VECTOR(l) xor STD_LOGIC_VECTOR(r)); END;
   FUNCTION "/="(l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN or_s(STD_LOGIC_VECTOR(l) xor STD_LOGIC_VECTOR(r)); END;

   FUNCTION "<" (l, r: UNSIGNED) RETURN STD_LOGIC IS
     VARIABLE diff: UNSIGNED(l'LENGTH DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT l'LENGTH = r'LENGTH SEVERITY FAILURE;
     --synopsys translate_on
     diff := ('0'&l) - ('0'&r);
     RETURN diff(l'LENGTH);
   END;
   FUNCTION "<"(l, r: SIGNED  ) RETURN STD_LOGIC IS
   BEGIN
     RETURN (UNSIGNED(l) < UNSIGNED(r)) xor (l(l'LEFT) xor r(r'LEFT));
   END;

   FUNCTION "<="(l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN not STD_LOGIC'(r < l); END;
   FUNCTION "<=" (l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN not STD_LOGIC'(r < l); END;
   FUNCTION ">" (l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN r < l; END;
   FUNCTION ">"(l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN r < l; END;
   FUNCTION ">="(l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN not STD_LOGIC'(l < r); END;
   FUNCTION ">=" (l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN not STD_LOGIC'(l < r); END;

   FUNCTION cmp (l, r: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
   BEGIN
     --synopsys translate_off
     ASSERT l'LENGTH = r'LENGTH SEVERITY FAILURE;
     --synopsys translate_on
     RETURN not or_s(l xor r);
   END;

-----------------------------------------------------------------
-- Vectorized Overloaded Arithmetic Operators
-----------------------------------------------------------------

   --some functions to placate spyglass
   FUNCTION mult_natural(a,b : NATURAL) RETURN NATURAL IS
   BEGIN
     return a*b;
   END mult_natural;

   FUNCTION div_natural(a,b : NATURAL) RETURN NATURAL IS
   BEGIN
     return a/b;
   END div_natural;

   FUNCTION mod_natural(a,b : NATURAL) RETURN NATURAL IS
   BEGIN
     return a mod b;
   END mod_natural;

   FUNCTION add_unsigned(a,b : UNSIGNED) RETURN UNSIGNED IS
   BEGIN
     return a+b;
   END add_unsigned;

   FUNCTION sub_unsigned(a,b : UNSIGNED) RETURN UNSIGNED IS
   BEGIN
     return a-b;
   END sub_unsigned;

   FUNCTION sub_int(a,b : INTEGER) RETURN INTEGER IS
   BEGIN
     return a-b;
   END sub_int;

   FUNCTION concat_0(b : UNSIGNED) RETURN UNSIGNED IS
   BEGIN
     return '0' & b;
   END concat_0;

   FUNCTION concat_uns(a,b : UNSIGNED) RETURN UNSIGNED IS
   BEGIN
     return a&b;
   END concat_uns;

   FUNCTION concat_vect(a,b : STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR IS
   BEGIN
     return a&b;
   END concat_vect;





   FUNCTION faccu(arg: UNSIGNED; width: NATURAL) RETURN UNSIGNED IS
     CONSTANT ninps : NATURAL := arg'LENGTH / width;
     ALIAS    arg0  : UNSIGNED(arg'LENGTH-1 DOWNTO 0) IS arg;
     VARIABLE result: UNSIGNED(width-1 DOWNTO 0);
     VARIABLE from  : INTEGER;
     VARIABLE dto   : INTEGER;
   BEGIN
     --synopsys translate_off
     ASSERT arg'LENGTH = width * ninps SEVERITY FAILURE;
     --synopsys translate_on
     result := (OTHERS => '0');
     FOR i IN ninps-1 DOWNTO 0 LOOP
       --result := result + arg0((i+1)*width-1 DOWNTO i*width);
       from := mult_natural((i+1), width)-1; --2.1.6.3
       dto  := mult_natural(i,width); --2.1.6.3
       result := add_unsigned(result , arg0(from DOWNTO dto) );
     END LOOP;
     RETURN result;
   END faccu;

   FUNCTION  fabs (arg1: SIGNED) RETURN UNSIGNED IS
   BEGIN
     CASE arg1(arg1'LEFT) IS
     WHEN '1'
     --synopsys translate_off
          | 'H'
     --synopsys translate_on
       =>
       RETURN UNSIGNED'("0") - UNSIGNED(arg1);
     WHEN '0'
     --synopsys translate_off
          | 'L'
     --synopsys translate_on
       =>
       RETURN UNSIGNED(arg1);
     WHEN others =>
       RETURN resolve_unsigned(UNSIGNED(arg1), UNSIGNED'("0") - UNSIGNED(arg1));
     END CASE;
   END;

   PROCEDURE divmod(l, r: UNSIGNED; rdiv, rmod: OUT UNSIGNED) IS
     CONSTANT llen: INTEGER := l'LENGTH;
     CONSTANT rlen: INTEGER := r'LENGTH;
     CONSTANT llen_plus_rlen: INTEGER := llen + rlen;
     VARIABLE lbuf: UNSIGNED(llen+rlen-1 DOWNTO 0);
     VARIABLE diff: UNSIGNED(rlen DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT rdiv'LENGTH = llen AND rmod'LENGTH = rlen SEVERITY FAILURE;
     --synopsys translate_on
     lbuf := (others => '0');
     lbuf(llen-1 DOWNTO 0) := l;
     FOR i IN rdiv'range LOOP
       diff := sub_unsigned(lbuf(llen_plus_rlen-1 DOWNTO llen-1) ,(concat_0(r)));
       rdiv(i) := not diff(rlen);
       IF diff(rlen) = '0' THEN
         lbuf(llen_plus_rlen-1 DOWNTO llen-1) := diff;
       END IF;
       lbuf(llen_plus_rlen-1 DOWNTO 1) := lbuf(llen_plus_rlen-2 DOWNTO 0);
     END LOOP;
     rmod := lbuf(llen_plus_rlen-1 DOWNTO llen);
   END divmod;

   FUNCTION "/"  (l, r: UNSIGNED) RETURN UNSIGNED IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
   BEGIN
     divmod(l, r, rdiv, rmod);
     RETURN rdiv;
   END "/";

   FUNCTION "MOD"(l, r: UNSIGNED) RETURN UNSIGNED IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
   BEGIN
     divmod(l, r, rdiv, rmod);
     RETURN rmod;
   END;

   FUNCTION "REM"(l, r: UNSIGNED) RETURN UNSIGNED IS
     BEGIN RETURN l MOD r; END;

   FUNCTION "/"  (l, r: SIGNED  ) RETURN SIGNED  IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
   BEGIN
     divmod(fabs(l), fabs(r), rdiv, rmod);
     IF to_X01(l(l'LEFT)) /= to_X01(r(r'LEFT)) THEN
       rdiv := UNSIGNED'("0") - rdiv;
     END IF;
     RETURN SIGNED(rdiv); -- overflow problem "1000" / "11"
   END "/";

   FUNCTION "MOD"(l, r: SIGNED  ) RETURN SIGNED  IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
     CONSTANT rnul: UNSIGNED(r'LENGTH-1 DOWNTO 0) := (others => '0');
   BEGIN
     divmod(fabs(l), fabs(r), rdiv, rmod);
     IF to_X01(l(l'LEFT)) = '1' THEN
       rmod := UNSIGNED'("0") - rmod;
     END IF;
     IF rmod /= rnul AND to_X01(l(l'LEFT)) /= to_X01(r(r'LEFT)) THEN
       rmod := UNSIGNED(r) + rmod;
     END IF;
     RETURN SIGNED(rmod);
   END "MOD";

   FUNCTION "REM"(l, r: SIGNED  ) RETURN SIGNED  IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
   BEGIN
     divmod(fabs(l), fabs(r), rdiv, rmod);
     IF to_X01(l(l'LEFT)) = '1' THEN
       rmod := UNSIGNED'("0") - rmod;
     END IF;
     RETURN SIGNED(rmod);
   END "REM";

   FUNCTION mult_unsigned(l,r : UNSIGNED) return UNSIGNED is
   BEGIN
     return l*r; 
   END mult_unsigned;

   FUNCTION "**" (l, r : UNSIGNED) RETURN UNSIGNED IS
     CONSTANT llen  : NATURAL := l'LENGTH;
     VARIABLE result: UNSIGNED(llen-1 DOWNTO 0);
     VARIABLE fak   : UNSIGNED(llen-1 DOWNTO 0);
   BEGIN
     fak := l;
     result := (others => '0'); result(0) := '1';
     FOR i IN r'reverse_range LOOP
       --was:result := UNSIGNED(mux_v(STD_LOGIC_VECTOR(result & (result*fak)), r(i)));
       result := UNSIGNED(mux_v(STD_LOGIC_VECTOR( concat_uns(result , mult_unsigned(result,fak) )), r(i)));

       fak := mult_unsigned(fak , fak);
     END LOOP;
     RETURN result;
   END "**";

   FUNCTION "**" (l, r : SIGNED) RETURN SIGNED IS
     CONSTANT rlen  : NATURAL := r'LENGTH;
     ALIAS    r0    : SIGNED(0 TO r'LENGTH-1) IS r;
     VARIABLE result: SIGNED(l'range);
   BEGIN
     CASE r(r'LEFT) IS
     WHEN '0'
   --synopsys translate_off
          | 'L'
   --synopsys translate_on
     =>
       result := SIGNED(UNSIGNED(l) ** UNSIGNED(r0(1 TO r'LENGTH-1)));
     WHEN '1'
   --synopsys translate_off
          | 'H'
   --synopsys translate_on
     =>
       result := (others => '0');
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END "**";

-----------------------------------------------------------------
--               S H I F T   F U C T I O N S
-- negative shift shifts the opposite direction
-----------------------------------------------------------------

   FUNCTION add_nat(arg1 : NATURAL; arg2 : NATURAL ) RETURN NATURAL IS
   BEGIN
     return (arg1 + arg2);
   END;
   
--   FUNCTION UNSIGNED_2_BIT_VECTOR(arg1 : NATURAL; arg2 : NATURAL ) RETURN BIT_VECTOR IS
--   BEGIN
--     return (arg1 + arg2);
--   END;
   
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
     CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
   BEGIN
     result := (others => sbit);
     result(ilenub DOWNTO 0) := arg1;
     result := shl(result, arg2);
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshl_stdar(arg1: SIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
     CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: SIGNED(len-1 DOWNTO 0);
   BEGIN
     result := (others => sbit);
     result(ilenub DOWNTO 0) := arg1;
     result := shl(SIGNED(result), arg2);
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
     CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
   BEGIN
     result := (others => sbit);
     result(ilenub DOWNTO 0) := arg1;
     result := shr(result, arg2);
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshr_stdar(arg1: SIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
     CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: SIGNED(len-1 DOWNTO 0);
   BEGIN
     result := (others => sbit);
     result(ilenub DOWNTO 0) := arg1;
     result := shr(result, arg2);
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT arg1l: NATURAL := arg1'LENGTH - 1;
     ALIAS    arg1x: UNSIGNED(arg1l DOWNTO 0) IS arg1;
     CONSTANT arg2l: NATURAL := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE arg1x_pad: UNSIGNED(arg1l+1 DOWNTO 0);
     VARIABLE result: UNSIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others=>'0');
     arg1x_pad(arg1l+1) := sbit;
     arg1x_pad(arg1l downto 0) := arg1x;
     IF arg2l = 0 THEN
       RETURN fshr_stdar(arg1x_pad, UNSIGNED(arg2x), sbit, olen);
     -- ELSIF arg1l = 0 THEN
     --   RETURN fshl(sbit & arg1x, arg2x, sbit, olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
     --synopsys translate_off
            | 'L'
     --synopsys translate_on
       =>
         RETURN fshl_stdar(arg1x_pad, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN '1'
     --synopsys translate_off
            | 'H'
     --synopsys translate_on
       =>
         RETURN fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_unsigned(
           fshl_stdar(arg1x, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit,  olen),
           fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen)
         );
         --synopsys translate_on
         RETURN result;
       END CASE;
     END IF;
   END;

   FUNCTION fshl_stdar(arg1: SIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
     CONSTANT arg1l: NATURAL := arg1'LENGTH - 1;
     ALIAS    arg1x: SIGNED(arg1l DOWNTO 0) IS arg1;
     CONSTANT arg2l: NATURAL := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE arg1x_pad: SIGNED(arg1l+1 DOWNTO 0);
     VARIABLE result: SIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others=>'0');
     arg1x_pad(arg1l+1) := sbit;
     arg1x_pad(arg1l downto 0) := arg1x;
     IF arg2l = 0 THEN
       RETURN fshr_stdar(arg1x_pad, UNSIGNED(arg2x), sbit, olen);
     -- ELSIF arg1l = 0 THEN
     --   RETURN fshl(sbit & arg1x, arg2x, sbit, olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
       =>
         RETURN fshl_stdar(arg1x_pad, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
       =>
         RETURN fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_signed(
           fshl_stdar(arg1x, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit,  olen),
           fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen)
         );
         --synopsys translate_on
         RETURN result;
       END CASE;
     END IF;
   END;

   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT arg2l: INTEGER := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE result: UNSIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others => '0');
     IF arg2l = 0 THEN
       RETURN fshl_stdar(arg1, UNSIGNED(arg2x), olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
        =>
         RETURN fshr_stdar(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
        =>
         RETURN fshl_stdar(arg1 & '0', '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_unsigned(
           fshr_stdar(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen),
           fshl_stdar(arg1 & '0', '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen)
         );
         --synopsys translate_on
	 return result;
       END CASE;
     END IF;
   END;

   FUNCTION fshr_stdar(arg1: SIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
     CONSTANT arg2l: INTEGER := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE result: SIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others => '0');
     IF arg2l = 0 THEN
       RETURN fshl_stdar(arg1, UNSIGNED(arg2x), olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
       =>
         RETURN fshr_stdar(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
       =>
         RETURN fshl_stdar(arg1 & '0', '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_signed(
           fshr_stdar(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen),
           fshl_stdar(arg1 & '0', '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen)
         );
         --synopsys translate_on
	 return result;
       END CASE;
     END IF;
   END;

   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshl_stdar(arg1, arg2, '0', olen); END;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshr_stdar(arg1, arg2, '0', olen); END;
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshl_stdar(arg1, arg2, '0', olen); END;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshr_stdar(arg1, arg2, '0', olen); END;

   FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN fshl_stdar(arg1, arg2, arg1(arg1'LEFT), olen); END;
   FUNCTION fshr_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN fshr_stdar(arg1, arg2, arg1(arg1'LEFT), olen); END;
   FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN fshl_stdar(arg1, arg2, arg1(arg1'LEFT), olen); END;
   FUNCTION fshr_stdar(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN fshr_stdar(arg1, arg2, arg1(arg1'LEFT), olen); END;


   FUNCTION fshl(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
     VARIABLE temp: UNSIGNED(len-1 DOWNTO 0);
     --SUBTYPE  sw_range IS NATURAL range 1 TO len;
     VARIABLE sw: NATURAL range 1 TO len;
     VARIABLE temp_idx : INTEGER; --2.1.6.3
   BEGIN
     sw := 1;
     result := (others => sbit);
     result(ilen-1 DOWNTO 0) := arg1;
     FOR i IN arg2'reverse_range LOOP
       temp := (others => '0');
       FOR i2 IN len-1-sw DOWNTO 0 LOOP
         --was:temp(i2+sw) := result(i2);
         temp_idx := add_nat(i2,sw);
         temp(temp_idx) := result(i2);
       END LOOP;
       result := UNSIGNED(mux_v(STD_LOGIC_VECTOR(concat_uns(result,temp)), arg2(i)));
       sw := minimum(mult_natural(sw,2), len);
     END LOOP;
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshr(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
     VARIABLE temp: UNSIGNED(len-1 DOWNTO 0);
     SUBTYPE  sw_range IS NATURAL range 1 TO len;
     VARIABLE sw: sw_range;
     VARIABLE result_idx : INTEGER; --2.1.6.3
   BEGIN
     sw := 1;
     result := (others => sbit);
     result(ilen-1 DOWNTO 0) := arg1;
     FOR i IN arg2'reverse_range LOOP
       temp := (others => sbit);
       FOR i2 IN len-1-sw DOWNTO 0 LOOP
         -- was: temp(i2) := result(i2+sw);
         result_idx := add_nat(i2,sw);
         temp(i2) := result(result_idx);
       END LOOP;
       result := UNSIGNED(mux_v(STD_LOGIC_VECTOR(concat_uns(result,temp)), arg2(i)));
       sw := minimum(mult_natural(sw,2), len);
     END LOOP;
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshl(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT arg1l: NATURAL := arg1'LENGTH - 1;
     ALIAS    arg1x: UNSIGNED(arg1l DOWNTO 0) IS arg1;
     CONSTANT arg2l: NATURAL := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE arg1x_pad: UNSIGNED(arg1l+1 DOWNTO 0);
     VARIABLE result: UNSIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others=>'0');
     arg1x_pad(arg1l+1) := sbit;
     arg1x_pad(arg1l downto 0) := arg1x;
     IF arg2l = 0 THEN
       RETURN fshr(arg1x_pad, UNSIGNED(arg2x), sbit, olen);
     -- ELSIF arg1l = 0 THEN
     --   RETURN fshl(sbit & arg1x, arg2x, sbit, olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
       =>
         RETURN fshl(arg1x_pad, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);

       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
       =>
         RETURN fshr(arg1x_pad(arg1l+1 DOWNTO 1), not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);

       WHEN others =>
         --synopsys translate_off
         result := resolve_unsigned(
           fshl(arg1x_pad, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit,  olen),
           fshr(arg1x_pad(arg1l+1 DOWNTO 1), not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen)
         );
         --synopsys translate_on
         RETURN result;
       END CASE;
     END IF;
   END;

   FUNCTION fshr(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT arg2l: INTEGER := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE result: UNSIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others => '0');
     IF arg2l = 0 THEN
       RETURN fshl(arg1, UNSIGNED(arg2x), olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
       =>
         RETURN fshr(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);

       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
       =>
         RETURN fshl(arg1 & '0', not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_unsigned(
           fshr(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen),
           fshl(arg1 & '0', not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen)
         );
         --synopsys translate_on
	 return result;
       END CASE;
     END IF;
   END;

   FUNCTION fshl(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshl(arg1, arg2, '0', olen); END;
   FUNCTION fshr(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshr(arg1, arg2, '0', olen); END;
   FUNCTION fshl(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshl(arg1, arg2, '0', olen); END;
   FUNCTION fshr(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshr(arg1, arg2, '0', olen); END;

   FUNCTION fshl(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN SIGNED(fshl(UNSIGNED(arg1), arg2, arg1(arg1'LEFT), olen)); END;
   FUNCTION fshr(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN SIGNED(fshr(UNSIGNED(arg1), arg2, arg1(arg1'LEFT), olen)); END;
   FUNCTION fshl(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN SIGNED(fshl(UNSIGNED(arg1), arg2, arg1(arg1'LEFT), olen)); END;
   FUNCTION fshr(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN SIGNED(fshr(UNSIGNED(arg1), arg2, arg1(arg1'LEFT), olen)); END;


   FUNCTION frot(arg1: STD_LOGIC_VECTOR; arg2: STD_LOGIC_VECTOR; signd2: BOOLEAN; sdir: INTEGER range -1 TO 1) RETURN STD_LOGIC_VECTOR IS
     CONSTANT len: INTEGER := arg1'LENGTH;
     VARIABLE result: STD_LOGIC_VECTOR(len-1 DOWNTO 0);
     VARIABLE temp: STD_LOGIC_VECTOR(len-1 DOWNTO 0);
     SUBTYPE sw_range IS NATURAL range 0 TO len-1;
     VARIABLE sw: sw_range;
     VARIABLE temp_idx : INTEGER; --2.1.6.3
   BEGIN
     result := (others=>'0');
     result := arg1;
     sw := sdir MOD len;
     FOR i IN arg2'reverse_range LOOP
       EXIT WHEN sw = 0;
       IF signd2 AND i = arg2'LEFT THEN 
         sw := sub_int(len,sw); 
       END IF;
       -- temp := result(len-sw-1 DOWNTO 0) & result(len-1 DOWNTO len-sw)
       FOR i2 IN len-1 DOWNTO 0 LOOP
         --was: temp((i2+sw) MOD len) := result(i2);
         temp_idx := add_nat(i2,sw) MOD len;
         temp(temp_idx) := result(i2);
       END LOOP;
       result := mux_v(STD_LOGIC_VECTOR(concat_vect(result,temp)), arg2(i));
       sw := mod_natural(mult_natural(sw,2), len);
     END LOOP;
     RETURN result;
   END frot;

   FUNCTION frol(arg1: STD_LOGIC_VECTOR; arg2: UNSIGNED) RETURN STD_LOGIC_VECTOR IS
     BEGIN RETURN frot(arg1, STD_LOGIC_VECTOR(arg2), FALSE, 1); END;
   FUNCTION fror(arg1: STD_LOGIC_VECTOR; arg2: UNSIGNED) RETURN STD_LOGIC_VECTOR IS
     BEGIN RETURN frot(arg1, STD_LOGIC_VECTOR(arg2), FALSE, -1); END;
   FUNCTION frol(arg1: STD_LOGIC_VECTOR; arg2: SIGNED  ) RETURN STD_LOGIC_VECTOR IS
     BEGIN RETURN frot(arg1, STD_LOGIC_VECTOR(arg2), TRUE, 1); END;
   FUNCTION fror(arg1: STD_LOGIC_VECTOR; arg2: SIGNED  ) RETURN STD_LOGIC_VECTOR IS
     BEGIN RETURN frot(arg1, STD_LOGIC_VECTOR(arg2), TRUE, -1); END;

-----------------------------------------------------------------
-- indexing functions: LSB always has index 0
-----------------------------------------------------------------

   FUNCTION readindex(vec: STD_LOGIC_VECTOR; index: INTEGER                 ) RETURN STD_LOGIC IS
     CONSTANT len : INTEGER := vec'LENGTH;
     ALIAS    vec0: STD_LOGIC_VECTOR(len-1 DOWNTO 0) IS vec;
   BEGIN
     IF index >= len OR index < 0 THEN
       RETURN 'X';
     END IF;
     RETURN vec0(index);
   END;

   FUNCTION readslice(vec: STD_LOGIC_VECTOR; index: INTEGER; width: POSITIVE) RETURN STD_LOGIC_VECTOR IS
     CONSTANT len : INTEGER := vec'LENGTH;
     CONSTANT indexPwidthM1 : INTEGER := index+width-1; --2.1.6.3
     ALIAS    vec0: STD_LOGIC_VECTOR(len-1 DOWNTO 0) IS vec;
     CONSTANT xxx : STD_LOGIC_VECTOR(width-1 DOWNTO 0) := (others => 'X');
   BEGIN
     IF index+width > len OR index < 0 THEN
       RETURN xxx;
     END IF;
     RETURN vec0(indexPwidthM1 DOWNTO index);
   END;

   FUNCTION writeindex(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC       ; index: INTEGER) RETURN STD_LOGIC_VECTOR IS
     CONSTANT len : INTEGER := vec'LENGTH;
     VARIABLE vec0: STD_LOGIC_VECTOR(len-1 DOWNTO 0);
     CONSTANT xxx : STD_LOGIC_VECTOR(len-1 DOWNTO 0) := (others => 'X');
   BEGIN
     vec0 := vec;
     IF index >= len OR index < 0 THEN
       RETURN xxx;
     END IF;
     vec0(index) := dinput;
     RETURN vec0;
   END;

   FUNCTION n_bits(p: NATURAL) RETURN POSITIVE IS
     VARIABLE n_b : POSITIVE;
     VARIABLE p_v : NATURAL;
   BEGIN
     p_v := p;
     FOR i IN 1 TO 32 LOOP
       p_v := div_natural(p_v,2);
       n_b := i;
       EXIT WHEN (p_v = 0);
     END LOOP;
     RETURN n_b;
   END;


--   FUNCTION writeslice(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC_VECTOR; index: INTEGER) RETURN STD_LOGIC_VECTOR IS
--
--     CONSTANT vlen: INTEGER := vec'LENGTH;
--     CONSTANT ilen: INTEGER := dinput'LENGTH;
--     CONSTANT max_shift: INTEGER := vlen-ilen;
--     CONSTANT ones: UNSIGNED(ilen-1 DOWNTO 0) := (others => '1');
--     CONSTANT xxx : STD_LOGIC_VECTOR(vlen-1 DOWNTO 0) := (others => 'X');
--     VARIABLE shift : UNSIGNED(n_bits(max_shift)-1 DOWNTO 0);
--     VARIABLE vec0: STD_LOGIC_VECTOR(vlen-1 DOWNTO 0);
--     VARIABLE inp: UNSIGNED(vlen-1 DOWNTO 0);
--     VARIABLE mask: UNSIGNED(vlen-1 DOWNTO 0);
--   BEGIN
--     inp := (others => '0');
--     mask := (others => '0');
--
--     IF index > max_shift OR index < 0 THEN
--       RETURN xxx;
--     END IF;
--
--     shift := CONV_UNSIGNED(index, shift'LENGTH);
--     inp(ilen-1 DOWNTO 0) := UNSIGNED(dinput);
--     mask(ilen-1 DOWNTO 0) := ones;
--     inp := fshl(inp, shift, vlen);
--     mask := fshl(mask, shift, vlen);
--     vec0 := (vec and (not STD_LOGIC_VECTOR(mask))) or STD_LOGIC_VECTOR(inp);
--     RETURN vec0;
--   END;

   FUNCTION writeslice(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC_VECTOR; enable: STD_LOGIC_VECTOR; byte_width: INTEGER;  index: INTEGER) RETURN STD_LOGIC_VECTOR IS

     type enable_matrix is array (0 to enable'LENGTH-1 ) of std_logic_vector(byte_width-1 downto 0);
     CONSTANT vlen: INTEGER := vec'LENGTH;
     CONSTANT ilen: INTEGER := dinput'LENGTH;
     CONSTANT max_shift: INTEGER := vlen-ilen;
     CONSTANT ones: UNSIGNED(ilen-1 DOWNTO 0) := (others => '1');
     CONSTANT xxx : STD_LOGIC_VECTOR(vlen-1 DOWNTO 0) := (others => 'X');
     VARIABLE shift : UNSIGNED(n_bits(max_shift)-1 DOWNTO 0);
     VARIABLE vec0: STD_LOGIC_VECTOR(vlen-1 DOWNTO 0);
     VARIABLE inp: UNSIGNED(vlen-1 DOWNTO 0);
     VARIABLE mask: UNSIGNED(vlen-1 DOWNTO 0);
     VARIABLE mask2: UNSIGNED(vlen-1 DOWNTO 0);
     VARIABLE enables: enable_matrix;
     VARIABLE cat_enables: STD_LOGIC_VECTOR(ilen-1 DOWNTO 0 );
     VARIABLE lsbi : INTEGER;
     VARIABLE msbi : INTEGER;

   BEGIN
     cat_enables := (others => '0');
     lsbi := 0;
     msbi := byte_width-1;
     inp := (others => '0');
     mask := (others => '0');

     IF index > max_shift OR index < 0 THEN
       RETURN xxx;
     END IF;

     --initialize enables
     for i in 0 TO (enable'LENGTH-1) loop
       enables(i)  := (others => enable(i));
       cat_enables(msbi downto lsbi) := enables(i) ;
       lsbi := msbi+1;
       msbi := msbi+byte_width;
     end loop;


     shift := CONV_UNSIGNED(index, shift'LENGTH);
     inp(ilen-1 DOWNTO 0) := UNSIGNED(dinput);
     mask(ilen-1 DOWNTO 0) := UNSIGNED((STD_LOGIC_VECTOR(ones) AND cat_enables));
     inp := fshl(inp, shift, vlen);
     mask := fshl(mask, shift, vlen);
     vec0 := (vec and (not STD_LOGIC_VECTOR(mask))) or STD_LOGIC_VECTOR(inp);
     RETURN vec0;
   END;


   FUNCTION ceil_log2(size : NATURAL) return NATURAL is
     VARIABLE cnt : NATURAL;
     VARIABLE res : NATURAL;
   begin
     cnt := 1;
     res := 0;
     while (cnt < size) loop
       res := res + 1;
       cnt := 2 * cnt;
     end loop;
     return res;
   END;
   
   FUNCTION bits(size : NATURAL) return NATURAL is
   begin
     return ceil_log2(size);
   END;

   PROCEDURE csa(a, b, c: IN INTEGER; s, cout: OUT STD_LOGIC_VECTOR) IS
   BEGIN
     s    := conv_std_logic_vector(a, s'LENGTH) xor conv_std_logic_vector(b, s'LENGTH) xor conv_std_logic_vector(c, s'LENGTH);
     cout := ( (conv_std_logic_vector(a, cout'LENGTH) and conv_std_logic_vector(b, cout'LENGTH)) or (conv_std_logic_vector(a, cout'LENGTH) and conv_std_logic_vector(c, cout'LENGTH)) or (conv_std_logic_vector(b, cout'LENGTH) and conv_std_logic_vector(c, cout'LENGTH)) );
   END PROCEDURE csa;

   PROCEDURE csha(a, b: IN INTEGER; s, cout: OUT STD_LOGIC_VECTOR) IS
   BEGIN
     s    := conv_std_logic_vector(a, s'LENGTH) xor conv_std_logic_vector(b, s'LENGTH);
     cout := (conv_std_logic_vector(a, cout'LENGTH) and conv_std_logic_vector(b, cout'LENGTH));
   END PROCEDURE csha;

END funcs;

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_comps.vhd 
LIBRARY ieee;

USE ieee.std_logic_1164.all;

PACKAGE mgc_comps IS
 
FUNCTION ifeqsel(arg1, arg2, seleq, selne : INTEGER) RETURN INTEGER;
FUNCTION ceil_log2(size : NATURAL) return NATURAL;
 

COMPONENT mgc_not
  GENERIC (
    width  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    z: out std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_and
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_nand
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_or
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_nor
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_xor
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_xnor
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mux
  GENERIC (
    width  :  NATURAL;
    ctrlw  :  NATURAL;
    p2ctrlw : NATURAL := 0
  );
  PORT (
    a: in  std_logic_vector(width*(2**ctrlw) - 1 DOWNTO 0);
    c: in  std_logic_vector(ctrlw            - 1 DOWNTO 0);
    z: out std_logic_vector(width            - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mux1hot
  GENERIC (
    width  : NATURAL;
    ctrlw  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ctrlw - 1 DOWNTO 0);
    c: in  std_logic_vector(ctrlw       - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_reg_pos
  GENERIC (
    width  : NATURAL;
    has_a_rst : NATURAL;  -- 0 to 1
    a_rst_on  : NATURAL;  -- 0 to 1
    has_s_rst : NATURAL;  -- 0 to 1
    s_rst_on  : NATURAL;  -- 0 to 1
    has_enable : NATURAL; -- 0 to 1
    enable_on  : NATURAL  -- 0 to 1
  );
  PORT (
    clk: in  std_logic;
    d  : in  std_logic_vector(width-1 DOWNTO 0);
    z  : out std_logic_vector(width-1 DOWNTO 0);
    sync_rst_val : in std_logic_vector(width-1 DOWNTO 0);
    sync_rst : in std_logic;
    async_rst_val : in std_logic_vector(width-1 DOWNTO 0);
    async_rst : in std_logic;
    en : in std_logic
  );
END COMPONENT;

COMPONENT mgc_reg_neg
  GENERIC (
    width  : NATURAL;
    has_a_rst : NATURAL;  -- 0 to 1
    a_rst_on  : NATURAL;  -- 0 to 1
    has_s_rst : NATURAL;  -- 0 to 1
    s_rst_on  : NATURAL;   -- 0 to 1
    has_enable : NATURAL; -- 0 to 1
    enable_on  : NATURAL -- 0 to 1
  );
  PORT (
    clk: in  std_logic;
    d  : in  std_logic_vector(width-1 DOWNTO 0);
    z  : out std_logic_vector(width-1 DOWNTO 0);
    sync_rst_val : in std_logic_vector(width-1 DOWNTO 0);
    sync_rst : in std_logic;
    async_rst_val : in std_logic_vector(width-1 DOWNTO 0);
    async_rst : in std_logic;
    en : in std_logic
  );
END COMPONENT;

COMPONENT mgc_generic_reg
  GENERIC(
   width: natural := 8;
   ph_clk: integer range 0 to 1 := 1; -- clock polarity, 1=rising_edge
   ph_en: integer range 0 to 1 := 1;
   ph_a_rst: integer range 0 to 1 := 1;   --  0 to 1 IGNORED
   ph_s_rst: integer range 0 to 1 := 1;   --  0 to 1 IGNORED
   a_rst_used: integer range 0 to 1 := 1;
   s_rst_used: integer range 0 to 1 := 0;
   en_used: integer range 0 to 1 := 1
  );
  PORT(
   d: std_logic_vector(width-1 downto 0);
   clk: in std_logic;
   en: in std_logic;
   a_rst: in std_logic;
   s_rst: in std_logic;
   q: out std_logic_vector(width-1 downto 0)
  );
END COMPONENT;

COMPONENT mgc_equal
  GENERIC (
    width  : NATURAL
  );
  PORT (
    a : in  std_logic_vector(width-1 DOWNTO 0);
    b : in  std_logic_vector(width-1 DOWNTO 0);
    eq: out std_logic;
    ne: out std_logic
  );
END COMPONENT;

COMPONENT mgc_shift_l
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_r
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_bl
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_br
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_rot
  GENERIC (
    width  : NATURAL;
    width_s: NATURAL;
    signd_s: NATURAL;      -- 0:unsigned 1:signed
    sleft  : NATURAL;      -- 0:right 1:left;
    log2w  : NATURAL := 0; -- LOG2(width)
    l2wp2  : NATURAL := 0  --2**LOG2(width)
  );
  PORT (
    a : in  std_logic_vector(width  -1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width  -1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_add
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_sub
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_add_ci
  GENERIC (
    width_a : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width_a, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width_a, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width_a,width_b)-1 DOWNTO 0);
    c: in  std_logic_vector(0 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width_a,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_addc
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    c: in  std_logic_vector(0 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_add3
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_c : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_c : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    c: in  std_logic_vector(ifeqsel(width_c,0,width,width_c)-1 DOWNTO 0);
    d: in  std_logic_vector(0 DOWNTO 0);
    e: in  std_logic_vector(0 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_add_pipe
  GENERIC (
     width_a : natural := 16;
     signd_a : integer range 0 to 1 := 0;
     width_b : natural := 3;
     signd_b : integer range 0 to 1 := 0;
     width_z : natural := 18;
     ph_clk : integer range 0 to 1 := 1;
     ph_en : integer range 0 to 1 := 1;
     ph_a_rst : integer range 0 to 1 := 1;
     ph_s_rst : integer range 0 to 1 := 1;
     n_outreg : natural := 2;
     stages : natural := 2; -- Default value is minimum required value
     a_rst_used: integer range 0 to 1 := 1;
     s_rst_used: integer range 0 to 1 := 0;
     en_used: integer range 0 to 1 := 1
     );
  PORT(
     a: in std_logic_vector(width_a-1 downto 0);
     b: in std_logic_vector(width_b-1 downto 0);
     clk: in std_logic;
     en: in std_logic;
     a_rst: in std_logic;
     s_rst: in std_logic;
     z: out std_logic_vector(width_z-1 downto 0)
     );
END COMPONENT;

COMPONENT mgc_sub_pipe
  GENERIC (
     width_a : natural := 16;
     signd_a : integer range 0 to 1 := 0;
     width_b : natural := 3;
     signd_b : integer range 0 to 1 := 0;
     width_z : natural := 18;
     ph_clk : integer range 0 to 1 := 1;
     ph_en : integer range 0 to 1 := 1;
     ph_a_rst : integer range 0 to 1 := 1;
     ph_s_rst : integer range 0 to 1 := 1;
     n_outreg : natural := 2;
     stages : natural := 2; -- Default value is minimum required value
     a_rst_used: integer range 0 to 1 := 1;
     s_rst_used: integer range 0 to 1 := 0;
     en_used: integer range 0 to 1 := 1
     );
  PORT(
     a: in std_logic_vector(width_a-1 downto 0);
     b: in std_logic_vector(width_b-1 downto 0);
     clk: in std_logic;
     en: in std_logic;
     a_rst: in std_logic;
     s_rst: in std_logic;
     z: out std_logic_vector(width_z-1 downto 0)
     );
END COMPONENT;

COMPONENT mgc_addc_pipe
  GENERIC (
     width_a : natural := 16;
     signd_a : integer range 0 to 1 := 0;
     width_b : natural := 3;
     signd_b : integer range 0 to 1 := 0;
     width_z : natural := 18;
     ph_clk : integer range 0 to 1 := 1;
     ph_en : integer range 0 to 1 := 1;
     ph_a_rst : integer range 0 to 1 := 1;
     ph_s_rst : integer range 0 to 1 := 1;
     n_outreg : natural := 2;
     stages : natural := 2; -- Default value is minimum required value
     a_rst_used: integer range 0 to 1 := 1;
     s_rst_used: integer range 0 to 1 := 0;
     en_used: integer range 0 to 1 := 1
     );
  PORT(
     a: in std_logic_vector(width_a-1 downto 0);
     b: in std_logic_vector(width_b-1 downto 0);
     c: in std_logic_vector(0 downto 0);
     clk: in std_logic;
     en: in std_logic;
     a_rst: in std_logic;
     s_rst: in std_logic;
     z: out std_logic_vector(width_z-1 downto 0)
     );
END COMPONENT;

COMPONENT mgc_addsub
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    add: in  std_logic;
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_accu
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps-1 DOWNTO 0);
    z: out std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_abs
  GENERIC (
    width  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    z: out std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_z : NATURAL    -- <= width_a + width_b
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul_fast
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_z : NATURAL    -- <= width_a + width_b
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul_pipe
  GENERIC (
    width_a       : NATURAL;
    signd_a       : NATURAL;
    width_b       : NATURAL;
    signd_b       : NATURAL;
    width_z       : NATURAL; -- <= width_a + width_b
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 

  );
  PORT (
    a     : in  std_logic_vector(width_a-1 DOWNTO 0);
    b     : in  std_logic_vector(width_b-1 DOWNTO 0);
    clk   : in  std_logic;
    en    : in  std_logic;
    a_rst : in  std_logic;
    s_rst : in  std_logic;
    z     : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul2add1
  GENERIC (
    gentype : NATURAL;
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_b2 : NATURAL;
    signd_b2 : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_d2 : NATURAL;
    signd_d2 : NATURAL;
    width_e : NATURAL;
    signd_e : NATURAL;
    width_z : NATURAL;   -- <= max(width_a + width_b, width_c + width_d)+1
    isadd   : NATURAL;
    add_b2  : NATURAL;
    add_d2  : NATURAL
  );
  PORT (
    a   : in  std_logic_vector(width_a-1 DOWNTO 0);
    b   : in  std_logic_vector(width_b-1 DOWNTO 0);
    b2  : in  std_logic_vector(width_b2-1 DOWNTO 0);
    c   : in  std_logic_vector(width_c-1 DOWNTO 0);
    d   : in  std_logic_vector(width_d-1 DOWNTO 0);
    d2  : in  std_logic_vector(width_d2-1 DOWNTO 0);
    cst : in  std_logic_vector(width_e-1 DOWNTO 0);
    z   : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul2add1_pipe
  GENERIC (
    gentype : NATURAL;
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_b2 : NATURAL;
    signd_b2 : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_d2 : NATURAL;
    signd_d2 : NATURAL;
    width_e : NATURAL;
    signd_e : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c + width_d)+1
    isadd   : NATURAL;
    add_b2   : NATURAL;
    add_d2   : NATURAL;
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 
  );
  PORT (
    a     : in  std_logic_vector(width_a-1 DOWNTO 0);
    b     : in  std_logic_vector(width_b-1 DOWNTO 0);
    b2     : in  std_logic_vector(width_b2-1 DOWNTO 0);
    c     : in  std_logic_vector(width_c-1 DOWNTO 0);
    d     : in  std_logic_vector(width_d-1 DOWNTO 0);
    d2     : in  std_logic_vector(width_d2-1 DOWNTO 0);
    cst   : in  std_logic_vector(width_e-1 DOWNTO 0);
    clk   : in  std_logic;
    en    : in  std_logic;
    a_rst : in  std_logic;
    s_rst : in  std_logic;
    z     : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_muladd1
  -- operation is z = a * (b + d) + c + cst
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_cst : NATURAL;
    signd_cst : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c, width_cst)+1
    add_axb : NATURAL;
    add_c   : NATURAL;
    add_d   : NATURAL
  );
  PORT (
    a:   in  std_logic_vector(width_a-1 DOWNTO 0);
    b:   in  std_logic_vector(width_b-1 DOWNTO 0);
    c:   in  std_logic_vector(width_c-1 DOWNTO 0);
    cst: in  std_logic_vector(width_cst-1 DOWNTO 0);
    d:   in  std_logic_vector(width_d-1 DOWNTO 0);
    z:   out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_muladd1_pipe
  -- operation is z = a * (b + d) + c + cst
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_cst : NATURAL;
    signd_cst : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c, width_cst)+1
    add_axb : NATURAL;
    add_c   : NATURAL;
    add_d   : NATURAL;
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 
  );
  PORT (
    a     : in  std_logic_vector(width_a-1 DOWNTO 0);
    b     : in  std_logic_vector(width_b-1 DOWNTO 0);
    c     : in  std_logic_vector(width_c-1 DOWNTO 0);
    cst   : in  std_logic_vector(width_cst-1 DOWNTO 0);
    d     : in  std_logic_vector(width_d-1 DOWNTO 0);
    clk   : in  std_logic;
    en    : in  std_logic;
    a_rst : in  std_logic;
    s_rst : in  std_logic;
    z     : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mulacc_pipe
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c)+1
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 
  );
  PORT (
    a         : in  std_logic_vector(width_a-1 DOWNTO 0);
    b         : in  std_logic_vector(width_b-1 DOWNTO 0);
    c         : in  std_logic_vector(width_c-1 DOWNTO 0);
    load      : in  std_logic;
    datavalid : in  std_logic;
    clk       : in  std_logic;
    en        : in  std_logic;
    a_rst     : in  std_logic;
    s_rst     : in  std_logic;
    z         : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul2acc_pipe
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_e : NATURAL;
    signd_e : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c)+1
    add_cxd : NATURAL;
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 
  );
  PORT (
    a         : in  std_logic_vector(width_a-1 DOWNTO 0);
    b         : in  std_logic_vector(width_b-1 DOWNTO 0);
    c         : in  std_logic_vector(width_c-1 DOWNTO 0);
    d         : in  std_logic_vector(width_d-1 DOWNTO 0);
    e         : in  std_logic_vector(width_e-1 DOWNTO 0);
    load      : in  std_logic;
    datavalid : in  std_logic;
    clk       : in  std_logic;
    en        : in  std_logic;
    a_rst     : in  std_logic;
    s_rst     : in  std_logic;
    z         : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_div
  GENERIC (
    width_a : NATURAL;
    width_b : NATURAL;
    signd   : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_a-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mod
  GENERIC (
    width_a : NATURAL;
    width_b : NATURAL;
    signd   : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_b-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_rem
  GENERIC (
    width_a : NATURAL;
    width_b : NATURAL;
    signd   : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_b-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_csa
  GENERIC (
     width : NATURAL
  );
  PORT (
     a: in std_logic_vector(width-1 downto 0);
     b: in std_logic_vector(width-1 downto 0);
     c: in std_logic_vector(width-1 downto 0);
     s: out std_logic_vector(width-1 downto 0);
     cout: out std_logic_vector(width-1 downto 0)
  );
END COMPONENT;

COMPONENT mgc_csha
  GENERIC (
     width : NATURAL
  );
  PORT (
     a: in std_logic_vector(width-1 downto 0);
     b: in std_logic_vector(width-1 downto 0);
     s: out std_logic_vector(width-1 downto 0);
     cout: out std_logic_vector(width-1 downto 0)
  );
END COMPONENT;

COMPONENT mgc_rom
    GENERIC (
      rom_id : natural := 1;
      size : natural := 33;
      width : natural := 32
      );
    PORT (
      data_in : std_logic_vector((size*width)-1 downto 0);
      addr : std_logic_vector(ceil_log2(size)-1 downto 0);
      data_out : out std_logic_vector(width-1 downto 0)
    );
END COMPONENT;

END mgc_comps;

PACKAGE BODY mgc_comps IS
 
   FUNCTION ceil_log2(size : NATURAL) return NATURAL is
     VARIABLE cnt : NATURAL;
     VARIABLE res : NATURAL;
   begin
     cnt := 1;
     res := 0;
     while (cnt < size) loop
       res := res + 1;
       cnt := 2 * cnt;
     end loop;
     return res;
   END;

   FUNCTION ifeqsel(arg1, arg2, seleq, selne : INTEGER) RETURN INTEGER IS
   BEGIN
     IF(arg1 = arg2) THEN
       RETURN(seleq) ;
     ELSE
       RETURN(selne) ;
     END IF;
   END;
 
END mgc_comps;

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_mul_pipe_beh.vhd 

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY mgc_mul_pipe IS
  GENERIC (
    width_a       : NATURAL;
    signd_a       : NATURAL;
    width_b       : NATURAL;
    signd_b       : NATURAL;
    width_z       : NATURAL; -- <= width_a + width_b
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 

  );
  PORT (
    a     : in  std_logic_vector(width_a-1 DOWNTO 0);
    b     : in  std_logic_vector(width_b-1 DOWNTO 0);
    clk   : in  std_logic;
    en    : in  std_logic;
    a_rst : in  std_logic;
    s_rst : in  std_logic;
    z     : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END mgc_mul_pipe;

LIBRARY IEEE;

USE ieee.std_logic_arith.all;

ARCHITECTURE beh OF mgc_mul_pipe IS
  TYPE reg_array_type is array(natural range<>) of std_logic_vector(width_z-1 DOWNTO 0); 
  SIGNAL xz : std_logic_vector(width_a+width_b DOWNTO 0);

--MF Added pipelined input
    signal a_f     : STD_LOGIC_VECTOR(width_a-1 downto 0); 
    signal b_f     : STD_LOGIC_VECTOR(width_b-1 downto 0);
   type a_array is array (natural range <>) of STD_LOGIC_VECTOR(width_a-1 downto 0);
   type b_array is array (natural range <>) of STD_LOGIC_VECTOR(width_b-1 downto 0);
BEGIN
  n_inreg_gt_0: if n_inreg > 0 generate
    GENPOS_INREG: IF clock_edge = 1 GENERATE
     I0: process(clk)
        variable a_in_reg: a_array(n_inreg-1 downto 0);
        variable b_in_reg: b_array(n_inreg-1 downto 0);
      begin
        if (clk'event and clk = '1' ) then
          if (conv_integer(en) = enable_active) then
            for i in n_inreg - 2 downto 0 loop
              a_in_reg(i+1) := a_in_reg(i);
              b_in_reg(i+1) := b_in_reg(i);
            end loop;                                                                                                                             
            a_in_reg(0) := a;
            b_in_reg(0) := b;

            a_f <= a_in_reg(n_inreg-1);             
            b_f <= b_in_reg(n_inreg-1);    
                                                   
          end if;
        end if;
      end process;
    END GENERATE;
  
   GENNEG_INREG: IF clock_edge = 0 GENERATE
     I0: process(clk)
        variable a_in_reg: a_array(n_inreg-1 downto 0);
        variable b_in_reg: b_array(n_inreg-1 downto 0);
      begin
        if (clk'event and clk = '0' ) then
          if (conv_integer(en) = enable_active) then
            for i in n_inreg - 2 downto 0 loop
              a_in_reg(i+1) := a_in_reg(i);
              b_in_reg(i+1) := b_in_reg(i);
            end loop;                                                                                                                             
            a_in_reg(0) := a;
            b_in_reg(0) := b;            
                                 
            a_f <= a_in_reg(n_inreg-1);             
            b_f <= b_in_reg(n_inreg-1);
                                                        
          end if;
        end if;
      end process;
    END GENERATE;
  END GENERATE;

  n_inreg_eq_0: if n_inreg = 0 generate
    a_f <= a;
    b_f <= b;
  end generate n_inreg_eq_0;

  xz <= '0'&(unsigned(a_f) * unsigned(b_f)) WHEN signd_a = 0 AND signd_b = 0 ELSE
            (  signed(a_f) * unsigned(b_f)) WHEN signd_a = 1 AND signd_b = 0 ELSE
            (unsigned(a_f) *   signed(b_f)) WHEN signd_a = 0 AND signd_b = 1 ELSE
        '0'&(  signed(a_f) *   signed(b_f));

  GENPOS: IF clock_edge = 1 GENERATE
    PROCESS (clk)
    VARIABLE reg_array: reg_array_type(stages-2 DOWNTO 0);
    BEGIN
      IF ( clk'EVENT AND clk = '1') THEN
        IF ( conv_integer(en) = enable_active) THEN
          FOR I IN stages-2 DOWNTO 1 LOOP
            reg_array(I) := reg_array(I-1);
          END LOOP;
          reg_array(0) := xz(width_z-1 DOWNTO 0);
          z <= reg_array(stages-2);
        END IF;
      END IF;
    END PROCESS;
  END GENERATE;

  GENNEG: IF clock_edge = 0 GENERATE
    PROCESS (clk)
    VARIABLE reg_array: reg_array_type(stages-2 DOWNTO 0);
    BEGIN
      IF ( clk'EVENT AND clk = '0') THEN
        IF ( conv_integer(en) = enable_active) THEN
          FOR I IN stages-2 DOWNTO 1 LOOP
            reg_array(I) := reg_array(I-1);
          END LOOP;
          reg_array(0) := xz(width_z-1 DOWNTO 0);
          z <= reg_array(stages-2);
        END IF;
      END IF;
    END PROCESS;
  END GENERATE;
END beh;

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_shift_comps_v5.vhd 
LIBRARY ieee;

USE ieee.std_logic_1164.all;

PACKAGE mgc_shift_comps_v5 IS

COMPONENT mgc_shift_l_v5
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_r_v5
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_bl_v5
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_br_v5
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

END mgc_shift_comps_v5;

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_shift_bl_beh_v5.vhd 
LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY mgc_shift_bl_v5 IS
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END mgc_shift_bl_v5;

LIBRARY ieee;

USE ieee.std_logic_arith.all;

ARCHITECTURE beh OF mgc_shift_bl_v5 IS

  FUNCTION resolve_std_logic_vector(input1: STD_LOGIC_VECTOR; input2: STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR IS
    CONSTANT len: INTEGER := input1'LENGTH;
    ALIAS input1a: STD_LOGIC_VECTOR(len-1 DOWNTO 0) IS input1;
    ALIAS input2a: STD_LOGIC_VECTOR(len-1 DOWNTO 0) IS input2;
    VARIABLE result: STD_LOGIC_VECTOR(len-1 DOWNTO 0);
  BEGIN
    result := (others => '0');
    --synopsys translate_off
    FOR i IN len-1 DOWNTO 0 LOOP
      result(i) := resolved(input1a(i) & input2a(i));
    END LOOP;
    --synopsys translate_on
    RETURN result;
  END;

  FUNCTION resolve_unsigned(input1: UNSIGNED; input2: UNSIGNED)
  RETURN UNSIGNED IS
  BEGIN
    RETURN UNSIGNED(resolve_std_logic_vector(STD_LOGIC_VECTOR(input1),
                                             STD_LOGIC_VECTOR(input2)));
  END;

  FUNCTION resolve_signed(input1: SIGNED; input2: SIGNED)
  RETURN SIGNED IS
  BEGIN
    RETURN SIGNED(resolve_std_logic_vector(STD_LOGIC_VECTOR(input1),
                                           STD_LOGIC_VECTOR(input2)));
  END;

  FUNCTION "not"(arg1: UNSIGNED) RETURN UNSIGNED IS
    BEGIN RETURN UNSIGNED(not STD_LOGIC_VECTOR(arg1)); END;

  FUNCTION maximum (arg1,arg2: INTEGER) RETURN INTEGER IS
  BEGIN
    IF(arg1 > arg2) THEN
      RETURN(arg1) ;
    ELSE
      RETURN(arg2) ;
    END IF;
  END;

  FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
    CONSTANT ilen: INTEGER := arg1'LENGTH;
    CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
    CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
    CONSTANT len: INTEGER := maximum(ilen, olen);
    VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
  BEGIN
    result := (others => sbit);
    result(ilenub DOWNTO 0) := arg1;
    result := shl(result, arg2);
    RETURN result(olenM1 DOWNTO 0);
  END;

  FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
    CONSTANT ilen: INTEGER := arg1'LENGTH;
    CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
    CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
    CONSTANT len: INTEGER := maximum(ilen, olen);
    VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
  BEGIN
    result := (others => sbit);
    result(ilenub DOWNTO 0) := arg1;
    result := shr(result, arg2);
    RETURN result(olenM1 DOWNTO 0);
  END;

  FUNCTION fshl_stdar(arg1: SIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
    CONSTANT ilen: INTEGER := arg1'LENGTH;
    CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
    CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
    CONSTANT len: INTEGER := maximum(ilen, olen);
    VARIABLE result: SIGNED(len-1 DOWNTO 0);
  BEGIN
    result := (others => sbit);
    result(ilenub DOWNTO 0) := arg1;
    result := shl(SIGNED(result), arg2);
    RETURN result(olenM1 DOWNTO 0);
  END;

  FUNCTION fshr_stdar(arg1: SIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
    CONSTANT ilen: INTEGER := arg1'LENGTH;
    CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
    CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
    CONSTANT len: INTEGER := maximum(ilen, olen);
    VARIABLE result: SIGNED(len-1 DOWNTO 0);
  BEGIN
    result := (others => sbit);
    result(ilenub DOWNTO 0) := arg1;
    result := shr(result, arg2);
    RETURN result(olenM1 DOWNTO 0);
  END;

 FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
    CONSTANT arg1l: NATURAL := arg1'LENGTH - 1;
    ALIAS    arg1x: UNSIGNED(arg1l DOWNTO 0) IS arg1;
    CONSTANT arg2l: NATURAL := arg2'LENGTH - 1;
    ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
    VARIABLE arg1x_pad: UNSIGNED(arg1l+1 DOWNTO 0);
    VARIABLE result: UNSIGNED(olen-1 DOWNTO 0);
  BEGIN
    result := (others=>'0');
    arg1x_pad(arg1l+1) := sbit;
    arg1x_pad(arg1l downto 0) := arg1x;
    IF arg2l = 0 THEN
      RETURN fshr_stdar(arg1x_pad, UNSIGNED(arg2x), sbit, olen);
    -- ELSIF arg1l = 0 THEN
    --   RETURN fshl(sbit & arg1x, arg2x, sbit, olen);
    ELSE
      CASE arg2x(arg2l) IS
      WHEN '0'
    --synopsys translate_off
           | 'L'
    --synopsys translate_on
      =>
        RETURN fshl_stdar(arg1x_pad, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
      WHEN '1'
    --synopsys translate_off
           | 'H'
    --synopsys translate_on
      =>
        RETURN fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
      WHEN others =>
        --synopsys translate_off
        result := resolve_unsigned(
          fshl_stdar(arg1x, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit,  olen),
          fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen)
        );
        --synopsys translate_on
        RETURN result;
      END CASE;
    END IF;
  END;

  FUNCTION fshl_stdar(arg1: SIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
    CONSTANT arg1l: NATURAL := arg1'LENGTH - 1;
    ALIAS    arg1x: SIGNED(arg1l DOWNTO 0) IS arg1;
    CONSTANT arg2l: NATURAL := arg2'LENGTH - 1;
    ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
    VARIABLE arg1x_pad: SIGNED(arg1l+1 DOWNTO 0);
    VARIABLE result: SIGNED(olen-1 DOWNTO 0);
  BEGIN
    result := (others=>'0');
    arg1x_pad(arg1l+1) := sbit;
    arg1x_pad(arg1l downto 0) := arg1x;
    IF arg2l = 0 THEN
      RETURN fshr_stdar(arg1x_pad, UNSIGNED(arg2x), sbit, olen);
    -- ELSIF arg1l = 0 THEN
    --   RETURN fshl(sbit & arg1x, arg2x, sbit, olen);
    ELSE
      CASE arg2x(arg2l) IS
      WHEN '0'
      --synopsys translate_off
           | 'L'
      --synopsys translate_on
      =>
        RETURN fshl_stdar(arg1x_pad, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
      WHEN '1'
      --synopsys translate_off
           | 'H'
      --synopsys translate_on
      =>
        RETURN fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
      WHEN others =>
        --synopsys translate_off
        result := resolve_signed(
          fshl_stdar(arg1x, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit,  olen),
          fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen)
        );
        --synopsys translate_on
        RETURN result;
      END CASE;
    END IF;
  END;

  FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE)
  RETURN UNSIGNED IS
  BEGIN
    RETURN fshl_stdar(arg1, arg2, '0', olen);
  END;

  FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE)
  RETURN SIGNED IS
  BEGIN
    RETURN fshl_stdar(arg1, arg2, arg1(arg1'LEFT), olen);
  END;

BEGIN
UNSGNED:  IF signd_a = 0 GENERATE
    z <= std_logic_vector(fshl_stdar(unsigned(a), signed(s), width_z));
  END GENERATE;
SGNED:  IF signd_a /= 0 GENERATE
    z <= std_logic_vector(fshl_stdar(  signed(a), signed(s), width_z));
  END GENERATE;
END beh;

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_shift_l_beh_v5.vhd 
LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY mgc_shift_l_v5 IS
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END mgc_shift_l_v5;

LIBRARY ieee;

USE ieee.std_logic_arith.all;

ARCHITECTURE beh OF mgc_shift_l_v5 IS

  FUNCTION maximum (arg1,arg2: INTEGER) RETURN INTEGER IS
  BEGIN
    IF(arg1 > arg2) THEN
      RETURN(arg1) ;
    ELSE
      RETURN(arg2) ;
    END IF;
  END;

  FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
    CONSTANT ilen: INTEGER := arg1'LENGTH;
    CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
    CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
    CONSTANT len: INTEGER := maximum(ilen, olen);
    VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
  BEGIN
    result := (others => sbit);
    result(ilenub DOWNTO 0) := arg1;
    result := shl(result, arg2);
    RETURN result(olenM1 DOWNTO 0);
  END;

  FUNCTION fshl_stdar(arg1: SIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
    CONSTANT ilen: INTEGER := arg1'LENGTH;
    CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
    CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
    CONSTANT len: INTEGER := maximum(ilen, olen);
    VARIABLE result: SIGNED(len-1 DOWNTO 0);
  BEGIN
    result := (others => sbit);
    result(ilenub DOWNTO 0) := arg1;
    result := shl(SIGNED(result), arg2);
    RETURN result(olenM1 DOWNTO 0);
  END;

  FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE)
  RETURN UNSIGNED IS
  BEGIN
    RETURN fshl_stdar(arg1, arg2, '0', olen);
  END;

  FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE)
  RETURN SIGNED IS
  BEGIN
    RETURN fshl_stdar(arg1, arg2, arg1(arg1'LEFT), olen);
  END;

BEGIN
UNSGNED:  IF signd_a = 0 GENERATE
    z <= std_logic_vector(fshl_stdar(unsigned(a), unsigned(s), width_z));
  END GENERATE;
SGNED:  IF signd_a /= 0 GENERATE
    z <= std_logic_vector(fshl_stdar(  signed(a), unsigned(s), width_z));
  END GENERATE;
END beh;

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/ccs_xilinx/hdl/BLOCK_1R1W_RBW_DUAL.vhd 
-- Memory Type:            BLOCK
-- Operating Mode:         Simple Dual Port (2-Port)
-- Clock Mode:             Dual Clock
-- 
-- RTL Code RW Resolution: RBW
-- Catapult RW Resolution: RBW
-- 
-- HDL Work Library:       Xilinx_RAMS_lib
-- Component Name:         BLOCK_1R1W_RBW_DUAL
-- Latency = 1:            RAM with no registers on inputs or outputs
--         = 2:            adds embedded register on RAM output
--         = 3:            adds fabric registers to non-clock input RAM pins
--         = 4:            adds fabric register to output (driven by embedded register from latency=2)

LIBRARY ieee;

  USE ieee.std_logic_1164.all;
  USE ieee.numeric_std.all;
PACKAGE BLOCK_1R1W_RBW_DUAL_pkg IS
  COMPONENT BLOCK_1R1W_RBW_DUAL IS
  GENERIC (
    addr_width : integer := 8 ;
    data_width : integer := 7 ;
    depth : integer := 256 ;
    latency : integer := 1 
    
  );
  PORT (
    clkr : in std_logic ;
    clkr_en : in std_logic ;
    clkw : in std_logic ;
    clkw_en : in std_logic ;
    d : in std_logic_vector(data_width-1 downto 0) ;
    q : out std_logic_vector(data_width-1 downto 0) ;
    radr : in std_logic_vector(addr_width-1 downto 0) ;
    wadr : in std_logic_vector(addr_width-1 downto 0) ;
    we : in std_logic 
    
  );
  END COMPONENT;
END BLOCK_1R1W_RBW_DUAL_pkg;
LIBRARY ieee;

  USE ieee.std_logic_1164.all;
  USE ieee.numeric_std.all;
ENTITY BLOCK_1R1W_RBW_DUAL IS
  GENERIC (
    addr_width : integer := 8 ;
    data_width : integer := 7 ;
    depth : integer := 256 ;
    latency : integer := 1 
    
  );
  PORT (
    clkr : in std_logic ;
    clkr_en : in std_logic ;
    clkw : in std_logic ;
    clkw_en : in std_logic ;
    d : in std_logic_vector(data_width-1 downto 0) ;
    q : out std_logic_vector(data_width-1 downto 0) ;
    radr : in std_logic_vector(addr_width-1 downto 0) ;
    wadr : in std_logic_vector(addr_width-1 downto 0) ;
    we : in std_logic 
    
  );
 END BLOCK_1R1W_RBW_DUAL;
ARCHITECTURE rtl OF BLOCK_1R1W_RBW_DUAL IS
  TYPE ram_t IS ARRAY (depth-1 DOWNTO 0) OF std_logic_vector(data_width-1 DOWNTO 0);
  SIGNAL mem : ram_t := (OTHERS => (OTHERS => '0'));
  ATTRIBUTE ram_style: STRING;
  ATTRIBUTE ram_style OF mem : SIGNAL IS "block";
  ATTRIBUTE syn_ramstyle: STRING;
  ATTRIBUTE syn_ramstyle OF mem : SIGNAL IS "block";
  
  SIGNAL ramq : std_logic_vector(data_width-1 downto 0);
  
BEGIN
-- Port Map
-- readA :: CLOCK clkr ENABLE clkr_en DATA_OUT q ADDRESS radr
-- writeA :: CLOCK clkw ENABLE clkw_en DATA_IN d ADDRESS wadr WRITE_ENABLE we

-- Access memory with non-registered inputs (latency = 1||2)
  IN_PIN :  IF latency < 3 GENERATE
  BEGIN
    PROCESS (clkr)
    BEGIN
      IF (rising_edge(clkr)) THEN
         IF (clkr_en = '1') THEN
          -- workaround for simulation when read address out-of-range during inactive cycle
          --pragma translate_off
          IF (to_integer(unsigned(radr)) < depth) THEN
          --pragma translate_on
          ramq <= mem(to_integer(unsigned(radr)));
          --pragma translate_off
          END IF;
          --pragma translate_on
        END IF;
      END IF;
    END PROCESS;
    PROCESS (clkw)
    BEGIN
      IF (rising_edge(clkw)) THEN
         IF (clkw_en = '1') THEN
          IF (we = '1') THEN
            mem(to_integer(unsigned(wadr))) <= d;
          END IF;
        END IF;
      END IF;
    END PROCESS;
    
  END GENERATE IN_PIN; 

-- Register all non-clock inputs (latency = 3||4)
  IN_REG :  IF latency > 2 GENERATE
    SIGNAL radr_reg : std_logic_vector(addr_width-1 downto 0);
    SIGNAL d_reg : std_logic_vector(data_width-1 downto 0);
    SIGNAL wadr_reg : std_logic_vector(addr_width-1 downto 0);
    SIGNAL we_reg : std_logic;
    
  BEGIN
    PROCESS (clkr)
    BEGIN
      IF (rising_edge(clkr)) THEN
        IF (clkr_en = '1') THEN
          radr_reg <= radr;
        END IF;
      END IF;
    END PROCESS;
    PROCESS (clkw)
    BEGIN
      IF (rising_edge(clkw)) THEN
        IF (clkw_en = '1') THEN
          d_reg <= d;
          wadr_reg <= wadr;
          we_reg <= we;
        END IF;
      END IF;
    END PROCESS;
    
    PROCESS (clkr)
    BEGIN
      IF (rising_edge(clkr)) THEN
         IF (clkr_en = '1') THEN
          -- workaround for simulation when read address out-of-range during inactive cycle
          --pragma translate_off
          IF (to_integer(unsigned(radr_reg)) < depth) THEN
          --pragma translate_on
          ramq <= mem(to_integer(unsigned(radr_reg)));
          --pragma translate_off
          END IF;
          --pragma translate_on
        END IF;
      END IF;
    END PROCESS;
    PROCESS (clkw)
    BEGIN
      IF (rising_edge(clkw)) THEN
         IF (clkw_en = '1') THEN
          IF (we_reg = '1') THEN
            mem(to_integer(unsigned(wadr_reg))) <= d_reg;
          END IF;
        END IF;
      END IF;
    END PROCESS;
    
  END GENERATE IN_REG;

  out_ram : IF latency = 1 GENERATE
  BEGIN
    q <= ramq;
    
  END GENERATE out_ram;

  out_reg1 : IF ((latency = 2) OR (latency = 3)) GENERATE
    SIGNAL tmpq : std_logic_vector(data_width-1 downto 0);
    
  BEGIN
    PROCESS (clkr)
    BEGIN
      IF (rising_edge(clkr)) THEN
        IF (clkr_en = '1') THEN
          tmpq <= ramq;
        END IF;
      END IF;
    END PROCESS;
    
    q <= tmpq;
    
  END GENERATE out_reg1;

  out_reg2 : IF latency = 4 GENERATE
    SIGNAL tmp1q : std_logic_vector(data_width-1 downto 0);
    
    SIGNAL tmp2q : std_logic_vector(data_width-1 downto 0);
    
  BEGIN
    PROCESS (clkr)
    BEGIN
      IF (rising_edge(clkr)) THEN
        IF (clkr_en = '1') THEN
          tmp1q <= ramq;
        END IF;
      END IF;
    END PROCESS;
    
    PROCESS (clkr)
    BEGIN
      IF (rising_edge(clkr)) THEN
        IF (clkr_en = '1') THEN
          tmp2q <= tmp1q;
        END IF;
      END IF;
    END PROCESS;
    
    q <= tmp2q;
    
  END GENERATE out_reg2;


END rtl;

--------> ./rtl.vhdl 
-- ----------------------------------------------------------------------
--  HLS HDL:        VHDL Netlister
--  HLS Version:    10.5c/896140 Production Release
--  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
-- 
--  Generated by:   yl7897@newnano.poly.edu
--  Generated date: Wed Sep 15 01:49:31 2021
-- ----------------------------------------------------------------------

-- 
-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_550_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_550_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_550_8_32_256_256_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_550_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_549_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_549_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_549_8_32_256_256_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_549_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_548_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_548_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_548_8_32_256_256_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_548_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_547_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_547_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_547_8_32_256_256_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_547_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_546_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_546_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_546_8_32_256_256_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_546_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_545_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_545_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_545_8_32_256_256_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_545_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_544_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_544_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_544_8_32_256_256_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_544_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_543_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_543_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_543_8_32_256_256_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_543_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_542_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_542_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_542_8_32_256_256_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_542_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_541_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_541_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_541_8_32_256_256_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_541_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_540_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_540_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_540_8_32_256_256_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_540_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_539_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_539_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_539_8_32_256_256_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_539_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_538_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_538_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_538_8_32_256_256_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_538_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_537_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_537_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_537_8_32_256_256_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_537_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_536_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_536_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_536_8_32_256_256_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_536_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_535_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_535_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_535_8_32_256_256_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_535_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_534_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_534_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_534_8_32_256_256_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_534_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_533_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_533_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_533_8_32_256_256_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_533_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_532_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_532_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_532_8_32_256_256_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_532_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_531_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_531_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_531_8_32_256_256_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_531_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_530_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_530_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_530_8_32_256_256_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_530_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_529_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_529_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_529_8_32_256_256_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_529_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_528_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_528_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_528_8_32_256_256_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_528_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_527_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_527_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_527_8_32_256_256_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_527_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_526_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_526_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_526_8_32_256_256_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_526_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_525_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_525_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_525_8_32_256_256_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_525_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_524_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_524_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_524_8_32_256_256_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_524_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_523_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_523_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_523_8_32_256_256_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_523_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_522_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_522_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_522_8_32_256_256_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_522_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_521_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_521_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_521_8_32_256_256_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_521_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_520_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_520_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_520_8_32_256_256_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_520_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_519_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_519_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_519_8_32_256_256_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_519_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_518_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_518_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_518_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_518_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_517_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_517_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_517_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_517_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_516_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_516_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_516_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_516_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_515_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_515_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_515_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_515_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_514_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_514_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_514_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_514_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_513_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_513_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_513_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_513_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_512_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_512_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_512_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_512_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_511_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_511_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_511_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_511_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_510_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_510_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_510_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_510_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_509_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_509_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_509_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_509_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_508_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_508_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_508_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_508_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_507_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_507_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_507_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_507_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_506_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_506_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_506_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_506_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_505_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_505_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_505_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_505_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_504_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_504_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_504_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_504_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_503_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_503_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_503_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_503_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_502_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_502_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_502_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_502_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_501_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_501_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_501_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_501_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_500_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_500_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_500_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_500_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_499_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_499_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_499_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_499_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_498_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_498_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_498_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_498_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_497_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_497_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_497_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_497_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_496_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_496_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_496_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_496_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_495_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_495_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_495_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_495_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_494_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_494_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_494_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_494_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_493_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_493_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_493_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_493_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_492_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_492_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_492_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_492_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_491_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_491_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_491_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_491_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_490_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_490_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_490_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_490_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_489_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_489_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_489_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_489_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_488_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_488_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_488_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_488_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_487_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_487_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_487_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_487_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_486_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_486_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_486_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_486_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_485_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_485_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_485_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_485_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_484_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_484_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_484_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_484_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_483_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_483_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_483_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_483_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_482_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_482_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_482_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_482_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_481_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_481_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_481_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_481_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_480_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_480_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_480_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_480_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_479_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_479_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_479_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_479_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_478_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_478_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_478_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_478_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_477_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_477_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_477_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_477_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_476_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_476_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_476_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_476_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_475_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_475_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_475_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_475_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_474_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_474_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_474_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_474_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_473_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_473_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_473_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_473_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_472_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_472_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_472_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_472_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_471_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_471_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_471_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_471_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_470_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_470_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_470_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_470_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_469_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_469_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_469_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_469_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_468_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_468_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_468_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_468_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_467_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_467_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_467_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_467_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_466_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_466_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_466_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_466_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_465_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_465_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_465_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_465_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_464_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_464_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_464_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_464_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_463_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_463_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_463_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_463_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_462_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_462_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_462_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_462_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_461_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_461_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_461_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_461_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_460_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_460_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_460_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_460_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_459_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_459_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_459_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_459_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_458_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_458_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_458_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_458_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_457_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_457_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_457_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_457_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_456_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_456_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_456_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_456_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_455_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_455_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_455_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_455_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_454_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_454_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_454_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_454_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_453_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_453_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_453_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_453_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_452_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_452_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_452_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_452_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_451_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_451_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_451_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_451_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_450_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_450_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_450_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_450_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_449_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_449_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_449_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_449_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_448_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_448_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_448_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_448_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_447_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_447_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_447_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_447_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_446_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_446_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_446_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_446_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_445_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_445_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_445_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_445_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_444_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_444_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_444_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_444_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_443_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_443_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_443_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_443_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_442_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_442_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_442_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_442_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_441_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_441_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_441_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_441_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_440_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_440_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_440_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_440_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_439_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_439_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_439_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_439_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_438_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_438_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_438_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_438_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_437_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_437_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_437_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_437_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_436_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_436_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_436_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_436_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_435_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_435_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_435_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_435_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_434_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_434_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_434_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_434_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_433_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_433_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_433_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_433_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_432_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_432_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_432_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_432_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_431_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_431_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_431_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_431_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_430_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_430_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_430_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_430_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_429_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_429_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_429_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_429_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_428_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_428_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_428_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_428_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_427_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_427_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_427_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_427_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_426_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_426_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_426_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_426_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_425_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_425_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_425_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_425_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_424_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_424_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_424_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_424_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_423_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_423_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_423_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_423_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_422_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_422_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_422_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_422_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_421_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_421_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_421_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_421_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_420_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_420_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_420_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_420_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_419_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_419_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_419_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_419_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_418_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_418_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_418_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_418_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_417_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_417_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_417_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_417_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_416_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_416_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_416_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_416_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_415_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_415_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_415_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_415_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_414_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_414_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_414_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_414_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_413_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_413_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_413_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_413_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_412_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_412_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_412_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_412_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_411_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_411_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_411_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_411_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_410_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_410_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_410_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_410_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_409_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_409_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_409_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_409_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_408_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_408_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_408_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_408_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_407_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_407_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_407_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_407_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_406_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_406_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_406_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_406_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_405_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_405_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_405_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_405_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_404_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_404_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_404_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_404_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_403_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_403_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_403_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_403_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_402_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_402_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_402_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_402_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_401_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_401_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_401_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_401_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_400_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_400_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_400_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_400_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_399_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_399_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_399_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_399_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_398_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_398_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_398_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_398_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_397_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_397_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_397_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_397_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_396_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_396_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_396_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_396_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_395_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_395_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_395_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_395_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_394_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_394_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_394_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_394_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_393_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_393_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_393_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_393_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_392_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_392_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_392_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_392_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_391_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_391_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_391_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_391_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_390_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_390_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_390_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_390_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_389_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_389_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_389_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_389_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_388_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_388_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_388_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_388_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_387_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_387_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_387_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_387_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_386_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_386_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_386_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_386_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_385_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_385_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_385_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_385_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_384_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_384_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_384_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_384_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_383_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_383_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_383_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_383_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_382_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_382_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_382_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_382_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_381_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_381_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_381_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_381_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_380_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_380_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_380_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_380_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_379_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_379_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_379_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_379_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_378_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_378_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_378_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_378_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_377_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_377_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_377_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_377_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_376_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_376_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_376_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_376_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_375_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_375_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_375_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_375_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_374_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_374_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_374_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_374_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_373_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_373_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_373_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_373_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_372_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_372_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_372_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_372_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_371_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_371_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_371_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_371_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_370_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_370_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_370_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_370_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_369_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_369_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_369_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_369_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_368_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_368_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_368_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_368_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_367_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_367_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_367_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_367_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_366_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_366_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_366_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_366_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_365_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_365_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_365_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_365_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_364_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_364_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_364_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_364_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_363_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_363_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_363_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_363_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_362_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_362_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_362_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_362_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_361_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_361_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_361_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_361_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_360_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_360_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_360_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_360_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_359_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_359_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_359_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_359_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_358_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_358_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_358_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_358_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_357_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_357_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_357_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_357_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_356_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_356_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_356_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_356_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_355_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_355_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_355_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_355_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_354_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_354_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_354_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_354_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_353_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_353_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_353_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_353_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_352_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_352_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_352_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_352_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_351_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_351_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_351_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_351_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_350_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_350_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_350_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_350_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_349_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_349_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_349_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_349_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_348_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_348_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_348_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_348_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_347_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_347_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_347_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_347_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_346_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_346_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_346_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_346_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_345_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_345_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_345_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_345_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_344_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_344_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_344_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_344_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_343_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_343_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_343_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_343_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_342_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_342_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_342_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_342_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_341_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_341_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_341_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_341_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_340_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_340_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_340_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_340_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_339_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_339_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_339_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_339_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_338_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_338_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_338_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_338_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_337_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_337_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_337_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_337_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_336_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_336_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_336_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_336_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_335_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_335_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_335_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_335_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_334_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_334_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_334_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_334_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_333_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_333_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_333_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_333_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_332_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_332_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_332_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_332_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_331_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_331_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_331_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_331_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_330_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_330_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_330_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_330_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_329_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_329_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_329_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_329_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_328_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_328_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_328_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_328_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_327_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_327_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_327_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_327_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_326_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_326_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_326_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_326_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_325_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_325_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_325_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_325_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_324_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_324_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_324_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_324_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_323_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_323_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_323_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_323_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_322_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_322_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_322_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_322_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_321_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_321_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_321_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_321_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_320_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_320_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_320_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_320_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_319_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_319_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_319_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_319_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_318_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_318_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_318_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_318_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_317_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_317_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_317_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_317_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_316_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_316_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_316_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_316_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_315_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_315_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_315_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_315_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_314_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_314_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_314_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_314_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_313_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_313_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_313_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_313_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_312_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_312_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_312_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_312_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_311_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_311_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_311_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_311_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_310_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_310_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_310_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_310_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_309_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_309_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_309_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_309_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_308_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_308_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_308_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_308_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_307_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_307_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_307_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_307_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_306_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_306_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_306_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_306_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_305_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_305_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_305_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_305_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_304_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_304_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_304_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_304_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_303_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_303_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_303_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_303_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_302_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_302_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_302_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_302_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_301_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_301_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_301_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_301_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_300_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_300_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_300_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_300_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_299_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_299_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_299_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_299_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_298_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_298_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_298_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_298_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_297_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_297_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_297_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_297_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_296_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_296_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_296_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_296_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_295_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_295_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_295_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_295_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_294_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_294_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_294_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_294_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_293_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_293_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_293_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_293_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_292_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_292_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_292_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_292_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_291_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_291_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_291_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_291_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_290_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_290_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_290_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_290_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_289_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_289_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_289_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_289_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_288_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_288_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_288_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_288_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_287_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_287_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_287_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_287_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_286_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_286_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_286_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_286_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_285_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_285_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_285_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_285_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_284_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_284_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_284_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_284_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_283_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_283_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_283_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_283_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_282_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_282_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_282_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_282_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_281_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_281_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_281_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_281_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_280_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_280_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_280_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_280_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_279_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_279_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_279_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_279_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_278_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_278_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_278_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_278_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_277_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_277_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_277_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_277_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_276_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_276_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_276_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_276_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_275_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_275_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_275_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_275_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_274_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_274_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_274_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_274_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_273_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_273_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_273_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_273_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_272_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_272_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_272_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_272_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_271_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_271_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_271_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_271_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_270_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_270_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_270_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_270_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_269_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_269_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_269_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_269_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_268_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_268_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_268_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_268_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_267_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_267_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_267_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_267_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_266_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_266_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_266_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_266_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_265_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_265_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_265_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_265_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_264_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_264_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_264_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_264_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_263_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_263_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_263_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_263_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_262_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_262_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_262_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_262_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_261_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_261_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_261_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_261_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_260_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_260_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_260_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_260_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_259_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_259_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_259_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_259_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_258_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_258_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_258_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_258_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_257_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_257_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_257_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_257_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_256_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_256_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_256_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_256_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_255_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_255_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_255_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_255_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_254_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_254_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_254_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_254_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_253_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_253_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_253_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_253_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_252_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_252_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_252_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_252_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_251_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_251_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_251_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_251_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_250_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_250_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_250_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_250_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_249_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_249_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_249_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_249_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_248_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_248_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_248_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_248_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_247_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_247_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_247_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_247_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_246_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_246_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_246_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_246_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_245_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_245_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_245_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_245_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_244_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_244_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_244_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_244_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_243_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_243_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_243_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_243_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_242_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_242_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_242_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_242_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_241_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_241_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_241_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_241_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_240_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_240_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_240_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_240_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_239_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_239_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_239_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_239_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_238_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_238_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_238_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_238_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_237_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_237_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_237_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_237_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_236_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_236_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_236_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_236_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_235_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_235_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_235_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_235_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_234_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_234_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_234_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_234_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_233_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_233_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_233_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_233_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_232_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_232_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_232_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_232_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_231_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_231_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_231_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_231_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_230_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_230_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_230_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_230_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_229_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_229_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_229_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_229_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_228_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_228_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_228_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_228_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_227_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_227_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_227_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_227_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_226_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_226_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_226_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_226_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_225_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_225_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_225_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_225_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_224_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_224_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_224_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_224_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_223_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_223_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_223_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_223_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_222_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_222_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_222_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_222_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_221_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_221_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_221_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_221_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_220_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_220_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_220_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_220_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_219_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_219_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_219_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_219_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_218_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_218_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_218_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_218_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_217_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_217_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_217_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_217_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_216_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_216_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_216_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_216_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_215_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_215_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_215_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_215_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_214_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_214_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_214_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_214_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_213_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_213_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_213_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_213_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_212_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_212_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_212_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_212_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_211_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_211_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_211_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_211_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_210_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_210_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_210_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_210_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_209_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_209_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_209_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_209_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_208_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_208_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_208_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_208_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_207_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_207_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_207_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_207_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_206_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_206_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_206_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_206_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_205_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_205_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_205_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_205_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_204_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_204_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_204_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_204_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_203_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_203_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_203_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_203_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_202_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_202_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_202_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_202_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_201_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_201_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_201_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_201_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_200_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_200_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_200_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_200_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_199_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_199_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_199_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_199_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_198_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_198_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_198_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_198_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_197_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_197_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_197_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_197_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_196_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_196_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_196_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_196_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_195_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_195_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_195_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_195_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_194_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_194_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_194_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_194_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_193_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_193_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_193_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_193_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_192_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_192_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_192_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_192_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_191_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_191_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_191_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_191_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_190_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_190_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_190_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_190_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_189_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_189_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_189_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_189_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_188_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_188_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_188_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_188_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_187_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_187_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_187_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_187_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_186_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_186_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_186_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_186_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_185_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_185_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_185_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_185_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_184_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_184_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_184_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_184_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_183_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_183_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_183_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_183_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_182_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_182_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_182_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_182_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_181_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_181_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_181_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_181_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_180_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_180_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_180_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_180_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_179_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_179_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_179_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_179_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_178_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_178_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_178_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_178_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_177_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_177_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_177_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_177_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_176_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_176_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_176_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_176_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_175_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_175_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_175_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_175_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_174_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_174_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_174_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_174_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_173_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_173_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_173_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_173_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_172_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_172_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_172_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_172_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_171_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_171_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_171_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_171_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_170_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_170_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_170_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_170_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_169_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_169_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_169_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_169_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_168_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_168_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_168_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_168_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_167_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_167_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_167_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_167_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_166_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_166_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_166_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_166_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_165_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_165_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_165_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_165_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_164_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_164_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_164_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_164_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_163_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_163_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_163_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_163_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_162_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_162_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_162_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_162_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_161_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_161_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_161_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_161_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_160_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_160_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_160_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_160_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_159_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_159_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_159_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_159_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_158_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_158_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_158_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_158_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_157_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_157_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_157_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_157_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_156_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_156_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_156_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_156_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_155_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_155_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_155_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_155_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_154_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_154_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_154_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_154_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_153_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_153_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_153_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_153_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_152_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_152_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_152_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_152_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_151_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_151_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_151_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_151_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_150_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_150_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_150_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_150_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_149_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_149_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_149_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_149_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_148_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_148_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_148_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_148_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_147_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_147_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_147_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_147_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_146_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_146_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_146_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_146_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_145_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_145_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_145_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_145_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_144_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_144_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_144_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_144_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_143_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_143_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_143_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_143_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_142_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_142_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_142_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_142_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_141_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_141_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_141_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_141_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_140_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_140_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_140_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_140_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_139_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_139_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_139_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_139_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_138_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_138_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_138_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_138_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_137_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_137_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_137_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_137_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_136_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_136_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_136_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_136_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_135_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_135_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_135_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_135_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_134_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_134_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_134_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_134_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_133_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_133_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_133_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_133_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_132_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_132_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_132_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_132_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_131_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_131_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_131_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_131_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_130_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_130_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_130_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_130_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_129_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_129_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_129_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_129_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_128_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_128_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_128_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_128_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_127_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_127_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_127_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_127_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_126_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_126_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_126_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_126_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_125_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_125_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_125_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_125_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_124_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_124_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_124_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_124_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_123_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_123_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_123_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_123_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_122_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_122_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_122_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_122_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_121_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_121_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_121_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_121_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_120_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_120_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_120_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_120_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_119_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_119_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_119_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_119_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_118_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_118_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_118_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_118_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_117_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_117_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_117_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_117_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_116_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_116_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_116_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_116_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_115_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_115_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_115_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_115_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_114_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_114_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_114_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_114_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_113_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_113_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_113_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_113_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_112_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_112_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_112_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_112_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_111_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_111_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_111_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_111_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_110_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_110_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_110_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_110_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_109_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_109_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_109_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_109_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_108_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_108_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_108_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_108_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_107_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_107_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_107_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_107_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_106_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_106_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_106_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_106_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_105_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_105_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_105_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_105_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_104_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_104_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_104_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_104_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_103_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_103_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_103_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_103_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_102_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_102_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_102_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_102_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_101_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_101_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_101_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_101_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_100_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_100_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_100_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_100_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_99_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_99_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_99_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_99_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_98_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_98_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_98_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_98_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_97_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_97_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_97_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_97_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_96_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_96_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_96_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_96_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_95_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_95_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_95_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_95_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_94_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_94_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_94_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_94_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_93_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_93_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_93_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_93_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_92_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_92_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_92_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_92_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_91_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_91_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_91_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_91_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_90_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_90_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_90_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_90_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_89_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_89_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_89_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_89_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_88_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_88_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_88_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_88_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_87_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_87_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_87_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_87_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_86_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_86_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_86_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_86_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_85_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_85_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_85_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_85_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_84_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_84_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_84_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_84_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_83_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_83_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_83_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_83_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_82_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_82_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_82_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_82_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_81_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_81_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_81_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_81_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_80_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_80_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_80_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_80_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_79_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_79_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_79_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_79_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_78_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_78_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_78_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_78_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_77_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_77_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_77_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_77_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_76_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_76_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_76_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_76_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_75_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_75_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_75_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_75_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_74_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_74_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_74_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_74_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_73_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_73_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_73_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_73_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_72_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_72_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_72_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_72_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_71_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_71_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_71_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_71_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_70_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_70_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_70_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_70_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_69_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_69_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_69_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_69_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_68_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_68_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_68_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_68_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_67_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_67_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_67_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_67_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_66_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_66_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_66_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_66_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_65_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_65_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_65_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_65_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_64_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_64_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_64_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_64_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_63_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_63_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_63_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_63_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_62_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_62_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_62_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_62_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_61_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_61_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_61_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_61_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_60_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_60_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_60_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_60_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_59_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_59_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_59_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_59_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_58_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_58_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_58_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_58_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_57_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_57_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_57_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_57_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_56_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_56_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_56_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_56_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_55_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_55_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_55_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_55_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_54_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_54_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_54_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_54_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_53_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_53_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_53_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_53_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_52_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_52_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_52_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_52_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_51_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_51_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_51_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_51_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_50_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_50_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_50_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_50_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_49_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_49_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_49_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_49_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_48_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_48_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_48_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_48_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_47_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_47_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_47_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_47_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_46_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_46_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_46_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_46_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_45_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_45_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_45_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_45_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_44_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_44_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_44_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_44_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_43_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_43_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_43_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_43_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_42_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_42_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_42_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_42_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_41_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_41_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_41_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_41_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_40_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_40_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_40_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_40_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_39_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_39_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_39_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_39_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_38_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_38_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_38_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_38_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_37_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_37_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_37_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_37_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_36_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_36_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_36_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_36_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_35_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_35_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_35_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_35_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_34_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_34_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_34_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_34_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_33_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_33_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_33_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_33_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_32_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_32_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_32_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_32_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_31_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_31_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_31_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_31_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_30_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_30_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_30_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_30_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_29_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_29_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_29_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_29_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_28_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_28_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_28_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_28_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_27_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_27_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_27_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_27_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_26_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_26_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_26_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_26_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_25_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_25_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_25_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_25_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_24_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_24_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_24_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_24_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_23_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_23_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_23_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_23_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_22_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_22_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_22_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_22_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_21_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_21_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_21_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_21_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_20_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_20_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_20_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_20_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_19_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_19_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_19_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_19_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_18_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_18_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_18_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_18_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_17_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_17_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_17_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_17_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_16_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_16_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_16_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_16_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_15_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_15_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_15_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_15_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_14_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_14_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_14_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_14_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_13_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_13_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_13_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_13_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_12_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_12_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_12_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_12_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_11_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_11_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_11_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_11_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_10_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_10_4_32_16_16_32_1_gen
    IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_10_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_10_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_9_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_9_4_32_16_16_32_1_gen IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_9_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_9_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_8_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_8_4_32_16_16_32_1_gen IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_8_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_8_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_7_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_7_4_32_16_16_32_1_gen IS
  PORT(
    clkr_en : OUT STD_LOGIC;
    clkw_en : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    clkr : IN STD_LOGIC;
    clkr_en_d : IN STD_LOGIC;
    clkw_en_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_7_4_32_16_16_32_1_gen;

ARCHITECTURE v14 OF peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_7_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkr_en <= (clkr_en_d);
  clkw_en <= (clkw_en_d);
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_core_fsm
--  FSM Module
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_core_core_fsm IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    fsm_output : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
    INNER_LOOP1_C_0_tr0 : IN STD_LOGIC;
    INNER_LOOP2_C_0_tr0 : IN STD_LOGIC;
    STAGE_LOOP_C_2_tr0 : IN STD_LOGIC;
    INNER_LOOP3_C_0_tr0 : IN STD_LOGIC;
    INNER_LOOP4_C_0_tr0 : IN STD_LOGIC;
    INNER_LOOP4_C_0_tr1 : IN STD_LOGIC
  );
END peaseNTT_core_core_fsm;

ARCHITECTURE v14 OF peaseNTT_core_core_fsm IS
  -- Default Constants

  -- FSM State Type Declaration for peaseNTT_core_core_fsm_1
  TYPE peaseNTT_core_core_fsm_1_ST IS (main_C_0, STAGE_LOOP_C_0, INNER_LOOP1_C_0,
      STAGE_LOOP_C_1, INNER_LOOP2_C_0, STAGE_LOOP_C_2, STAGE_LOOP1_C_0, INNER_LOOP3_C_0,
      STAGE_LOOP1_C_1, INNER_LOOP4_C_0, main_C_1);

  SIGNAL state_var : peaseNTT_core_core_fsm_1_ST;
  SIGNAL state_var_NS : peaseNTT_core_core_fsm_1_ST;

BEGIN
  peaseNTT_core_core_fsm_1 : PROCESS (INNER_LOOP1_C_0_tr0, INNER_LOOP2_C_0_tr0, STAGE_LOOP_C_2_tr0,
      INNER_LOOP3_C_0_tr0, INNER_LOOP4_C_0_tr0, INNER_LOOP4_C_0_tr1, state_var)
  BEGIN
    CASE state_var IS
      WHEN STAGE_LOOP_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000010");
        state_var_NS <= INNER_LOOP1_C_0;
      WHEN INNER_LOOP1_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000100");
        IF ( INNER_LOOP1_C_0_tr0 = '1' ) THEN
          state_var_NS <= STAGE_LOOP_C_1;
        ELSE
          state_var_NS <= INNER_LOOP1_C_0;
        END IF;
      WHEN STAGE_LOOP_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000001000");
        state_var_NS <= INNER_LOOP2_C_0;
      WHEN INNER_LOOP2_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000010000");
        IF ( INNER_LOOP2_C_0_tr0 = '1' ) THEN
          state_var_NS <= STAGE_LOOP_C_2;
        ELSE
          state_var_NS <= INNER_LOOP2_C_0;
        END IF;
      WHEN STAGE_LOOP_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000100000");
        IF ( STAGE_LOOP_C_2_tr0 = '1' ) THEN
          state_var_NS <= STAGE_LOOP1_C_0;
        ELSE
          state_var_NS <= STAGE_LOOP_C_0;
        END IF;
      WHEN STAGE_LOOP1_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001000000");
        state_var_NS <= INNER_LOOP3_C_0;
      WHEN INNER_LOOP3_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010000000");
        IF ( INNER_LOOP3_C_0_tr0 = '1' ) THEN
          state_var_NS <= STAGE_LOOP1_C_1;
        ELSE
          state_var_NS <= INNER_LOOP3_C_0;
        END IF;
      WHEN STAGE_LOOP1_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100000000");
        state_var_NS <= INNER_LOOP4_C_0;
      WHEN INNER_LOOP4_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000000000");
        IF ( INNER_LOOP4_C_0_tr0 = '1' ) THEN
          state_var_NS <= main_C_1;
        ELSIF ( INNER_LOOP4_C_0_tr1 = '1' ) THEN
          state_var_NS <= INNER_LOOP4_C_0;
        ELSE
          state_var_NS <= STAGE_LOOP1_C_0;
        END IF;
      WHEN main_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000000000");
        state_var_NS <= main_C_0;
      -- main_C_0
      WHEN OTHERS =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000001");
        state_var_NS <= STAGE_LOOP_C_0;
    END CASE;
  END PROCESS peaseNTT_core_core_fsm_1;

  peaseNTT_core_core_fsm_1_REG : PROCESS (clk)
  BEGIN
    IF clk'event AND ( clk = '1' ) THEN
      IF ( rst = '1' ) THEN
        state_var <= main_C_0;
      ELSE
        state_var <= state_var_NS;
      END IF;
    END IF;
  END PROCESS peaseNTT_core_core_fsm_1_REG;

END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_core_wait_dp IS
  PORT(
    yt_rsc_0_0_cgo_iro : IN STD_LOGIC;
    yt_rsc_0_0_i_clkr_en_d : OUT STD_LOGIC;
    yt_rsc_0_16_cgo_iro : IN STD_LOGIC;
    yt_rsc_0_16_i_clkr_en_d : OUT STD_LOGIC;
    yt_rsc_1_0_cgo_iro : IN STD_LOGIC;
    yt_rsc_1_0_i_clkr_en_d : OUT STD_LOGIC;
    yt_rsc_1_16_cgo_iro : IN STD_LOGIC;
    yt_rsc_1_16_i_clkr_en_d : OUT STD_LOGIC;
    yt_rsc_2_0_cgo_iro : IN STD_LOGIC;
    yt_rsc_2_0_i_clkr_en_d : OUT STD_LOGIC;
    yt_rsc_2_16_cgo_iro : IN STD_LOGIC;
    yt_rsc_2_16_i_clkr_en_d : OUT STD_LOGIC;
    yt_rsc_3_0_cgo_iro : IN STD_LOGIC;
    yt_rsc_3_0_i_clkr_en_d : OUT STD_LOGIC;
    yt_rsc_3_16_cgo_iro : IN STD_LOGIC;
    yt_rsc_3_16_i_clkr_en_d : OUT STD_LOGIC;
    yt_rsc_4_0_cgo_iro : IN STD_LOGIC;
    yt_rsc_4_0_i_clkr_en_d : OUT STD_LOGIC;
    yt_rsc_4_16_cgo_iro : IN STD_LOGIC;
    yt_rsc_4_16_i_clkr_en_d : OUT STD_LOGIC;
    yt_rsc_5_0_cgo_iro : IN STD_LOGIC;
    yt_rsc_5_0_i_clkr_en_d : OUT STD_LOGIC;
    yt_rsc_5_16_cgo_iro : IN STD_LOGIC;
    yt_rsc_5_16_i_clkr_en_d : OUT STD_LOGIC;
    yt_rsc_6_0_cgo_iro : IN STD_LOGIC;
    yt_rsc_6_0_i_clkr_en_d : OUT STD_LOGIC;
    yt_rsc_6_16_cgo_iro : IN STD_LOGIC;
    yt_rsc_6_16_i_clkr_en_d : OUT STD_LOGIC;
    yt_rsc_7_0_cgo_iro : IN STD_LOGIC;
    yt_rsc_7_0_i_clkr_en_d : OUT STD_LOGIC;
    yt_rsc_7_16_cgo_iro : IN STD_LOGIC;
    yt_rsc_7_16_i_clkr_en_d : OUT STD_LOGIC;
    ensig_cgo_iro : IN STD_LOGIC;
    ensig_cgo_iro_17 : IN STD_LOGIC;
    yt_rsc_0_0_cgo : IN STD_LOGIC;
    yt_rsc_0_16_cgo : IN STD_LOGIC;
    yt_rsc_1_0_cgo : IN STD_LOGIC;
    yt_rsc_1_16_cgo : IN STD_LOGIC;
    yt_rsc_2_0_cgo : IN STD_LOGIC;
    yt_rsc_2_16_cgo : IN STD_LOGIC;
    yt_rsc_3_0_cgo : IN STD_LOGIC;
    yt_rsc_3_16_cgo : IN STD_LOGIC;
    yt_rsc_4_0_cgo : IN STD_LOGIC;
    yt_rsc_4_16_cgo : IN STD_LOGIC;
    yt_rsc_5_0_cgo : IN STD_LOGIC;
    yt_rsc_5_16_cgo : IN STD_LOGIC;
    yt_rsc_6_0_cgo : IN STD_LOGIC;
    yt_rsc_6_16_cgo : IN STD_LOGIC;
    yt_rsc_7_0_cgo : IN STD_LOGIC;
    yt_rsc_7_16_cgo : IN STD_LOGIC;
    ensig_cgo : IN STD_LOGIC;
    mult_t_mul_cmp_en : OUT STD_LOGIC;
    ensig_cgo_17 : IN STD_LOGIC;
    mult_z_mul_cmp_1_en : OUT STD_LOGIC
  );
END peaseNTT_core_wait_dp;

ARCHITECTURE v14 OF peaseNTT_core_wait_dp IS
  -- Default Constants

BEGIN
  yt_rsc_0_0_i_clkr_en_d <= yt_rsc_0_0_cgo OR yt_rsc_0_0_cgo_iro;
  yt_rsc_0_16_i_clkr_en_d <= yt_rsc_0_16_cgo OR yt_rsc_0_16_cgo_iro;
  yt_rsc_1_0_i_clkr_en_d <= yt_rsc_1_0_cgo OR yt_rsc_1_0_cgo_iro;
  yt_rsc_1_16_i_clkr_en_d <= yt_rsc_1_16_cgo OR yt_rsc_1_16_cgo_iro;
  yt_rsc_2_0_i_clkr_en_d <= yt_rsc_2_0_cgo OR yt_rsc_2_0_cgo_iro;
  yt_rsc_2_16_i_clkr_en_d <= yt_rsc_2_16_cgo OR yt_rsc_2_16_cgo_iro;
  yt_rsc_3_0_i_clkr_en_d <= yt_rsc_3_0_cgo OR yt_rsc_3_0_cgo_iro;
  yt_rsc_3_16_i_clkr_en_d <= yt_rsc_3_16_cgo OR yt_rsc_3_16_cgo_iro;
  yt_rsc_4_0_i_clkr_en_d <= yt_rsc_4_0_cgo OR yt_rsc_4_0_cgo_iro;
  yt_rsc_4_16_i_clkr_en_d <= yt_rsc_4_16_cgo OR yt_rsc_4_16_cgo_iro;
  yt_rsc_5_0_i_clkr_en_d <= yt_rsc_5_0_cgo OR yt_rsc_5_0_cgo_iro;
  yt_rsc_5_16_i_clkr_en_d <= yt_rsc_5_16_cgo OR yt_rsc_5_16_cgo_iro;
  yt_rsc_6_0_i_clkr_en_d <= yt_rsc_6_0_cgo OR yt_rsc_6_0_cgo_iro;
  yt_rsc_6_16_i_clkr_en_d <= yt_rsc_6_16_cgo OR yt_rsc_6_16_cgo_iro;
  yt_rsc_7_0_i_clkr_en_d <= yt_rsc_7_0_cgo OR yt_rsc_7_0_cgo_iro;
  yt_rsc_7_16_i_clkr_en_d <= yt_rsc_7_16_cgo OR yt_rsc_7_16_cgo_iro;
  mult_t_mul_cmp_en <= ensig_cgo OR ensig_cgo_iro;
  mult_z_mul_cmp_1_en <= ensig_cgo_17 OR ensig_cgo_iro_17;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_core IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_triosy_0_0_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_1_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_2_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_3_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_4_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_5_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_6_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_7_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_8_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_9_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_10_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_11_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_12_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_13_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_14_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_15_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_16_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_17_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_18_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_19_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_20_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_21_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_22_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_23_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_24_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_25_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_26_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_27_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_28_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_29_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_30_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_31_lz : OUT STD_LOGIC;
    xt_rsc_triosy_1_0_lz : OUT STD_LOGIC;
    xt_rsc_triosy_1_1_lz : OUT STD_LOGIC;
    xt_rsc_triosy_1_2_lz : OUT STD_LOGIC;
    xt_rsc_triosy_1_3_lz : OUT STD_LOGIC;
    xt_rsc_triosy_1_4_lz : OUT STD_LOGIC;
    xt_rsc_triosy_1_5_lz : OUT STD_LOGIC;
    xt_rsc_triosy_1_6_lz : OUT STD_LOGIC;
    xt_rsc_triosy_1_7_lz : OUT STD_LOGIC;
    xt_rsc_triosy_1_8_lz : OUT STD_LOGIC;
    xt_rsc_triosy_1_9_lz : OUT STD_LOGIC;
    xt_rsc_triosy_1_10_lz : OUT STD_LOGIC;
    xt_rsc_triosy_1_11_lz : OUT STD_LOGIC;
    xt_rsc_triosy_1_12_lz : OUT STD_LOGIC;
    xt_rsc_triosy_1_13_lz : OUT STD_LOGIC;
    xt_rsc_triosy_1_14_lz : OUT STD_LOGIC;
    xt_rsc_triosy_1_15_lz : OUT STD_LOGIC;
    xt_rsc_triosy_1_16_lz : OUT STD_LOGIC;
    xt_rsc_triosy_1_17_lz : OUT STD_LOGIC;
    xt_rsc_triosy_1_18_lz : OUT STD_LOGIC;
    xt_rsc_triosy_1_19_lz : OUT STD_LOGIC;
    xt_rsc_triosy_1_20_lz : OUT STD_LOGIC;
    xt_rsc_triosy_1_21_lz : OUT STD_LOGIC;
    xt_rsc_triosy_1_22_lz : OUT STD_LOGIC;
    xt_rsc_triosy_1_23_lz : OUT STD_LOGIC;
    xt_rsc_triosy_1_24_lz : OUT STD_LOGIC;
    xt_rsc_triosy_1_25_lz : OUT STD_LOGIC;
    xt_rsc_triosy_1_26_lz : OUT STD_LOGIC;
    xt_rsc_triosy_1_27_lz : OUT STD_LOGIC;
    xt_rsc_triosy_1_28_lz : OUT STD_LOGIC;
    xt_rsc_triosy_1_29_lz : OUT STD_LOGIC;
    xt_rsc_triosy_1_30_lz : OUT STD_LOGIC;
    xt_rsc_triosy_1_31_lz : OUT STD_LOGIC;
    xt_rsc_triosy_2_0_lz : OUT STD_LOGIC;
    xt_rsc_triosy_2_1_lz : OUT STD_LOGIC;
    xt_rsc_triosy_2_2_lz : OUT STD_LOGIC;
    xt_rsc_triosy_2_3_lz : OUT STD_LOGIC;
    xt_rsc_triosy_2_4_lz : OUT STD_LOGIC;
    xt_rsc_triosy_2_5_lz : OUT STD_LOGIC;
    xt_rsc_triosy_2_6_lz : OUT STD_LOGIC;
    xt_rsc_triosy_2_7_lz : OUT STD_LOGIC;
    xt_rsc_triosy_2_8_lz : OUT STD_LOGIC;
    xt_rsc_triosy_2_9_lz : OUT STD_LOGIC;
    xt_rsc_triosy_2_10_lz : OUT STD_LOGIC;
    xt_rsc_triosy_2_11_lz : OUT STD_LOGIC;
    xt_rsc_triosy_2_12_lz : OUT STD_LOGIC;
    xt_rsc_triosy_2_13_lz : OUT STD_LOGIC;
    xt_rsc_triosy_2_14_lz : OUT STD_LOGIC;
    xt_rsc_triosy_2_15_lz : OUT STD_LOGIC;
    xt_rsc_triosy_2_16_lz : OUT STD_LOGIC;
    xt_rsc_triosy_2_17_lz : OUT STD_LOGIC;
    xt_rsc_triosy_2_18_lz : OUT STD_LOGIC;
    xt_rsc_triosy_2_19_lz : OUT STD_LOGIC;
    xt_rsc_triosy_2_20_lz : OUT STD_LOGIC;
    xt_rsc_triosy_2_21_lz : OUT STD_LOGIC;
    xt_rsc_triosy_2_22_lz : OUT STD_LOGIC;
    xt_rsc_triosy_2_23_lz : OUT STD_LOGIC;
    xt_rsc_triosy_2_24_lz : OUT STD_LOGIC;
    xt_rsc_triosy_2_25_lz : OUT STD_LOGIC;
    xt_rsc_triosy_2_26_lz : OUT STD_LOGIC;
    xt_rsc_triosy_2_27_lz : OUT STD_LOGIC;
    xt_rsc_triosy_2_28_lz : OUT STD_LOGIC;
    xt_rsc_triosy_2_29_lz : OUT STD_LOGIC;
    xt_rsc_triosy_2_30_lz : OUT STD_LOGIC;
    xt_rsc_triosy_2_31_lz : OUT STD_LOGIC;
    xt_rsc_triosy_3_0_lz : OUT STD_LOGIC;
    xt_rsc_triosy_3_1_lz : OUT STD_LOGIC;
    xt_rsc_triosy_3_2_lz : OUT STD_LOGIC;
    xt_rsc_triosy_3_3_lz : OUT STD_LOGIC;
    xt_rsc_triosy_3_4_lz : OUT STD_LOGIC;
    xt_rsc_triosy_3_5_lz : OUT STD_LOGIC;
    xt_rsc_triosy_3_6_lz : OUT STD_LOGIC;
    xt_rsc_triosy_3_7_lz : OUT STD_LOGIC;
    xt_rsc_triosy_3_8_lz : OUT STD_LOGIC;
    xt_rsc_triosy_3_9_lz : OUT STD_LOGIC;
    xt_rsc_triosy_3_10_lz : OUT STD_LOGIC;
    xt_rsc_triosy_3_11_lz : OUT STD_LOGIC;
    xt_rsc_triosy_3_12_lz : OUT STD_LOGIC;
    xt_rsc_triosy_3_13_lz : OUT STD_LOGIC;
    xt_rsc_triosy_3_14_lz : OUT STD_LOGIC;
    xt_rsc_triosy_3_15_lz : OUT STD_LOGIC;
    xt_rsc_triosy_3_16_lz : OUT STD_LOGIC;
    xt_rsc_triosy_3_17_lz : OUT STD_LOGIC;
    xt_rsc_triosy_3_18_lz : OUT STD_LOGIC;
    xt_rsc_triosy_3_19_lz : OUT STD_LOGIC;
    xt_rsc_triosy_3_20_lz : OUT STD_LOGIC;
    xt_rsc_triosy_3_21_lz : OUT STD_LOGIC;
    xt_rsc_triosy_3_22_lz : OUT STD_LOGIC;
    xt_rsc_triosy_3_23_lz : OUT STD_LOGIC;
    xt_rsc_triosy_3_24_lz : OUT STD_LOGIC;
    xt_rsc_triosy_3_25_lz : OUT STD_LOGIC;
    xt_rsc_triosy_3_26_lz : OUT STD_LOGIC;
    xt_rsc_triosy_3_27_lz : OUT STD_LOGIC;
    xt_rsc_triosy_3_28_lz : OUT STD_LOGIC;
    xt_rsc_triosy_3_29_lz : OUT STD_LOGIC;
    xt_rsc_triosy_3_30_lz : OUT STD_LOGIC;
    xt_rsc_triosy_3_31_lz : OUT STD_LOGIC;
    xt_rsc_triosy_4_0_lz : OUT STD_LOGIC;
    xt_rsc_triosy_4_1_lz : OUT STD_LOGIC;
    xt_rsc_triosy_4_2_lz : OUT STD_LOGIC;
    xt_rsc_triosy_4_3_lz : OUT STD_LOGIC;
    xt_rsc_triosy_4_4_lz : OUT STD_LOGIC;
    xt_rsc_triosy_4_5_lz : OUT STD_LOGIC;
    xt_rsc_triosy_4_6_lz : OUT STD_LOGIC;
    xt_rsc_triosy_4_7_lz : OUT STD_LOGIC;
    xt_rsc_triosy_4_8_lz : OUT STD_LOGIC;
    xt_rsc_triosy_4_9_lz : OUT STD_LOGIC;
    xt_rsc_triosy_4_10_lz : OUT STD_LOGIC;
    xt_rsc_triosy_4_11_lz : OUT STD_LOGIC;
    xt_rsc_triosy_4_12_lz : OUT STD_LOGIC;
    xt_rsc_triosy_4_13_lz : OUT STD_LOGIC;
    xt_rsc_triosy_4_14_lz : OUT STD_LOGIC;
    xt_rsc_triosy_4_15_lz : OUT STD_LOGIC;
    xt_rsc_triosy_4_16_lz : OUT STD_LOGIC;
    xt_rsc_triosy_4_17_lz : OUT STD_LOGIC;
    xt_rsc_triosy_4_18_lz : OUT STD_LOGIC;
    xt_rsc_triosy_4_19_lz : OUT STD_LOGIC;
    xt_rsc_triosy_4_20_lz : OUT STD_LOGIC;
    xt_rsc_triosy_4_21_lz : OUT STD_LOGIC;
    xt_rsc_triosy_4_22_lz : OUT STD_LOGIC;
    xt_rsc_triosy_4_23_lz : OUT STD_LOGIC;
    xt_rsc_triosy_4_24_lz : OUT STD_LOGIC;
    xt_rsc_triosy_4_25_lz : OUT STD_LOGIC;
    xt_rsc_triosy_4_26_lz : OUT STD_LOGIC;
    xt_rsc_triosy_4_27_lz : OUT STD_LOGIC;
    xt_rsc_triosy_4_28_lz : OUT STD_LOGIC;
    xt_rsc_triosy_4_29_lz : OUT STD_LOGIC;
    xt_rsc_triosy_4_30_lz : OUT STD_LOGIC;
    xt_rsc_triosy_4_31_lz : OUT STD_LOGIC;
    xt_rsc_triosy_5_0_lz : OUT STD_LOGIC;
    xt_rsc_triosy_5_1_lz : OUT STD_LOGIC;
    xt_rsc_triosy_5_2_lz : OUT STD_LOGIC;
    xt_rsc_triosy_5_3_lz : OUT STD_LOGIC;
    xt_rsc_triosy_5_4_lz : OUT STD_LOGIC;
    xt_rsc_triosy_5_5_lz : OUT STD_LOGIC;
    xt_rsc_triosy_5_6_lz : OUT STD_LOGIC;
    xt_rsc_triosy_5_7_lz : OUT STD_LOGIC;
    xt_rsc_triosy_5_8_lz : OUT STD_LOGIC;
    xt_rsc_triosy_5_9_lz : OUT STD_LOGIC;
    xt_rsc_triosy_5_10_lz : OUT STD_LOGIC;
    xt_rsc_triosy_5_11_lz : OUT STD_LOGIC;
    xt_rsc_triosy_5_12_lz : OUT STD_LOGIC;
    xt_rsc_triosy_5_13_lz : OUT STD_LOGIC;
    xt_rsc_triosy_5_14_lz : OUT STD_LOGIC;
    xt_rsc_triosy_5_15_lz : OUT STD_LOGIC;
    xt_rsc_triosy_5_16_lz : OUT STD_LOGIC;
    xt_rsc_triosy_5_17_lz : OUT STD_LOGIC;
    xt_rsc_triosy_5_18_lz : OUT STD_LOGIC;
    xt_rsc_triosy_5_19_lz : OUT STD_LOGIC;
    xt_rsc_triosy_5_20_lz : OUT STD_LOGIC;
    xt_rsc_triosy_5_21_lz : OUT STD_LOGIC;
    xt_rsc_triosy_5_22_lz : OUT STD_LOGIC;
    xt_rsc_triosy_5_23_lz : OUT STD_LOGIC;
    xt_rsc_triosy_5_24_lz : OUT STD_LOGIC;
    xt_rsc_triosy_5_25_lz : OUT STD_LOGIC;
    xt_rsc_triosy_5_26_lz : OUT STD_LOGIC;
    xt_rsc_triosy_5_27_lz : OUT STD_LOGIC;
    xt_rsc_triosy_5_28_lz : OUT STD_LOGIC;
    xt_rsc_triosy_5_29_lz : OUT STD_LOGIC;
    xt_rsc_triosy_5_30_lz : OUT STD_LOGIC;
    xt_rsc_triosy_5_31_lz : OUT STD_LOGIC;
    xt_rsc_triosy_6_0_lz : OUT STD_LOGIC;
    xt_rsc_triosy_6_1_lz : OUT STD_LOGIC;
    xt_rsc_triosy_6_2_lz : OUT STD_LOGIC;
    xt_rsc_triosy_6_3_lz : OUT STD_LOGIC;
    xt_rsc_triosy_6_4_lz : OUT STD_LOGIC;
    xt_rsc_triosy_6_5_lz : OUT STD_LOGIC;
    xt_rsc_triosy_6_6_lz : OUT STD_LOGIC;
    xt_rsc_triosy_6_7_lz : OUT STD_LOGIC;
    xt_rsc_triosy_6_8_lz : OUT STD_LOGIC;
    xt_rsc_triosy_6_9_lz : OUT STD_LOGIC;
    xt_rsc_triosy_6_10_lz : OUT STD_LOGIC;
    xt_rsc_triosy_6_11_lz : OUT STD_LOGIC;
    xt_rsc_triosy_6_12_lz : OUT STD_LOGIC;
    xt_rsc_triosy_6_13_lz : OUT STD_LOGIC;
    xt_rsc_triosy_6_14_lz : OUT STD_LOGIC;
    xt_rsc_triosy_6_15_lz : OUT STD_LOGIC;
    xt_rsc_triosy_6_16_lz : OUT STD_LOGIC;
    xt_rsc_triosy_6_17_lz : OUT STD_LOGIC;
    xt_rsc_triosy_6_18_lz : OUT STD_LOGIC;
    xt_rsc_triosy_6_19_lz : OUT STD_LOGIC;
    xt_rsc_triosy_6_20_lz : OUT STD_LOGIC;
    xt_rsc_triosy_6_21_lz : OUT STD_LOGIC;
    xt_rsc_triosy_6_22_lz : OUT STD_LOGIC;
    xt_rsc_triosy_6_23_lz : OUT STD_LOGIC;
    xt_rsc_triosy_6_24_lz : OUT STD_LOGIC;
    xt_rsc_triosy_6_25_lz : OUT STD_LOGIC;
    xt_rsc_triosy_6_26_lz : OUT STD_LOGIC;
    xt_rsc_triosy_6_27_lz : OUT STD_LOGIC;
    xt_rsc_triosy_6_28_lz : OUT STD_LOGIC;
    xt_rsc_triosy_6_29_lz : OUT STD_LOGIC;
    xt_rsc_triosy_6_30_lz : OUT STD_LOGIC;
    xt_rsc_triosy_6_31_lz : OUT STD_LOGIC;
    xt_rsc_triosy_7_0_lz : OUT STD_LOGIC;
    xt_rsc_triosy_7_1_lz : OUT STD_LOGIC;
    xt_rsc_triosy_7_2_lz : OUT STD_LOGIC;
    xt_rsc_triosy_7_3_lz : OUT STD_LOGIC;
    xt_rsc_triosy_7_4_lz : OUT STD_LOGIC;
    xt_rsc_triosy_7_5_lz : OUT STD_LOGIC;
    xt_rsc_triosy_7_6_lz : OUT STD_LOGIC;
    xt_rsc_triosy_7_7_lz : OUT STD_LOGIC;
    xt_rsc_triosy_7_8_lz : OUT STD_LOGIC;
    xt_rsc_triosy_7_9_lz : OUT STD_LOGIC;
    xt_rsc_triosy_7_10_lz : OUT STD_LOGIC;
    xt_rsc_triosy_7_11_lz : OUT STD_LOGIC;
    xt_rsc_triosy_7_12_lz : OUT STD_LOGIC;
    xt_rsc_triosy_7_13_lz : OUT STD_LOGIC;
    xt_rsc_triosy_7_14_lz : OUT STD_LOGIC;
    xt_rsc_triosy_7_15_lz : OUT STD_LOGIC;
    xt_rsc_triosy_7_16_lz : OUT STD_LOGIC;
    xt_rsc_triosy_7_17_lz : OUT STD_LOGIC;
    xt_rsc_triosy_7_18_lz : OUT STD_LOGIC;
    xt_rsc_triosy_7_19_lz : OUT STD_LOGIC;
    xt_rsc_triosy_7_20_lz : OUT STD_LOGIC;
    xt_rsc_triosy_7_21_lz : OUT STD_LOGIC;
    xt_rsc_triosy_7_22_lz : OUT STD_LOGIC;
    xt_rsc_triosy_7_23_lz : OUT STD_LOGIC;
    xt_rsc_triosy_7_24_lz : OUT STD_LOGIC;
    xt_rsc_triosy_7_25_lz : OUT STD_LOGIC;
    xt_rsc_triosy_7_26_lz : OUT STD_LOGIC;
    xt_rsc_triosy_7_27_lz : OUT STD_LOGIC;
    xt_rsc_triosy_7_28_lz : OUT STD_LOGIC;
    xt_rsc_triosy_7_29_lz : OUT STD_LOGIC;
    xt_rsc_triosy_7_30_lz : OUT STD_LOGIC;
    xt_rsc_triosy_7_31_lz : OUT STD_LOGIC;
    p_rsc_dat : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    p_rsc_triosy_lz : OUT STD_LOGIC;
    r_rsc_triosy_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_0_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_1_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_2_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_3_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_4_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_5_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_6_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_7_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_8_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_9_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_10_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_11_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_12_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_13_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_14_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_15_lz : OUT STD_LOGIC;
    twiddle_h_rsc_triosy_0_0_lz : OUT STD_LOGIC;
    twiddle_h_rsc_triosy_0_1_lz : OUT STD_LOGIC;
    twiddle_h_rsc_triosy_0_2_lz : OUT STD_LOGIC;
    twiddle_h_rsc_triosy_0_3_lz : OUT STD_LOGIC;
    twiddle_h_rsc_triosy_0_4_lz : OUT STD_LOGIC;
    twiddle_h_rsc_triosy_0_5_lz : OUT STD_LOGIC;
    twiddle_h_rsc_triosy_0_6_lz : OUT STD_LOGIC;
    twiddle_h_rsc_triosy_0_7_lz : OUT STD_LOGIC;
    twiddle_h_rsc_triosy_0_8_lz : OUT STD_LOGIC;
    twiddle_h_rsc_triosy_0_9_lz : OUT STD_LOGIC;
    twiddle_h_rsc_triosy_0_10_lz : OUT STD_LOGIC;
    twiddle_h_rsc_triosy_0_11_lz : OUT STD_LOGIC;
    twiddle_h_rsc_triosy_0_12_lz : OUT STD_LOGIC;
    twiddle_h_rsc_triosy_0_13_lz : OUT STD_LOGIC;
    twiddle_h_rsc_triosy_0_14_lz : OUT STD_LOGIC;
    twiddle_h_rsc_triosy_0_15_lz : OUT STD_LOGIC;
    yt_rsc_0_0_i_clkr_en_d : OUT STD_LOGIC;
    yt_rsc_0_0_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_1_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_2_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_3_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_4_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_5_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_6_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_7_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_8_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_9_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_10_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_11_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_12_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_13_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_14_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_15_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_16_i_clkr_en_d : OUT STD_LOGIC;
    yt_rsc_0_16_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_17_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_18_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_19_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_20_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_21_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_22_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_23_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_24_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_25_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_26_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_27_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_28_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_29_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_30_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_31_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_0_i_clkr_en_d : OUT STD_LOGIC;
    yt_rsc_1_0_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_1_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_2_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_3_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_4_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_5_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_6_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_7_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_8_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_9_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_10_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_11_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_12_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_13_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_14_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_15_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_16_i_clkr_en_d : OUT STD_LOGIC;
    yt_rsc_1_16_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_17_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_18_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_19_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_20_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_21_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_22_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_23_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_24_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_25_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_26_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_27_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_28_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_29_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_30_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_31_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_2_0_i_clkr_en_d : OUT STD_LOGIC;
    yt_rsc_2_0_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_2_1_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_2_2_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_2_3_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_2_4_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_2_5_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_2_6_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_2_7_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_2_8_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_2_9_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_2_10_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_2_11_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_2_12_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_2_13_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_2_14_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_2_15_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_2_16_i_clkr_en_d : OUT STD_LOGIC;
    yt_rsc_2_16_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_2_17_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_2_18_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_2_19_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_2_20_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_2_21_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_2_22_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_2_23_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_2_24_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_2_25_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_2_26_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_2_27_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_2_28_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_2_29_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_2_30_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_2_31_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_3_0_i_clkr_en_d : OUT STD_LOGIC;
    yt_rsc_3_0_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_3_1_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_3_2_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_3_3_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_3_4_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_3_5_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_3_6_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_3_7_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_3_8_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_3_9_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_3_10_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_3_11_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_3_12_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_3_13_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_3_14_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_3_15_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_3_16_i_clkr_en_d : OUT STD_LOGIC;
    yt_rsc_3_16_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_3_17_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_3_18_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_3_19_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_3_20_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_3_21_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_3_22_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_3_23_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_3_24_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_3_25_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_3_26_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_3_27_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_3_28_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_3_29_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_3_30_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_3_31_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_4_0_i_clkr_en_d : OUT STD_LOGIC;
    yt_rsc_4_0_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_4_1_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_4_2_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_4_3_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_4_4_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_4_5_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_4_6_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_4_7_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_4_8_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_4_9_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_4_10_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_4_11_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_4_12_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_4_13_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_4_14_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_4_15_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_4_16_i_clkr_en_d : OUT STD_LOGIC;
    yt_rsc_4_16_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_4_17_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_4_18_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_4_19_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_4_20_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_4_21_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_4_22_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_4_23_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_4_24_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_4_25_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_4_26_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_4_27_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_4_28_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_4_29_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_4_30_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_4_31_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_5_0_i_clkr_en_d : OUT STD_LOGIC;
    yt_rsc_5_0_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_5_1_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_5_2_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_5_3_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_5_4_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_5_5_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_5_6_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_5_7_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_5_8_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_5_9_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_5_10_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_5_11_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_5_12_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_5_13_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_5_14_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_5_15_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_5_16_i_clkr_en_d : OUT STD_LOGIC;
    yt_rsc_5_16_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_5_17_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_5_18_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_5_19_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_5_20_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_5_21_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_5_22_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_5_23_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_5_24_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_5_25_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_5_26_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_5_27_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_5_28_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_5_29_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_5_30_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_5_31_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_6_0_i_clkr_en_d : OUT STD_LOGIC;
    yt_rsc_6_0_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_6_1_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_6_2_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_6_3_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_6_4_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_6_5_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_6_6_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_6_7_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_6_8_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_6_9_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_6_10_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_6_11_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_6_12_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_6_13_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_6_14_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_6_15_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_6_16_i_clkr_en_d : OUT STD_LOGIC;
    yt_rsc_6_16_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_6_17_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_6_18_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_6_19_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_6_20_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_6_21_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_6_22_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_6_23_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_6_24_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_6_25_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_6_26_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_6_27_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_6_28_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_6_29_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_6_30_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_6_31_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_7_0_i_clkr_en_d : OUT STD_LOGIC;
    yt_rsc_7_0_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_7_1_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_7_2_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_7_3_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_7_4_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_7_5_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_7_6_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_7_7_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_7_8_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_7_9_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_7_10_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_7_11_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_7_12_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_7_13_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_7_14_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_7_15_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_7_16_i_clkr_en_d : OUT STD_LOGIC;
    yt_rsc_7_16_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_7_17_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_7_18_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_7_19_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_7_20_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_7_21_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_7_22_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_7_23_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_7_24_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_7_25_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_7_26_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_7_27_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_7_28_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_7_29_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_7_30_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_7_31_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_0_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_1_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_2_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_3_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_4_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_5_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_6_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_7_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_8_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_9_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_10_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_11_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_12_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_13_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_14_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_15_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_16_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_17_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_18_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_19_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_20_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_21_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_22_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_23_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_24_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_25_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_26_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_27_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_28_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_29_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_30_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_31_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_0_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_1_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_2_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_3_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_4_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_5_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_6_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_7_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_8_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_9_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_10_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_11_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_12_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_13_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_14_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_15_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_16_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_17_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_18_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_19_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_20_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_21_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_22_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_23_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_24_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_25_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_26_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_27_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_28_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_29_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_30_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_31_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_2_0_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_2_1_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_2_2_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_2_3_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_2_4_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_2_5_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_2_6_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_2_7_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_2_8_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_2_9_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_2_10_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_2_11_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_2_12_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_2_13_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_2_14_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_2_15_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_2_16_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_2_17_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_2_18_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_2_19_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_2_20_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_2_21_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_2_22_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_2_23_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_2_24_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_2_25_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_2_26_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_2_27_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_2_28_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_2_29_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_2_30_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_2_31_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_3_0_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_3_1_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_3_2_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_3_3_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_3_4_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_3_5_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_3_6_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_3_7_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_3_8_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_3_9_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_3_10_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_3_11_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_3_12_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_3_13_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_3_14_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_3_15_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_3_16_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_3_17_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_3_18_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_3_19_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_3_20_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_3_21_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_3_22_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_3_23_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_3_24_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_3_25_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_3_26_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_3_27_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_3_28_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_3_29_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_3_30_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_3_31_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_0_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_1_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_2_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_3_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_4_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_5_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_6_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_7_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_8_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_9_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_10_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_11_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_12_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_13_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_14_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_15_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_16_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_17_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_18_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_19_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_20_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_21_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_22_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_23_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_24_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_25_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_26_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_27_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_28_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_29_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_30_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_31_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_5_0_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_5_1_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_5_2_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_5_3_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_5_4_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_5_5_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_5_6_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_5_7_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_5_8_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_5_9_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_5_10_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_5_11_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_5_12_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_5_13_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_5_14_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_5_15_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_5_16_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_5_17_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_5_18_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_5_19_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_5_20_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_5_21_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_5_22_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_5_23_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_5_24_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_5_25_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_5_26_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_5_27_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_5_28_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_5_29_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_5_30_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_5_31_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_6_0_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_6_1_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_6_2_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_6_3_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_6_4_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_6_5_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_6_6_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_6_7_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_6_8_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_6_9_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_6_10_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_6_11_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_6_12_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_6_13_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_6_14_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_6_15_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_6_16_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_6_17_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_6_18_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_6_19_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_6_20_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_6_21_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_6_22_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_6_23_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_6_24_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_6_25_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_6_26_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_6_27_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_6_28_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_6_29_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_6_30_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_6_31_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_7_0_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_7_1_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_7_2_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_7_3_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_7_4_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_7_5_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_7_6_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_7_7_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_7_8_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_7_9_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_7_10_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_7_11_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_7_12_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_7_13_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_7_14_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_7_15_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_7_16_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_7_17_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_7_18_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_7_19_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_7_20_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_7_21_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_7_22_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_7_23_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_7_24_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_7_25_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_7_26_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_7_27_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_7_28_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_7_29_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_7_30_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_7_31_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_0_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
        DOWNTO 0);
    twiddle_rsc_0_1_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_1_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
        DOWNTO 0);
    twiddle_rsc_0_2_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_2_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
        DOWNTO 0);
    twiddle_rsc_0_3_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_3_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
        DOWNTO 0);
    twiddle_rsc_0_4_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_4_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
        DOWNTO 0);
    twiddle_rsc_0_5_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_5_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
        DOWNTO 0);
    twiddle_rsc_0_6_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_6_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
        DOWNTO 0);
    twiddle_rsc_0_7_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_7_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
        DOWNTO 0);
    twiddle_rsc_0_8_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_8_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
        DOWNTO 0);
    twiddle_rsc_0_9_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_9_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
        DOWNTO 0);
    twiddle_rsc_0_10_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_10_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
        DOWNTO 0);
    twiddle_rsc_0_11_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_11_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
        DOWNTO 0);
    twiddle_rsc_0_12_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_12_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
        DOWNTO 0);
    twiddle_rsc_0_13_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_13_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
        DOWNTO 0);
    twiddle_rsc_0_14_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_14_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
        DOWNTO 0);
    twiddle_rsc_0_15_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_15_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
        DOWNTO 0);
    twiddle_h_rsc_0_0_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_h_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
        DOWNTO 0);
    twiddle_h_rsc_0_1_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_1_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_h_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
        DOWNTO 0);
    twiddle_h_rsc_0_2_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_2_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_h_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
        DOWNTO 0);
    twiddle_h_rsc_0_3_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_3_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_h_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
        DOWNTO 0);
    twiddle_h_rsc_0_4_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_4_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_h_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
        DOWNTO 0);
    twiddle_h_rsc_0_5_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_5_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_h_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
        DOWNTO 0);
    twiddle_h_rsc_0_6_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_6_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_h_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
        DOWNTO 0);
    twiddle_h_rsc_0_7_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_7_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_h_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
        DOWNTO 0);
    twiddle_h_rsc_0_8_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_8_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_h_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
        DOWNTO 0);
    twiddle_h_rsc_0_9_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_9_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_h_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
        DOWNTO 0);
    twiddle_h_rsc_0_10_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_10_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_h_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    twiddle_h_rsc_0_11_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_11_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_h_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    twiddle_h_rsc_0_12_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_12_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_h_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    twiddle_h_rsc_0_13_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_13_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_h_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    twiddle_h_rsc_0_14_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_14_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_h_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    twiddle_h_rsc_0_15_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_15_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_h_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    yt_rsc_0_0_i_d_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_0_i_radr_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    yt_rsc_0_0_i_wadr_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    yt_rsc_0_0_i_we_d_pff : OUT STD_LOGIC;
    yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_pff : OUT STD_LOGIC;
    yt_rsc_0_1_i_d_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_1_i_wadr_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    yt_rsc_0_2_i_d_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_2_i_wadr_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    yt_rsc_0_3_i_d_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_3_i_wadr_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    yt_rsc_0_4_i_d_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_4_i_wadr_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    yt_rsc_0_5_i_d_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_5_i_wadr_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    yt_rsc_0_6_i_d_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_6_i_wadr_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    yt_rsc_0_7_i_d_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_8_i_d_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_9_i_d_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_10_i_d_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_10_i_wadr_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    yt_rsc_0_11_i_d_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_11_i_wadr_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    yt_rsc_0_12_i_d_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_13_i_d_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_14_i_d_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_15_i_d_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_16_i_we_d_pff : OUT STD_LOGIC;
    yt_rsc_1_0_i_we_d_pff : OUT STD_LOGIC;
    yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_pff : OUT STD_LOGIC;
    yt_rsc_1_16_i_we_d_pff : OUT STD_LOGIC;
    yt_rsc_2_0_i_we_d_pff : OUT STD_LOGIC;
    yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_pff : OUT STD_LOGIC;
    yt_rsc_2_16_i_we_d_pff : OUT STD_LOGIC;
    yt_rsc_3_0_i_we_d_pff : OUT STD_LOGIC;
    yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_pff : OUT STD_LOGIC;
    yt_rsc_3_16_i_we_d_pff : OUT STD_LOGIC;
    yt_rsc_4_0_i_d_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_4_0_i_wadr_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    yt_rsc_4_0_i_we_d_pff : OUT STD_LOGIC;
    yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_pff : OUT STD_LOGIC;
    yt_rsc_4_1_i_d_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_4_1_i_wadr_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    yt_rsc_4_2_i_d_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_4_2_i_wadr_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    yt_rsc_4_3_i_d_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_4_3_i_wadr_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    yt_rsc_4_4_i_d_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_4_4_i_wadr_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    yt_rsc_4_5_i_d_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_4_5_i_wadr_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    yt_rsc_4_6_i_d_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_4_6_i_wadr_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    yt_rsc_4_7_i_d_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_4_8_i_d_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_4_9_i_d_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_4_9_i_wadr_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    yt_rsc_4_10_i_d_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_4_10_i_wadr_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    yt_rsc_4_11_i_d_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_4_11_i_wadr_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    yt_rsc_4_12_i_d_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_4_13_i_d_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_4_14_i_d_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_4_15_i_d_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_4_16_i_we_d_pff : OUT STD_LOGIC;
    yt_rsc_5_0_i_we_d_pff : OUT STD_LOGIC;
    yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_pff : OUT STD_LOGIC;
    yt_rsc_5_16_i_we_d_pff : OUT STD_LOGIC;
    yt_rsc_6_0_i_we_d_pff : OUT STD_LOGIC;
    yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_pff : OUT STD_LOGIC;
    yt_rsc_6_16_i_we_d_pff : OUT STD_LOGIC;
    yt_rsc_7_0_i_we_d_pff : OUT STD_LOGIC;
    yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_pff : OUT STD_LOGIC;
    yt_rsc_7_16_i_we_d_pff : OUT STD_LOGIC;
    xt_rsc_0_0_i_adra_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_0_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_0_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff : OUT STD_LOGIC;
    xt_rsc_0_1_i_adra_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_1_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_2_i_adra_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_2_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_3_i_adra_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_3_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_4_i_adra_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_4_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_5_i_adra_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_5_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_6_i_adra_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_6_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_7_i_adra_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_7_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_8_i_adra_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_8_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_9_i_adra_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_9_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_10_i_adra_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_10_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_11_i_adra_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_11_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_12_i_adra_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_12_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_13_i_adra_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_13_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_14_i_adra_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_14_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_15_i_adra_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_15_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_16_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_1_0_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff : OUT STD_LOGIC;
    xt_rsc_1_16_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_2_0_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff : OUT STD_LOGIC;
    xt_rsc_2_16_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_3_0_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff : OUT STD_LOGIC;
    xt_rsc_3_16_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_4_0_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff : OUT STD_LOGIC;
    xt_rsc_4_1_i_adra_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_4_1_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_2_i_adra_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_4_2_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_3_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_4_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_5_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_6_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_7_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_8_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_9_i_adra_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_4_9_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_10_i_adra_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_4_10_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_11_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_12_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_13_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_14_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_15_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff : OUT STD_LOGIC;
    xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff : OUT STD_LOGIC;
    xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff : OUT STD_LOGIC
  );
END peaseNTT_core;

ARCHITECTURE v14 OF peaseNTT_core IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';

  -- Interconnect Declarations
  SIGNAL p_rsci_idat : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_en : STD_LOGIC;
  SIGNAL mult_t_mul_cmp_z : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_1_z : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_2_z : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_3_z : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_4_z : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_5_z : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_6_z : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_7_z : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_8_z : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_9_z : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_10_z : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_11_z : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_12_z : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_13_z : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_14_z : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_15_z : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_1_en : STD_LOGIC;
  SIGNAL mult_z_mul_cmp_1_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_2_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_3_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_4_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_5_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_6_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_7_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_8_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_9_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_10_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_11_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_12_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_13_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_14_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_15_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_16_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_17_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_18_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_19_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_20_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_21_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_22_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_23_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_24_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_25_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_26_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_27_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_28_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_29_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_30_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_31_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL fsm_output : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL INNER_LOOP4_nor_tmp : STD_LOGIC;
  SIGNAL or_dcpl : STD_LOGIC;
  SIGNAL or_dcpl_2 : STD_LOGIC;
  SIGNAL or_dcpl_8 : STD_LOGIC;
  SIGNAL or_dcpl_10 : STD_LOGIC;
  SIGNAL or_dcpl_12 : STD_LOGIC;
  SIGNAL or_dcpl_19 : STD_LOGIC;
  SIGNAL or_dcpl_22 : STD_LOGIC;
  SIGNAL or_dcpl_25 : STD_LOGIC;
  SIGNAL or_dcpl_30 : STD_LOGIC;
  SIGNAL or_dcpl_33 : STD_LOGIC;
  SIGNAL or_dcpl_36 : STD_LOGIC;
  SIGNAL or_dcpl_63 : STD_LOGIC;
  SIGNAL or_dcpl_70 : STD_LOGIC;
  SIGNAL or_dcpl_72 : STD_LOGIC;
  SIGNAL or_dcpl_76 : STD_LOGIC;
  SIGNAL or_dcpl_78 : STD_LOGIC;
  SIGNAL or_dcpl_80 : STD_LOGIC;
  SIGNAL or_dcpl_82 : STD_LOGIC;
  SIGNAL or_dcpl_88 : STD_LOGIC;
  SIGNAL or_dcpl_89 : STD_LOGIC;
  SIGNAL or_dcpl_94 : STD_LOGIC;
  SIGNAL or_dcpl_105 : STD_LOGIC;
  SIGNAL or_dcpl_107 : STD_LOGIC;
  SIGNAL or_dcpl_109 : STD_LOGIC;
  SIGNAL or_dcpl_111 : STD_LOGIC;
  SIGNAL or_dcpl_116 : STD_LOGIC;
  SIGNAL or_dcpl_117 : STD_LOGIC;
  SIGNAL or_dcpl_119 : STD_LOGIC;
  SIGNAL or_dcpl_121 : STD_LOGIC;
  SIGNAL or_dcpl_125 : STD_LOGIC;
  SIGNAL or_dcpl_133 : STD_LOGIC;
  SIGNAL or_dcpl_135 : STD_LOGIC;
  SIGNAL or_dcpl_139 : STD_LOGIC;
  SIGNAL or_dcpl_141 : STD_LOGIC;
  SIGNAL or_dcpl_146 : STD_LOGIC;
  SIGNAL or_dcpl_148 : STD_LOGIC;
  SIGNAL or_dcpl_150 : STD_LOGIC;
  SIGNAL or_dcpl_152 : STD_LOGIC;
  SIGNAL or_dcpl_161 : STD_LOGIC;
  SIGNAL or_dcpl_163 : STD_LOGIC;
  SIGNAL or_dcpl_165 : STD_LOGIC;
  SIGNAL or_dcpl_167 : STD_LOGIC;
  SIGNAL or_dcpl_171 : STD_LOGIC;
  SIGNAL or_dcpl_173 : STD_LOGIC;
  SIGNAL or_dcpl_180 : STD_LOGIC;
  SIGNAL or_dcpl_181 : STD_LOGIC;
  SIGNAL or_dcpl_185 : STD_LOGIC;
  SIGNAL or_dcpl_187 : STD_LOGIC;
  SIGNAL or_dcpl_189 : STD_LOGIC;
  SIGNAL or_dcpl_197 : STD_LOGIC;
  SIGNAL or_dcpl_199 : STD_LOGIC;
  SIGNAL or_dcpl_201 : STD_LOGIC;
  SIGNAL or_dcpl_203 : STD_LOGIC;
  SIGNAL or_dcpl_205 : STD_LOGIC;
  SIGNAL or_dcpl_207 : STD_LOGIC;
  SIGNAL or_dcpl_210 : STD_LOGIC;
  SIGNAL or_dcpl_215 : STD_LOGIC;
  SIGNAL or_dcpl_218 : STD_LOGIC;
  SIGNAL or_dcpl_220 : STD_LOGIC;
  SIGNAL or_dcpl_224 : STD_LOGIC;
  SIGNAL or_dcpl_234 : STD_LOGIC;
  SIGNAL or_dcpl_238 : STD_LOGIC;
  SIGNAL or_dcpl_242 : STD_LOGIC;
  SIGNAL or_dcpl_246 : STD_LOGIC;
  SIGNAL or_dcpl_274 : STD_LOGIC;
  SIGNAL and_dcpl_62 : STD_LOGIC;
  SIGNAL or_tmp_26 : STD_LOGIC;
  SIGNAL or_tmp_29 : STD_LOGIC;
  SIGNAL mux_tmp : STD_LOGIC;
  SIGNAL or_tmp_35 : STD_LOGIC;
  SIGNAL not_tmp_25 : STD_LOGIC;
  SIGNAL or_tmp_38 : STD_LOGIC;
  SIGNAL or_tmp_40 : STD_LOGIC;
  SIGNAL not_tmp_29 : STD_LOGIC;
  SIGNAL and_dcpl_66 : STD_LOGIC;
  SIGNAL and_dcpl_67 : STD_LOGIC;
  SIGNAL and_dcpl_68 : STD_LOGIC;
  SIGNAL and_dcpl_69 : STD_LOGIC;
  SIGNAL and_dcpl_70 : STD_LOGIC;
  SIGNAL and_dcpl_73 : STD_LOGIC;
  SIGNAL and_dcpl_76 : STD_LOGIC;
  SIGNAL nor_tmp_1 : STD_LOGIC;
  SIGNAL or_tmp_48 : STD_LOGIC;
  SIGNAL or_tmp_50 : STD_LOGIC;
  SIGNAL mux_tmp_7 : STD_LOGIC;
  SIGNAL or_tmp_53 : STD_LOGIC;
  SIGNAL or_tmp_55 : STD_LOGIC;
  SIGNAL not_tmp_50 : STD_LOGIC;
  SIGNAL and_dcpl_78 : STD_LOGIC;
  SIGNAL and_dcpl_79 : STD_LOGIC;
  SIGNAL or_tmp_64 : STD_LOGIC;
  SIGNAL and_dcpl_81 : STD_LOGIC;
  SIGNAL and_dcpl_82 : STD_LOGIC;
  SIGNAL and_dcpl_83 : STD_LOGIC;
  SIGNAL or_tmp_72 : STD_LOGIC;
  SIGNAL and_dcpl_89 : STD_LOGIC;
  SIGNAL or_tmp_75 : STD_LOGIC;
  SIGNAL or_tmp_77 : STD_LOGIC;
  SIGNAL mux_tmp_22 : STD_LOGIC;
  SIGNAL nor_tmp_6 : STD_LOGIC;
  SIGNAL or_tmp_82 : STD_LOGIC;
  SIGNAL nor_tmp_10 : STD_LOGIC;
  SIGNAL or_tmp_84 : STD_LOGIC;
  SIGNAL or_tmp_86 : STD_LOGIC;
  SIGNAL not_tmp_67 : STD_LOGIC;
  SIGNAL not_tmp_69 : STD_LOGIC;
  SIGNAL or_tmp_90 : STD_LOGIC;
  SIGNAL and_dcpl_92 : STD_LOGIC;
  SIGNAL and_dcpl_93 : STD_LOGIC;
  SIGNAL nor_tmp_14 : STD_LOGIC;
  SIGNAL nor_tmp_15 : STD_LOGIC;
  SIGNAL or_tmp_93 : STD_LOGIC;
  SIGNAL or_tmp_94 : STD_LOGIC;
  SIGNAL nor_tmp_19 : STD_LOGIC;
  SIGNAL and_dcpl_96 : STD_LOGIC;
  SIGNAL or_tmp_99 : STD_LOGIC;
  SIGNAL or_tmp_102 : STD_LOGIC;
  SIGNAL or_tmp_104 : STD_LOGIC;
  SIGNAL and_dcpl_99 : STD_LOGIC;
  SIGNAL nor_tmp_22 : STD_LOGIC;
  SIGNAL or_tmp_112 : STD_LOGIC;
  SIGNAL not_tmp_87 : STD_LOGIC;
  SIGNAL mux_tmp_45 : STD_LOGIC;
  SIGNAL or_tmp_120 : STD_LOGIC;
  SIGNAL or_tmp_122 : STD_LOGIC;
  SIGNAL not_tmp_91 : STD_LOGIC;
  SIGNAL mux_tmp_50 : STD_LOGIC;
  SIGNAL and_dcpl_101 : STD_LOGIC;
  SIGNAL and_dcpl_102 : STD_LOGIC;
  SIGNAL and_dcpl_104 : STD_LOGIC;
  SIGNAL and_dcpl_105 : STD_LOGIC;
  SIGNAL and_dcpl_107 : STD_LOGIC;
  SIGNAL nor_tmp_25 : STD_LOGIC;
  SIGNAL mux_tmp_53 : STD_LOGIC;
  SIGNAL mux_tmp_56 : STD_LOGIC;
  SIGNAL or_tmp_133 : STD_LOGIC;
  SIGNAL and_dcpl_112 : STD_LOGIC;
  SIGNAL and_dcpl_114 : STD_LOGIC;
  SIGNAL and_dcpl_116 : STD_LOGIC;
  SIGNAL and_dcpl_123 : STD_LOGIC;
  SIGNAL mux_tmp_70 : STD_LOGIC;
  SIGNAL nor_tmp_32 : STD_LOGIC;
  SIGNAL or_tmp_153 : STD_LOGIC;
  SIGNAL not_tmp_115 : STD_LOGIC;
  SIGNAL or_tmp_156 : STD_LOGIC;
  SIGNAL and_dcpl_125 : STD_LOGIC;
  SIGNAL nor_tmp_36 : STD_LOGIC;
  SIGNAL mux_tmp_78 : STD_LOGIC;
  SIGNAL or_tmp_160 : STD_LOGIC;
  SIGNAL nor_tmp_43 : STD_LOGIC;
  SIGNAL nor_tmp_45 : STD_LOGIC;
  SIGNAL nor_tmp_46 : STD_LOGIC;
  SIGNAL and_dcpl_135 : STD_LOGIC;
  SIGNAL and_dcpl_138 : STD_LOGIC;
  SIGNAL and_dcpl_141 : STD_LOGIC;
  SIGNAL and_dcpl_145 : STD_LOGIC;
  SIGNAL and_dcpl_147 : STD_LOGIC;
  SIGNAL and_dcpl_150 : STD_LOGIC;
  SIGNAL and_dcpl_152 : STD_LOGIC;
  SIGNAL and_dcpl_154 : STD_LOGIC;
  SIGNAL and_dcpl_161 : STD_LOGIC;
  SIGNAL and_dcpl_163 : STD_LOGIC;
  SIGNAL and_dcpl_167 : STD_LOGIC;
  SIGNAL and_dcpl_169 : STD_LOGIC;
  SIGNAL or_dcpl_298 : STD_LOGIC;
  SIGNAL or_dcpl_300 : STD_LOGIC;
  SIGNAL and_dcpl_173 : STD_LOGIC;
  SIGNAL and_dcpl_175 : STD_LOGIC;
  SIGNAL and_dcpl_176 : STD_LOGIC;
  SIGNAL or_dcpl_315 : STD_LOGIC;
  SIGNAL and_dcpl_239 : STD_LOGIC;
  SIGNAL or_dcpl_353 : STD_LOGIC;
  SIGNAL or_dcpl_361 : STD_LOGIC;
  SIGNAL or_tmp_3231 : STD_LOGIC;
  SIGNAL or_tmp_3239 : STD_LOGIC;
  SIGNAL or_tmp_3242 : STD_LOGIC;
  SIGNAL or_tmp_3250 : STD_LOGIC;
  SIGNAL or_tmp_3252 : STD_LOGIC;
  SIGNAL or_tmp_3269 : STD_LOGIC;
  SIGNAL or_tmp_3279 : STD_LOGIC;
  SIGNAL or_tmp_3345 : STD_LOGIC;
  SIGNAL or_tmp_3354 : STD_LOGIC;
  SIGNAL or_tmp_3597 : STD_LOGIC;
  SIGNAL or_tmp_3600 : STD_LOGIC;
  SIGNAL or_tmp_3650 : STD_LOGIC;
  SIGNAL or_tmp_3666 : STD_LOGIC;
  SIGNAL or_tmp_3717 : STD_LOGIC;
  SIGNAL or_tmp_3723 : STD_LOGIC;
  SIGNAL or_tmp_3732 : STD_LOGIC;
  SIGNAL or_tmp_3755 : STD_LOGIC;
  SIGNAL or_tmp_3842 : STD_LOGIC;
  SIGNAL and_344_cse : STD_LOGIC;
  SIGNAL and_346_cse : STD_LOGIC;
  SIGNAL and_715_cse : STD_LOGIC;
  SIGNAL and_717_cse : STD_LOGIC;
  SIGNAL and_1022_cse : STD_LOGIC;
  SIGNAL and_1024_cse : STD_LOGIC;
  SIGNAL and_1329_cse : STD_LOGIC;
  SIGNAL and_1331_cse : STD_LOGIC;
  SIGNAL and_1636_cse : STD_LOGIC;
  SIGNAL and_1638_cse : STD_LOGIC;
  SIGNAL and_2007_cse : STD_LOGIC;
  SIGNAL and_2009_cse : STD_LOGIC;
  SIGNAL and_2314_cse : STD_LOGIC;
  SIGNAL and_2316_cse : STD_LOGIC;
  SIGNAL and_2621_cse : STD_LOGIC;
  SIGNAL and_2623_cse : STD_LOGIC;
  SIGNAL and_6834_cse : STD_LOGIC;
  SIGNAL and_6843_cse : STD_LOGIC;
  SIGNAL and_6852_cse : STD_LOGIC;
  SIGNAL and_7090_cse : STD_LOGIC;
  SIGNAL and_7109_cse : STD_LOGIC;
  SIGNAL and_7115_cse : STD_LOGIC;
  SIGNAL and_7153_cse : STD_LOGIC;
  SIGNAL and_7173_cse : STD_LOGIC;
  SIGNAL INNER_LOOP4_r_11_4_sva_6_0 : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL INNER_LOOP3_r_11_4_sva_6_0 : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL INNER_LOOP2_r_11_4_sva_6_0 : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_11_4_sva_6_0 : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL butterFly1_15_conc_2_itm_2_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL c_1_sva : STD_LOGIC;
  SIGNAL INNER_LOOP1_stage_0 : STD_LOGIC;
  SIGNAL butterFly1_15_conc_2_itm_3_0 : STD_LOGIC;
  SIGNAL butterFly1_15_conc_2_itm_8_0 : STD_LOGIC;
  SIGNAL butterFly1_15_conc_2_itm_5_0 : STD_LOGIC;
  SIGNAL butterFly1_15_conc_2_itm_4_0 : STD_LOGIC;
  SIGNAL butterFly1_15_conc_2_itm_2_0 : STD_LOGIC;
  SIGNAL butterFly2_15_conc_itm_10_2_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL butterFly2_15_conc_2_itm_9_2_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL butterFly1_15_f1_equal_tmp_1_1 : STD_LOGIC;
  SIGNAL butterFly1_15_conc_2_itm_0 : STD_LOGIC;
  SIGNAL butterFly1_15_f1_equal_tmp_2_1 : STD_LOGIC;
  SIGNAL butterFly1_15_conc_2_itm_1_0 : STD_LOGIC;
  SIGNAL butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1 : STD_LOGIC_VECTOR (2
      DOWNTO 0);
  SIGNAL butterFly2_15_conc_2_itm_6_2_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL butterFly1_15_conc_2_itm_9_2_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL butterFly1_15_conc_2_itm_9_0 : STD_LOGIC;
  SIGNAL INNER_LOOP1_stage_0_10 : STD_LOGIC;
  SIGNAL butterFly2_15_conc_2_itm_7_0 : STD_LOGIC;
  SIGNAL INNER_LOOP1_stage_0_11 : STD_LOGIC;
  SIGNAL INNER_LOOP2_stage_0_10 : STD_LOGIC;
  SIGNAL butterFly2_15_conc_2_itm_8_2_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL butterFly2_15_conc_2_itm_8_0 : STD_LOGIC;
  SIGNAL butterFly1_15_conc_2_itm_8_2_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL butterFly2_15_conc_2_itm_5_0 : STD_LOGIC;
  SIGNAL operator_20_false_acc_cse_sva : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL operator_33_true_3_lshift_psp_1_0_sva : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL INNER_LOOP1_stage_0_3 : STD_LOGIC;
  SIGNAL INNER_LOOP1_stage_0_2 : STD_LOGIC;
  SIGNAL butterFly2_15_conc_2_itm_0 : STD_LOGIC;
  SIGNAL butterFly2_15_conc_2_itm_1_0 : STD_LOGIC;
  SIGNAL butterFly2_15_conc_2_itm_2_0 : STD_LOGIC;
  SIGNAL butterFly2_15_conc_2_itm_3_0 : STD_LOGIC;
  SIGNAL butterFly1_15_conc_2_itm_4_2_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL p_sva : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_15_and_ssc : STD_LOGIC;
  SIGNAL butterFly1_15_and_ssc_2 : STD_LOGIC;
  SIGNAL butterFly1_14_and_ssc : STD_LOGIC;
  SIGNAL butterFly1_14_and_ssc_2 : STD_LOGIC;
  SIGNAL butterFly1_14_and_ssc_3 : STD_LOGIC;
  SIGNAL butterFly1_13_and_ssc : STD_LOGIC;
  SIGNAL butterFly1_13_and_ssc_2 : STD_LOGIC;
  SIGNAL butterFly1_13_and_ssc_3 : STD_LOGIC;
  SIGNAL butterFly1_12_and_ssc : STD_LOGIC;
  SIGNAL butterFly1_12_and_ssc_2 : STD_LOGIC;
  SIGNAL butterFly1_12_and_ssc_3 : STD_LOGIC;
  SIGNAL butterFly1_11_and_ssc : STD_LOGIC;
  SIGNAL butterFly1_11_and_ssc_2 : STD_LOGIC;
  SIGNAL butterFly1_11_and_ssc_3 : STD_LOGIC;
  SIGNAL butterFly1_10_and_ssc : STD_LOGIC;
  SIGNAL butterFly1_10_and_ssc_2 : STD_LOGIC;
  SIGNAL butterFly1_10_and_ssc_3 : STD_LOGIC;
  SIGNAL butterFly1_9_and_ssc : STD_LOGIC;
  SIGNAL butterFly1_9_and_ssc_2 : STD_LOGIC;
  SIGNAL butterFly1_9_and_ssc_3 : STD_LOGIC;
  SIGNAL butterFly1_8_and_ssc : STD_LOGIC;
  SIGNAL butterFly1_8_and_ssc_2 : STD_LOGIC;
  SIGNAL butterFly1_8_and_ssc_3 : STD_LOGIC;
  SIGNAL butterFly1_7_and_ssc : STD_LOGIC;
  SIGNAL butterFly1_7_and_ssc_2 : STD_LOGIC;
  SIGNAL butterFly1_7_and_ssc_3 : STD_LOGIC;
  SIGNAL butterFly1_6_and_ssc : STD_LOGIC;
  SIGNAL butterFly1_6_and_ssc_2 : STD_LOGIC;
  SIGNAL butterFly1_6_and_ssc_3 : STD_LOGIC;
  SIGNAL butterFly1_5_and_ssc : STD_LOGIC;
  SIGNAL butterFly1_5_and_ssc_2 : STD_LOGIC;
  SIGNAL butterFly1_5_and_ssc_3 : STD_LOGIC;
  SIGNAL butterFly1_4_and_ssc : STD_LOGIC;
  SIGNAL butterFly1_4_and_ssc_2 : STD_LOGIC;
  SIGNAL butterFly1_4_and_ssc_3 : STD_LOGIC;
  SIGNAL butterFly1_3_and_ssc : STD_LOGIC;
  SIGNAL butterFly1_3_and_ssc_2 : STD_LOGIC;
  SIGNAL butterFly1_3_and_ssc_3 : STD_LOGIC;
  SIGNAL butterFly1_2_and_ssc : STD_LOGIC;
  SIGNAL butterFly1_2_and_ssc_2 : STD_LOGIC;
  SIGNAL butterFly1_2_and_ssc_3 : STD_LOGIC;
  SIGNAL butterFly1_1_and_ssc : STD_LOGIC;
  SIGNAL butterFly1_1_and_ssc_2 : STD_LOGIC;
  SIGNAL butterFly1_1_and_ssc_3 : STD_LOGIC;
  SIGNAL butterFly1_and_ssc : STD_LOGIC;
  SIGNAL butterFly1_and_ssc_2 : STD_LOGIC;
  SIGNAL reg_yt_rsc_0_0_cgo_cse : STD_LOGIC;
  SIGNAL reg_yt_rsc_0_16_cgo_cse : STD_LOGIC;
  SIGNAL reg_yt_rsc_1_0_cgo_cse : STD_LOGIC;
  SIGNAL reg_yt_rsc_1_16_cgo_cse : STD_LOGIC;
  SIGNAL reg_yt_rsc_2_0_cgo_cse : STD_LOGIC;
  SIGNAL reg_yt_rsc_2_16_cgo_cse : STD_LOGIC;
  SIGNAL reg_yt_rsc_3_0_cgo_cse : STD_LOGIC;
  SIGNAL reg_yt_rsc_3_16_cgo_cse : STD_LOGIC;
  SIGNAL reg_yt_rsc_4_0_cgo_cse : STD_LOGIC;
  SIGNAL reg_yt_rsc_4_16_cgo_cse : STD_LOGIC;
  SIGNAL reg_yt_rsc_5_0_cgo_cse : STD_LOGIC;
  SIGNAL reg_yt_rsc_5_16_cgo_cse : STD_LOGIC;
  SIGNAL reg_yt_rsc_6_0_cgo_cse : STD_LOGIC;
  SIGNAL reg_yt_rsc_6_16_cgo_cse : STD_LOGIC;
  SIGNAL reg_yt_rsc_7_0_cgo_cse : STD_LOGIC;
  SIGNAL reg_yt_rsc_7_16_cgo_cse : STD_LOGIC;
  SIGNAL reg_xt_rsc_triosy_7_31_obj_ld_cse : STD_LOGIC;
  SIGNAL reg_ensig_cgo_cse : STD_LOGIC;
  SIGNAL mult_15_t_and_49_cse : STD_LOGIC;
  SIGNAL mult_15_t_and_51_cse : STD_LOGIC;
  SIGNAL mult_15_t_and_53_cse : STD_LOGIC;
  SIGNAL mult_15_t_and_55_cse : STD_LOGIC;
  SIGNAL mult_15_t_and_44_cse : STD_LOGIC;
  SIGNAL mult_15_t_and_45_cse : STD_LOGIC;
  SIGNAL mult_15_t_and_46_cse : STD_LOGIC;
  SIGNAL mult_15_t_and_47_cse : STD_LOGIC;
  SIGNAL mult_15_t_and_48_cse : STD_LOGIC;
  SIGNAL mult_15_t_and_50_cse : STD_LOGIC;
  SIGNAL mult_15_t_and_52_cse : STD_LOGIC;
  SIGNAL mult_15_t_and_54_cse : STD_LOGIC;
  SIGNAL reg_ensig_cgo_17_cse : STD_LOGIC;
  SIGNAL or_383_cse : STD_LOGIC;
  SIGNAL or_398_cse : STD_LOGIC;
  SIGNAL nor_27_cse : STD_LOGIC;
  SIGNAL and_8912_cse : STD_LOGIC;
  SIGNAL butterFly2_16_f1_nor_1_cse : STD_LOGIC;
  SIGNAL nand_7_cse : STD_LOGIC;
  SIGNAL and_8932_cse : STD_LOGIC;
  SIGNAL and_8913_cse : STD_LOGIC;
  SIGNAL and_8919_cse : STD_LOGIC;
  SIGNAL butterFly2_f1_nor_cse : STD_LOGIC;
  SIGNAL butterFly1_f1_nor_cse : STD_LOGIC;
  SIGNAL or_329_cse : STD_LOGIC;
  SIGNAL or_412_cse : STD_LOGIC;
  SIGNAL nand_24_cse : STD_LOGIC;
  SIGNAL butterFly2_16_f1_butterFly2_16_f1_and_6_cse : STD_LOGIC;
  SIGNAL and_8941_cse : STD_LOGIC;
  SIGNAL mult_15_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_14_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_13_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_12_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_11_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_10_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_9_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_8_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_7_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_6_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_5_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_4_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_3_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_2_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_1_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly2_7_tw_nor_cse : STD_LOGIC;
  SIGNAL butterFly2_7_tw_nor_1_cse : STD_LOGIC;
  SIGNAL butterFly2_7_tw_nor_2_cse : STD_LOGIC;
  SIGNAL mult_15_t_or_9_cse : STD_LOGIC;
  SIGNAL mult_15_t_or_10_cse : STD_LOGIC;
  SIGNAL mult_15_t_or_11_cse : STD_LOGIC;
  SIGNAL mult_15_t_or_12_cse : STD_LOGIC;
  SIGNAL mult_15_t_and_41_cse : STD_LOGIC;
  SIGNAL mult_15_t_and_42_cse : STD_LOGIC;
  SIGNAL mult_15_t_and_43_cse : STD_LOGIC;
  SIGNAL mult_15_t_and_37_cse : STD_LOGIC;
  SIGNAL mult_15_t_and_38_cse : STD_LOGIC;
  SIGNAL mult_15_t_and_39_cse : STD_LOGIC;
  SIGNAL mult_15_t_and_30_cse : STD_LOGIC;
  SIGNAL mult_15_t_and_31_cse : STD_LOGIC;
  SIGNAL mult_15_t_and_32_cse : STD_LOGIC;
  SIGNAL mult_15_t_or_3_cse : STD_LOGIC;
  SIGNAL mult_15_t_and_40_cse : STD_LOGIC;
  SIGNAL mult_15_t_and_36_cse : STD_LOGIC;
  SIGNAL mult_15_t_and_29_cse : STD_LOGIC;
  SIGNAL mult_15_t_or_1_cse : STD_LOGIC;
  SIGNAL mult_15_t_or_cse : STD_LOGIC;
  SIGNAL or_553_rmff : STD_LOGIC;
  SIGNAL or_652_rmff : STD_LOGIC;
  SIGNAL or_718_rmff : STD_LOGIC;
  SIGNAL or_785_rmff : STD_LOGIC;
  SIGNAL or_851_rmff : STD_LOGIC;
  SIGNAL or_918_rmff : STD_LOGIC;
  SIGNAL or_984_rmff : STD_LOGIC;
  SIGNAL or_1051_rmff : STD_LOGIC;
  SIGNAL or_1117_rmff : STD_LOGIC;
  SIGNAL or_1216_rmff : STD_LOGIC;
  SIGNAL or_1282_rmff : STD_LOGIC;
  SIGNAL or_1349_rmff : STD_LOGIC;
  SIGNAL or_1415_rmff : STD_LOGIC;
  SIGNAL or_1482_rmff : STD_LOGIC;
  SIGNAL or_1548_rmff : STD_LOGIC;
  SIGNAL or_1615_rmff : STD_LOGIC;
  SIGNAL INNER_LOOP1_tw_h_mux1h_4_rmff : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL and_6824_rmff : STD_LOGIC;
  SIGNAL butterFly2_1_tw_butterFly2_1_tw_mux_rmff : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL or_3498_rmff : STD_LOGIC;
  SIGNAL or_3502_rmff : STD_LOGIC;
  SIGNAL or_3506_rmff : STD_LOGIC;
  SIGNAL or_3510_rmff : STD_LOGIC;
  SIGNAL or_3514_rmff : STD_LOGIC;
  SIGNAL or_3518_rmff : STD_LOGIC;
  SIGNAL or_3522_rmff : STD_LOGIC;
  SIGNAL and_6895_rmff : STD_LOGIC;
  SIGNAL or_3599_rmff : STD_LOGIC;
  SIGNAL or_3759_rmff : STD_LOGIC;
  SIGNAL mult_4_t_mux1h_1_rmff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_5_a_mx0w1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_5_a_mx0w4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_11_a_mx0w3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_71_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_31_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_10_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_8450_itm_9 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_8833_itm_8 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL modulo_add_1_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_11_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_8961_itm_9 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_9344_itm_8 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL modulo_add_23_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_12_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_9472_itm_9 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_9855_itm_8 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL modulo_add_24_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_13_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_10015_itm_9 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_10366_itm_8 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL modulo_add_25_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_14_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_10494_itm_9 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_10877_itm_8 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL modulo_add_26_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_15_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_11005_itm_9 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_11388_itm_8 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL modulo_add_27_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_11516_itm_9 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_11899_itm_8 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL modulo_add_28_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_29_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_30_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13560_itm_9 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13943_itm_8 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14071_itm_9 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14454_itm_8 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12538_itm_8 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13049_itm_8 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14582_itm_8 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15093_itm_8 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15604_itm_8 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16115_itm_8 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12027_itm_8 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13560_itm_8 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14071_itm_8 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12538_itm_5 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12921_itm_5 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13049_itm_6 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13432_itm_6 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9472_itm_9 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9855_itm_9 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15093_itm_1 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15476_itm_1 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15604_itm_2 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15987_itm_2 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16115_itm_3 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16498_itm_3 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12027_itm_4 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12410_itm_4 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13560_itm_7 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13943_itm_7 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL z_out : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_9 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_10 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_11 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_12 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_13 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_14 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_15 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_16 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_17 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_18 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_19 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_20 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_21 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_22 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_23 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_24 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_25 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_26 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_27 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_28 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_29 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_30 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_31 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_32 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_33 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_34 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_35 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_36 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_37 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_38 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_39 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_40 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_41 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_42 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_43 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_44 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_45 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_46 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_47 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_48 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_49 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_50 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_51 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_52 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_53 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_54 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_55 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_56 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_57 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_58 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_59 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_60 : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL z_out_61 : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL z_out_62 : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL z_out_68 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_69 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_70 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_72 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_73 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_74 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_76 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_77 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_78 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_80 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_81 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_82 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_84 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_85 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_86 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_88 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_89 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_90 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_92 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_93 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_94 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_96 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_97 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_98 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_100 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_101 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_102 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_104 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_105 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_106 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_108 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_109 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_111 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_112 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_113 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_114 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_115 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_116 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_117 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_118 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_119 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_120 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_121 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_122 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_123 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_124 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_125 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_126 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_127 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_128 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_129 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_130 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_131 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_132 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_133 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_134 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_135 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_136 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_137 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_138 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_139 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_140 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_141 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_142 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL operator_33_true_1_lshift_psp_9_4_sva : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL tmp_64_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_66_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_68_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_70_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_72_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_74_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_76_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_78_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_80_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_82_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_84_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_86_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_88_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_90_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_92_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_15_f1_equal_tmp_1 : STD_LOGIC;
  SIGNAL butterFly1_15_f1_equal_tmp_3_1 : STD_LOGIC;
  SIGNAL butterFly1_15_f1_equal_tmp_4_1 : STD_LOGIC;
  SIGNAL butterFly1_15_f1_equal_tmp_5_1 : STD_LOGIC;
  SIGNAL butterFly1_15_f1_equal_tmp_6_1 : STD_LOGIC;
  SIGNAL butterFly1_15_f1_equal_tmp_7_1 : STD_LOGIC;
  SIGNAL tmp_94_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_1_z_asn_itm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_1_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12027_itm_1 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12027_itm_2 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12027_itm_3 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12027_itm_5 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12027_itm_6 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12027_itm_7 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12410_itm_1 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12410_itm_2 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12410_itm_3 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12410_itm_5 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12410_itm_6 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12410_itm_7 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12538_itm_1 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12538_itm_2 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12538_itm_3 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12538_itm_4 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12538_itm_6 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12538_itm_7 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12921_itm_1 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12921_itm_2 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12921_itm_3 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12921_itm_4 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12921_itm_6 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12921_itm_7 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13049_itm_1 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13049_itm_2 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13049_itm_3 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13049_itm_4 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13049_itm_5 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13049_itm_7 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13432_itm_1 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13432_itm_2 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13432_itm_3 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13432_itm_4 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13432_itm_5 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13432_itm_7 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL mult_10_z_asn_itm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_10_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_10_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13560_itm_1 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13560_itm_2 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13560_itm_3 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13560_itm_4 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13560_itm_5 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13560_itm_6 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13943_itm_1 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13943_itm_2 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13943_itm_3 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13943_itm_4 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13943_itm_5 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13943_itm_6 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL mult_11_z_asn_itm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_11_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_11_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14071_itm_1 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14071_itm_2 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14071_itm_3 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14071_itm_4 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14071_itm_5 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14071_itm_6 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14071_itm_7 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14454_itm_1 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14454_itm_2 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14454_itm_3 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14454_itm_4 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14454_itm_5 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14454_itm_6 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14454_itm_7 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL mult_12_z_asn_itm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_12_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_12_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14582_itm_1 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14582_itm_2 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14582_itm_3 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14582_itm_4 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14582_itm_5 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14582_itm_6 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14582_itm_7 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14965_itm_1 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14965_itm_2 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14965_itm_3 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14965_itm_4 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14965_itm_5 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14965_itm_6 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14965_itm_7 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL mult_13_z_asn_itm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_13_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_13_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15093_itm_2 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15093_itm_3 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15093_itm_4 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15093_itm_5 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15093_itm_6 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15093_itm_7 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15476_itm_2 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15476_itm_3 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15476_itm_4 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15476_itm_5 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15476_itm_6 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15476_itm_7 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL mult_14_z_asn_itm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_14_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_14_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15604_itm_1 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15604_itm_3 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15604_itm_4 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15604_itm_5 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15604_itm_6 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15604_itm_7 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15987_itm_1 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15987_itm_3 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15987_itm_4 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15987_itm_5 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15987_itm_6 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15987_itm_7 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL mult_15_z_asn_itm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_15_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_15_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16115_itm_1 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16115_itm_2 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16115_itm_4 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16115_itm_5 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16115_itm_6 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16115_itm_7 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16498_itm_1 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16498_itm_2 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16498_itm_4 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16498_itm_5 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16498_itm_6 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16498_itm_7 : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL tmp_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_2_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_4_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_6_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_8_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_10_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_10_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_10_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_10_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_10_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_10_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_10_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_12_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_14_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_16_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_18_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_20_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_22_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_24_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_26_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_28_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_30_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_16_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_17_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_18_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9472_itm_3 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9472_itm_4 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9472_itm_5 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9472_itm_6 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9472_itm_7 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9472_itm_8 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9855_itm_1 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9855_itm_2 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9855_itm_3 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9855_itm_4 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9855_itm_5 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9855_itm_6 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9855_itm_7 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9855_itm_8 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL mult_19_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_20_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_21_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_22_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_23_z_asn_itm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_23_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_23_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_24_z_asn_itm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_24_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_24_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_25_z_asn_itm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_25_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_25_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_26_z_asn_itm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_26_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_27_z_asn_itm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_27_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_28_z_asn_itm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_28_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_29_z_asn_itm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_29_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_30_z_asn_itm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_30_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_31_z_asn_itm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_31_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_96_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_98_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_100_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_102_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_102_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_102_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_102_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_102_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_102_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_102_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_104_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_104_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_104_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_104_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_104_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_104_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_104_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_106_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_106_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_106_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_106_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_106_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_106_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_106_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_108_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_108_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_108_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_108_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_108_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_108_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_108_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_110_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_110_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_110_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_110_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_110_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_110_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_110_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_112_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_112_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_112_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_112_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_112_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_112_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_112_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_114_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_114_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_114_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_114_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_114_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_114_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_114_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_116_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_116_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_116_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_116_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_116_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_116_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_116_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_118_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_118_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_118_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_118_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_118_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_118_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_118_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_120_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_120_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_120_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_120_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_120_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_120_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_120_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_122_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_122_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_122_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_122_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_122_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_122_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_122_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_124_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_124_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_124_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_124_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_124_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_124_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_124_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly2_15_f1_equal_tmp_1 : STD_LOGIC;
  SIGNAL butterFly2_15_f1_equal_tmp_7_1 : STD_LOGIC;
  SIGNAL tmp_126_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_126_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_126_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_126_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_126_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_126_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_126_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly2_15_tw_equal_tmp_1 : STD_LOGIC;
  SIGNAL butterFly2_15_tw_equal_tmp_3_1 : STD_LOGIC;
  SIGNAL butterFly2_15_tw_equal_tmp_5_1 : STD_LOGIC;
  SIGNAL butterFly2_15_tw_equal_tmp_6_1 : STD_LOGIC;
  SIGNAL butterFly2_15_tw_equal_tmp_7_1 : STD_LOGIC;
  SIGNAL tmp_32_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_34_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_36_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_38_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_40_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_42_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_44_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_46_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_48_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_50_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_52_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_54_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_56_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_58_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_60_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_60_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_60_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_60_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_60_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_60_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_60_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_62_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_62_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_62_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_62_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_62_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_62_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_62_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_15_conc_2_itm_1_2_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL butterFly1_15_conc_2_itm_2_2_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL butterFly1_15_conc_2_itm_3_2_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL butterFly1_15_conc_2_itm_5_2_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL butterFly1_15_conc_2_itm_6_2_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL butterFly1_15_conc_2_itm_6_0 : STD_LOGIC;
  SIGNAL butterFly1_15_conc_2_itm_7_2_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL butterFly1_15_conc_2_itm_7_0 : STD_LOGIC;
  SIGNAL butterFly2_15_conc_2_itm_4_0 : STD_LOGIC;
  SIGNAL butterFly2_15_conc_2_itm_7_2_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL operator_33_true_3_lshift_psp_1_0_sva_mx0w5 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL mult_15_res_lpi_3_dfm_1_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_14_res_lpi_3_dfm_1_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_13_res_lpi_3_dfm_1_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_12_res_lpi_3_dfm_1_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_11_res_lpi_3_dfm_1_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_10_res_lpi_3_dfm_1_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_9_res_lpi_3_dfm_1_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_8_res_lpi_3_dfm_1_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_7_res_lpi_3_dfm_1_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_6_res_lpi_3_dfm_1_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_5_res_lpi_3_dfm_1_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_4_res_lpi_3_dfm_1_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_3_res_lpi_3_dfm_1_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_2_res_lpi_3_dfm_1_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_1_res_lpi_3_dfm_1_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_res_lpi_3_dfm_1_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL INNER_LOOP2_r_11_4_sva_6_0_mx1 : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL operator_33_true_2_lshift_psp_2_0_sva_mx0 : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL modulo_sub_31_qelse_and_ssc : STD_LOGIC;
  SIGNAL modulo_sub_31_qelse_and_ssc_1 : STD_LOGIC;
  SIGNAL reg_modulo_sub_31_qr_lpi_3_dfm_1_ftd : STD_LOGIC;
  SIGNAL reg_modulo_sub_31_qr_lpi_3_dfm_1_ftd_1 : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_30_qelse_and_ssc : STD_LOGIC;
  SIGNAL modulo_sub_30_qelse_and_ssc_1 : STD_LOGIC;
  SIGNAL reg_modulo_sub_30_qr_lpi_3_dfm_1_ftd : STD_LOGIC;
  SIGNAL reg_modulo_sub_30_qr_lpi_3_dfm_1_ftd_1 : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_29_qelse_and_ssc : STD_LOGIC;
  SIGNAL modulo_sub_29_qelse_and_ssc_1 : STD_LOGIC;
  SIGNAL reg_modulo_sub_29_qr_lpi_3_dfm_1_ftd : STD_LOGIC;
  SIGNAL reg_modulo_sub_29_qr_lpi_3_dfm_1_ftd_1 : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_28_qelse_and_ssc : STD_LOGIC;
  SIGNAL modulo_sub_28_qelse_and_ssc_1 : STD_LOGIC;
  SIGNAL reg_modulo_sub_28_qr_lpi_3_dfm_1_ftd : STD_LOGIC;
  SIGNAL reg_modulo_sub_28_qr_lpi_3_dfm_1_ftd_1 : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_27_qelse_and_ssc : STD_LOGIC;
  SIGNAL modulo_sub_27_qelse_and_ssc_1 : STD_LOGIC;
  SIGNAL reg_modulo_sub_27_qr_lpi_3_dfm_1_ftd : STD_LOGIC;
  SIGNAL reg_modulo_sub_27_qr_lpi_3_dfm_1_ftd_1 : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_26_qelse_and_ssc : STD_LOGIC;
  SIGNAL modulo_sub_26_qelse_and_ssc_1 : STD_LOGIC;
  SIGNAL reg_modulo_sub_26_qr_lpi_3_dfm_1_ftd : STD_LOGIC;
  SIGNAL reg_modulo_sub_26_qr_lpi_3_dfm_1_ftd_1 : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_25_qelse_and_ssc : STD_LOGIC;
  SIGNAL modulo_sub_25_qelse_and_ssc_1 : STD_LOGIC;
  SIGNAL reg_modulo_sub_25_qr_lpi_3_dfm_1_ftd : STD_LOGIC;
  SIGNAL reg_modulo_sub_25_qr_lpi_3_dfm_1_ftd_1 : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_24_qelse_and_ssc : STD_LOGIC;
  SIGNAL modulo_sub_24_qelse_and_ssc_1 : STD_LOGIC;
  SIGNAL reg_modulo_sub_24_qr_lpi_3_dfm_1_ftd : STD_LOGIC;
  SIGNAL reg_modulo_sub_24_qr_lpi_3_dfm_1_ftd_1 : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_23_qelse_and_ssc : STD_LOGIC;
  SIGNAL modulo_sub_23_qelse_and_ssc_1 : STD_LOGIC;
  SIGNAL reg_modulo_sub_23_qr_lpi_3_dfm_1_ftd : STD_LOGIC;
  SIGNAL reg_modulo_sub_23_qr_lpi_3_dfm_1_ftd_1 : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_22_qelse_and_ssc : STD_LOGIC;
  SIGNAL modulo_sub_22_qelse_and_ssc_1 : STD_LOGIC;
  SIGNAL reg_modulo_sub_22_qr_lpi_3_dfm_1_ftd : STD_LOGIC;
  SIGNAL reg_modulo_sub_22_qr_lpi_3_dfm_1_ftd_1 : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_21_qelse_and_ssc : STD_LOGIC;
  SIGNAL modulo_sub_21_qelse_and_ssc_1 : STD_LOGIC;
  SIGNAL reg_modulo_sub_21_qr_lpi_3_dfm_1_ftd : STD_LOGIC;
  SIGNAL reg_modulo_sub_21_qr_lpi_3_dfm_1_ftd_1 : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_20_qelse_and_ssc : STD_LOGIC;
  SIGNAL modulo_sub_20_qelse_and_ssc_1 : STD_LOGIC;
  SIGNAL reg_modulo_sub_20_qr_lpi_3_dfm_1_ftd : STD_LOGIC;
  SIGNAL reg_modulo_sub_20_qr_lpi_3_dfm_1_ftd_1 : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_19_qelse_and_ssc : STD_LOGIC;
  SIGNAL modulo_sub_19_qelse_and_ssc_1 : STD_LOGIC;
  SIGNAL reg_modulo_sub_19_qr_lpi_3_dfm_1_ftd : STD_LOGIC;
  SIGNAL reg_modulo_sub_19_qr_lpi_3_dfm_1_ftd_1 : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_18_qelse_and_ssc : STD_LOGIC;
  SIGNAL modulo_sub_18_qelse_and_ssc_1 : STD_LOGIC;
  SIGNAL reg_modulo_sub_18_qr_lpi_3_dfm_1_ftd : STD_LOGIC;
  SIGNAL reg_modulo_sub_18_qr_lpi_3_dfm_1_ftd_1 : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_17_qelse_and_ssc : STD_LOGIC;
  SIGNAL modulo_sub_17_qelse_and_ssc_1 : STD_LOGIC;
  SIGNAL reg_modulo_sub_17_qr_lpi_3_dfm_1_ftd : STD_LOGIC;
  SIGNAL reg_modulo_sub_17_qr_lpi_3_dfm_1_ftd_1 : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_16_qelse_and_ssc : STD_LOGIC;
  SIGNAL modulo_sub_16_qelse_and_ssc_1 : STD_LOGIC;
  SIGNAL reg_modulo_sub_16_qr_lpi_3_dfm_1_ftd : STD_LOGIC;
  SIGNAL reg_modulo_sub_16_qr_lpi_3_dfm_1_ftd_1 : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_add_1_qelse_or_m1c : STD_LOGIC;
  SIGNAL reg_mult_15_res_lpi_3_dfm_1_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_mult_14_res_lpi_3_dfm_1_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_mult_13_res_lpi_3_dfm_1_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_mult_12_res_lpi_3_dfm_1_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_mult_11_res_lpi_3_dfm_1_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_mult_10_res_lpi_3_dfm_1_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_mult_9_res_lpi_3_dfm_1_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_mult_8_res_lpi_3_dfm_1_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_mult_7_res_lpi_3_dfm_1_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_mult_6_res_lpi_3_dfm_1_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_mult_5_res_lpi_3_dfm_1_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_mult_4_res_lpi_3_dfm_1_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_mult_3_res_lpi_3_dfm_1_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_mult_2_res_lpi_3_dfm_1_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_mult_1_res_lpi_3_dfm_1_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_mult_res_lpi_3_dfm_1_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_mult_32_res_lpi_3_dfm_1_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_mult_33_res_lpi_3_dfm_1_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_mult_34_res_lpi_3_dfm_1_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_mult_35_res_lpi_3_dfm_1_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_mult_36_res_lpi_3_dfm_1_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_mult_37_res_lpi_3_dfm_1_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_mult_38_res_lpi_3_dfm_1_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_mult_39_res_lpi_3_dfm_1_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_mult_40_res_lpi_3_dfm_1_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_mult_41_res_lpi_3_dfm_1_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_mult_42_res_lpi_3_dfm_1_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_mult_43_res_lpi_3_dfm_1_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_mult_44_res_lpi_3_dfm_1_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_mult_45_res_lpi_3_dfm_1_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_mult_46_res_lpi_3_dfm_1_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_mult_47_res_lpi_3_dfm_1_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_INNER_LOOP1_r_and_cse : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_INNER_LOOP1_r_and_3_cse : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_INNER_LOOP1_r_and_5_cse : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL butterFly1_15_f1_mux_cse : STD_LOGIC;
  SIGNAL butterFly1_15_f1_mux_1_cse : STD_LOGIC;
  SIGNAL butterFly1_15_f1_mux_2_cse : STD_LOGIC;
  SIGNAL butterFly1_15_f1_mux_3_cse : STD_LOGIC;
  SIGNAL butterFly1_15_f1_mux_4_cse : STD_LOGIC;
  SIGNAL butterFly1_15_f1_mux_5_cse : STD_LOGIC;
  SIGNAL butterFly1_15_f1_mux_6_cse : STD_LOGIC;
  SIGNAL butterFly1_15_f1_mux_7_cse : STD_LOGIC;
  SIGNAL butterFly1_31_f1_mux_cse : STD_LOGIC;
  SIGNAL butterFly1_31_f1_mux_1_cse : STD_LOGIC;
  SIGNAL butterFly1_31_f1_mux_2_cse : STD_LOGIC;
  SIGNAL butterFly1_31_f1_mux_3_cse : STD_LOGIC;
  SIGNAL butterFly1_31_f1_mux_4_cse : STD_LOGIC;
  SIGNAL butterFly1_31_f1_mux_5_cse : STD_LOGIC;
  SIGNAL butterFly1_31_f1_mux_6_cse : STD_LOGIC;
  SIGNAL butterFly1_31_f1_mux_7_cse : STD_LOGIC;
  SIGNAL butterFly2_f1_mux_cse : STD_LOGIC;
  SIGNAL butterFly2_f1_mux_1_cse : STD_LOGIC;
  SIGNAL butterFly2_f1_mux_2_cse : STD_LOGIC;
  SIGNAL butterFly2_f1_mux_3_cse : STD_LOGIC;
  SIGNAL butterFly2_f1_mux_4_cse : STD_LOGIC;
  SIGNAL butterFly2_f1_mux_5_cse : STD_LOGIC;
  SIGNAL butterFly2_f1_mux_6_cse : STD_LOGIC;
  SIGNAL butterFly2_f1_mux_7_cse : STD_LOGIC;
  SIGNAL butterFly2_21_f1_mux_cse : STD_LOGIC;
  SIGNAL butterFly2_21_f1_mux_1_cse : STD_LOGIC;
  SIGNAL butterFly2_21_f1_mux_2_cse : STD_LOGIC;
  SIGNAL butterFly2_21_f1_mux_3_cse : STD_LOGIC;
  SIGNAL butterFly2_21_f1_mux_4_cse : STD_LOGIC;
  SIGNAL butterFly2_21_f1_mux_5_cse : STD_LOGIC;
  SIGNAL butterFly2_21_f1_mux_6_cse : STD_LOGIC;
  SIGNAL butterFly2_21_f1_mux_7_cse : STD_LOGIC;
  SIGNAL or_4976_cse : STD_LOGIC;
  SIGNAL z_out_143_32 : STD_LOGIC;
  SIGNAL z_out_144_32 : STD_LOGIC;
  SIGNAL z_out_145_32 : STD_LOGIC;
  SIGNAL z_out_146_32 : STD_LOGIC;
  SIGNAL z_out_147_32 : STD_LOGIC;
  SIGNAL z_out_148_32 : STD_LOGIC;
  SIGNAL z_out_149_32 : STD_LOGIC;
  SIGNAL z_out_150_32 : STD_LOGIC;
  SIGNAL z_out_151_32 : STD_LOGIC;
  SIGNAL z_out_152_32 : STD_LOGIC;
  SIGNAL z_out_153_32 : STD_LOGIC;
  SIGNAL z_out_154_32 : STD_LOGIC;
  SIGNAL z_out_155_32 : STD_LOGIC;
  SIGNAL z_out_156_32 : STD_LOGIC;
  SIGNAL z_out_157_32 : STD_LOGIC;
  SIGNAL z_out_158_32 : STD_LOGIC;

  SIGNAL c_mux_nl : STD_LOGIC;
  SIGNAL butterFly2_21_tw_butterFly2_21_tw_or_nl : STD_LOGIC;
  SIGNAL mux_2_nl : STD_LOGIC;
  SIGNAL mux_1_nl : STD_LOGIC;
  SIGNAL or_322_nl : STD_LOGIC;
  SIGNAL mux_6_nl : STD_LOGIC;
  SIGNAL mux_5_nl : STD_LOGIC;
  SIGNAL or_337_nl : STD_LOGIC;
  SIGNAL mux_9_nl : STD_LOGIC;
  SIGNAL mux_8_nl : STD_LOGIC;
  SIGNAL or_344_nl : STD_LOGIC;
  SIGNAL mux_11_nl : STD_LOGIC;
  SIGNAL mux_10_nl : STD_LOGIC;
  SIGNAL or_352_nl : STD_LOGIC;
  SIGNAL mux_13_nl : STD_LOGIC;
  SIGNAL or_356_nl : STD_LOGIC;
  SIGNAL mux_12_nl : STD_LOGIC;
  SIGNAL mux_17_nl : STD_LOGIC;
  SIGNAL mux_16_nl : STD_LOGIC;
  SIGNAL or_360_nl : STD_LOGIC;
  SIGNAL mux_19_nl : STD_LOGIC;
  SIGNAL or_367_nl : STD_LOGIC;
  SIGNAL mux_18_nl : STD_LOGIC;
  SIGNAL mux_21_nl : STD_LOGIC;
  SIGNAL mux_20_nl : STD_LOGIC;
  SIGNAL or_368_nl : STD_LOGIC;
  SIGNAL mux_24_nl : STD_LOGIC;
  SIGNAL mux_23_nl : STD_LOGIC;
  SIGNAL or_372_nl : STD_LOGIC;
  SIGNAL mux_28_nl : STD_LOGIC;
  SIGNAL mux_27_nl : STD_LOGIC;
  SIGNAL mux_31_nl : STD_LOGIC;
  SIGNAL mux_30_nl : STD_LOGIC;
  SIGNAL nor_49_nl : STD_LOGIC;
  SIGNAL mux_32_nl : STD_LOGIC;
  SIGNAL nor_50_nl : STD_LOGIC;
  SIGNAL mux_34_nl : STD_LOGIC;
  SIGNAL nand_1_nl : STD_LOGIC;
  SIGNAL mux_33_nl : STD_LOGIC;
  SIGNAL mux_39_nl : STD_LOGIC;
  SIGNAL mux_38_nl : STD_LOGIC;
  SIGNAL mux_42_nl : STD_LOGIC;
  SIGNAL mux_41_nl : STD_LOGIC;
  SIGNAL mux_43_nl : STD_LOGIC;
  SIGNAL or_404_nl : STD_LOGIC;
  SIGNAL mux_47_nl : STD_LOGIC;
  SIGNAL mux_46_nl : STD_LOGIC;
  SIGNAL or_406_nl : STD_LOGIC;
  SIGNAL mux_52_nl : STD_LOGIC;
  SIGNAL mux_51_nl : STD_LOGIC;
  SIGNAL mux_55_nl : STD_LOGIC;
  SIGNAL mux_54_nl : STD_LOGIC;
  SIGNAL or_426_nl : STD_LOGIC;
  SIGNAL mux_58_nl : STD_LOGIC;
  SIGNAL mux_57_nl : STD_LOGIC;
  SIGNAL mux_60_nl : STD_LOGIC;
  SIGNAL or_433_nl : STD_LOGIC;
  SIGNAL mux_59_nl : STD_LOGIC;
  SIGNAL mux_64_nl : STD_LOGIC;
  SIGNAL mux_63_nl : STD_LOGIC;
  SIGNAL mux_66_nl : STD_LOGIC;
  SIGNAL or_442_nl : STD_LOGIC;
  SIGNAL mux_65_nl : STD_LOGIC;
  SIGNAL mux_68_nl : STD_LOGIC;
  SIGNAL mux_67_nl : STD_LOGIC;
  SIGNAL mux_72_nl : STD_LOGIC;
  SIGNAL mux_71_nl : STD_LOGIC;
  SIGNAL or_444_nl : STD_LOGIC;
  SIGNAL mux_76_nl : STD_LOGIC;
  SIGNAL mux_75_nl : STD_LOGIC;
  SIGNAL mux_80_nl : STD_LOGIC;
  SIGNAL mux_79_nl : STD_LOGIC;
  SIGNAL nor_48_nl : STD_LOGIC;
  SIGNAL mux_82_nl : STD_LOGIC;
  SIGNAL mux_81_nl : STD_LOGIC;
  SIGNAL mux_84_nl : STD_LOGIC;
  SIGNAL nand_nl : STD_LOGIC;
  SIGNAL mux_83_nl : STD_LOGIC;
  SIGNAL mux_88_nl : STD_LOGIC;
  SIGNAL mux_87_nl : STD_LOGIC;
  SIGNAL mux_90_nl : STD_LOGIC;
  SIGNAL mux_89_nl : STD_LOGIC;
  SIGNAL mux_92_nl : STD_LOGIC;
  SIGNAL mux_91_nl : STD_LOGIC;
  SIGNAL mult_4_t_and_nl : STD_LOGIC;
  SIGNAL mult_4_t_and_1_nl : STD_LOGIC;
  SIGNAL mult_4_t_and_2_nl : STD_LOGIC;
  SIGNAL mult_4_t_and_3_nl : STD_LOGIC;
  SIGNAL mult_4_t_and_4_nl : STD_LOGIC;
  SIGNAL mult_4_t_and_5_nl : STD_LOGIC;
  SIGNAL mult_4_t_and_6_nl : STD_LOGIC;
  SIGNAL mult_4_t_and_7_nl : STD_LOGIC;
  SIGNAL mult_4_t_and_8_nl : STD_LOGIC;
  SIGNAL mult_4_t_and_9_nl : STD_LOGIC;
  SIGNAL mult_4_t_and_10_nl : STD_LOGIC;
  SIGNAL mult_4_t_and_11_nl : STD_LOGIC;
  SIGNAL mult_4_t_and_12_nl : STD_LOGIC;
  SIGNAL mult_4_t_and_13_nl : STD_LOGIC;
  SIGNAL mult_4_t_and_14_nl : STD_LOGIC;
  SIGNAL mult_4_t_and_15_nl : STD_LOGIC;
  SIGNAL mult_4_t_and_16_nl : STD_LOGIC;
  SIGNAL mult_4_t_and_17_nl : STD_LOGIC;
  SIGNAL mult_4_t_and_18_nl : STD_LOGIC;
  SIGNAL mult_4_t_and_19_nl : STD_LOGIC;
  SIGNAL mult_4_t_and_20_nl : STD_LOGIC;
  SIGNAL mult_4_t_and_21_nl : STD_LOGIC;
  SIGNAL mult_4_t_and_22_nl : STD_LOGIC;
  SIGNAL mult_4_t_and_23_nl : STD_LOGIC;
  SIGNAL mult_4_t_and_24_nl : STD_LOGIC;
  SIGNAL mult_4_t_and_25_nl : STD_LOGIC;
  SIGNAL mult_4_t_and_26_nl : STD_LOGIC;
  SIGNAL mult_4_t_and_27_nl : STD_LOGIC;
  SIGNAL mult_4_t_and_28_nl : STD_LOGIC;
  SIGNAL mult_4_t_and_29_nl : STD_LOGIC;
  SIGNAL mult_4_t_and_30_nl : STD_LOGIC;
  SIGNAL mult_4_t_and_31_nl : STD_LOGIC;
  SIGNAL STAGE_LOOP_mux1h_nl : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL acc_2_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_1_qif_mux1h_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_1_qelse_and_nl : STD_LOGIC;
  SIGNAL modulo_add_1_qelse_or_1_nl : STD_LOGIC;
  SIGNAL modulo_add_1_qelse_and_4_nl : STD_LOGIC;
  SIGNAL modulo_add_1_qelse_and_5_nl : STD_LOGIC;
  SIGNAL acc_3_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_10_qif_mux1h_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_10_qelse_and_nl : STD_LOGIC;
  SIGNAL modulo_add_10_qelse_or_nl : STD_LOGIC;
  SIGNAL modulo_add_10_qelse_and_5_nl : STD_LOGIC;
  SIGNAL modulo_add_10_qelse_and_6_nl : STD_LOGIC;
  SIGNAL modulo_add_10_qelse_and_7_nl : STD_LOGIC;
  SIGNAL acc_4_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_11_qif_mux1h_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_11_qelse_and_nl : STD_LOGIC;
  SIGNAL modulo_add_11_qelse_or_nl : STD_LOGIC;
  SIGNAL modulo_add_11_qelse_and_5_nl : STD_LOGIC;
  SIGNAL modulo_add_11_qelse_and_6_nl : STD_LOGIC;
  SIGNAL modulo_add_11_qelse_and_7_nl : STD_LOGIC;
  SIGNAL acc_5_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_12_qif_mux1h_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_12_qelse_and_nl : STD_LOGIC;
  SIGNAL modulo_add_12_qelse_or_1_nl : STD_LOGIC;
  SIGNAL modulo_add_12_qelse_and_4_nl : STD_LOGIC;
  SIGNAL modulo_add_12_qelse_and_5_nl : STD_LOGIC;
  SIGNAL acc_6_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_13_qif_mux1h_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_13_qelse_and_nl : STD_LOGIC;
  SIGNAL modulo_add_13_qelse_or_1_nl : STD_LOGIC;
  SIGNAL modulo_add_13_qelse_and_4_nl : STD_LOGIC;
  SIGNAL modulo_add_13_qelse_and_5_nl : STD_LOGIC;
  SIGNAL acc_10_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_14_qif_mux1h_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_14_qelse_and_nl : STD_LOGIC;
  SIGNAL modulo_add_14_qelse_or_1_nl : STD_LOGIC;
  SIGNAL modulo_add_14_qelse_and_4_nl : STD_LOGIC;
  SIGNAL modulo_add_14_qelse_and_5_nl : STD_LOGIC;
  SIGNAL acc_14_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_15_qif_mux1h_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_15_qelse_and_nl : STD_LOGIC;
  SIGNAL modulo_add_15_qelse_or_nl : STD_LOGIC;
  SIGNAL modulo_add_15_qelse_and_5_nl : STD_LOGIC;
  SIGNAL modulo_add_15_qelse_and_6_nl : STD_LOGIC;
  SIGNAL modulo_add_15_qelse_and_7_nl : STD_LOGIC;
  SIGNAL butterFly1_f1_butterFly1_f1_nor_nl : STD_LOGIC;
  SIGNAL butterFly1_16_f1_butterFly1_16_f1_nor_nl : STD_LOGIC;
  SIGNAL butterFly2_f1_butterFly2_f1_and_5_nl : STD_LOGIC;
  SIGNAL butterFly2_16_f1_butterFly2_16_f1_and_5_nl : STD_LOGIC;
  SIGNAL butterFly1_f1_butterFly1_f1_and_nl : STD_LOGIC;
  SIGNAL butterFly1_16_f1_butterFly1_16_f1_and_nl : STD_LOGIC;
  SIGNAL butterFly1_f1_butterFly1_f1_and_1_nl : STD_LOGIC;
  SIGNAL butterFly1_16_f1_butterFly1_16_f1_and_1_nl : STD_LOGIC;
  SIGNAL butterFly1_f1_butterFly1_f1_and_2_nl : STD_LOGIC;
  SIGNAL butterFly1_16_f1_butterFly1_16_f1_and_2_nl : STD_LOGIC;
  SIGNAL butterFly2_f1_butterFly2_f1_and_nl : STD_LOGIC;
  SIGNAL butterFly2_16_f1_butterFly2_16_f1_and_nl : STD_LOGIC;
  SIGNAL butterFly1_f1_butterFly1_f1_and_3_nl : STD_LOGIC;
  SIGNAL butterFly1_16_f1_butterFly1_16_f1_and_3_nl : STD_LOGIC;
  SIGNAL butterFly2_f1_butterFly2_f1_and_1_nl : STD_LOGIC;
  SIGNAL butterFly2_16_f1_butterFly2_16_f1_and_1_nl : STD_LOGIC;
  SIGNAL butterFly1_f1_butterFly1_f1_and_4_nl : STD_LOGIC;
  SIGNAL butterFly1_16_f1_butterFly1_16_f1_and_4_nl : STD_LOGIC;
  SIGNAL butterFly2_f1_butterFly2_f1_and_2_nl : STD_LOGIC;
  SIGNAL butterFly2_16_f1_butterFly2_16_f1_and_2_nl : STD_LOGIC;
  SIGNAL butterFly1_f1_butterFly1_f1_and_5_nl : STD_LOGIC;
  SIGNAL butterFly1_16_f1_butterFly1_16_f1_and_5_nl : STD_LOGIC;
  SIGNAL butterFly2_f1_butterFly2_f1_and_3_nl : STD_LOGIC;
  SIGNAL butterFly2_16_f1_butterFly2_16_f1_and_3_nl : STD_LOGIC;
  SIGNAL butterFly1_f1_butterFly1_f1_and_6_nl : STD_LOGIC;
  SIGNAL butterFly1_16_f1_butterFly1_16_f1_and_6_nl : STD_LOGIC;
  SIGNAL butterFly2_f1_butterFly2_f1_and_4_nl : STD_LOGIC;
  SIGNAL butterFly2_16_f1_butterFly2_16_f1_and_4_nl : STD_LOGIC;
  SIGNAL INNER_LOOP1_mux_nl : STD_LOGIC;
  SIGNAL INNER_LOOP1_mux_4_nl : STD_LOGIC;
  SIGNAL INNER_LOOP1_mux_5_nl : STD_LOGIC;
  SIGNAL INNER_LOOP1_mux_6_nl : STD_LOGIC;
  SIGNAL butterFly1_15_mux_9_nl : STD_LOGIC;
  SIGNAL butterFly1_15_mux1h_47_nl : STD_LOGIC;
  SIGNAL butterFly2_15_mux1h_3_nl : STD_LOGIC;
  SIGNAL butterFly1_15_mux_10_nl : STD_LOGIC;
  SIGNAL STAGE_LOOP_base_STAGE_LOOP_base_mux_nl : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL INNER_LOOP2_r_or_nl : STD_LOGIC;
  SIGNAL acc_18_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_2_qif_mux1h_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_23_qelse_and_nl : STD_LOGIC;
  SIGNAL modulo_add_23_qelse_or_1_nl : STD_LOGIC;
  SIGNAL modulo_add_23_qelse_and_4_nl : STD_LOGIC;
  SIGNAL modulo_add_23_qelse_and_5_nl : STD_LOGIC;
  SIGNAL acc_22_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_3_qif_mux1h_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_24_qelse_and_nl : STD_LOGIC;
  SIGNAL modulo_add_24_qelse_or_1_nl : STD_LOGIC;
  SIGNAL modulo_add_24_qelse_and_4_nl : STD_LOGIC;
  SIGNAL modulo_add_24_qelse_and_5_nl : STD_LOGIC;
  SIGNAL acc_26_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_4_qif_mux1h_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_25_qelse_and_nl : STD_LOGIC;
  SIGNAL modulo_add_25_qelse_or_1_nl : STD_LOGIC;
  SIGNAL modulo_add_25_qelse_and_4_nl : STD_LOGIC;
  SIGNAL modulo_add_25_qelse_and_5_nl : STD_LOGIC;
  SIGNAL acc_30_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_5_qif_mux1h_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_26_qelse_and_nl : STD_LOGIC;
  SIGNAL modulo_add_26_qelse_or_nl : STD_LOGIC;
  SIGNAL modulo_add_26_qelse_and_5_nl : STD_LOGIC;
  SIGNAL modulo_add_26_qelse_and_6_nl : STD_LOGIC;
  SIGNAL modulo_add_26_qelse_and_7_nl : STD_LOGIC;
  SIGNAL acc_34_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_6_qif_mux1h_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_27_qelse_and_nl : STD_LOGIC;
  SIGNAL modulo_add_27_qelse_or_nl : STD_LOGIC;
  SIGNAL modulo_add_27_qelse_and_5_nl : STD_LOGIC;
  SIGNAL modulo_add_27_qelse_and_6_nl : STD_LOGIC;
  SIGNAL modulo_add_27_qelse_and_7_nl : STD_LOGIC;
  SIGNAL acc_38_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_7_qif_mux1h_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_28_qelse_and_nl : STD_LOGIC;
  SIGNAL modulo_add_28_qelse_or_nl : STD_LOGIC;
  SIGNAL modulo_add_28_qelse_and_5_nl : STD_LOGIC;
  SIGNAL modulo_add_28_qelse_and_6_nl : STD_LOGIC;
  SIGNAL modulo_add_28_qelse_and_7_nl : STD_LOGIC;
  SIGNAL acc_42_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_8_qif_mux1h_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_29_qelse_and_nl : STD_LOGIC;
  SIGNAL modulo_add_29_qelse_or_nl : STD_LOGIC;
  SIGNAL modulo_add_29_qelse_and_5_nl : STD_LOGIC;
  SIGNAL modulo_add_29_qelse_and_6_nl : STD_LOGIC;
  SIGNAL modulo_add_29_qelse_and_7_nl : STD_LOGIC;
  SIGNAL acc_46_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_9_qif_mux1h_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_30_qelse_and_nl : STD_LOGIC;
  SIGNAL modulo_add_30_qelse_or_nl : STD_LOGIC;
  SIGNAL modulo_add_30_qelse_and_5_nl : STD_LOGIC;
  SIGNAL modulo_add_30_qelse_and_6_nl : STD_LOGIC;
  SIGNAL modulo_add_30_qelse_and_7_nl : STD_LOGIC;
  SIGNAL acc_49_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_qif_mux1h_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_31_qelse_and_nl : STD_LOGIC;
  SIGNAL modulo_add_31_qelse_or_nl : STD_LOGIC;
  SIGNAL modulo_add_31_qelse_and_5_nl : STD_LOGIC;
  SIGNAL modulo_add_31_qelse_and_6_nl : STD_LOGIC;
  SIGNAL modulo_add_31_qelse_and_7_nl : STD_LOGIC;
  SIGNAL modulo_sub_16_qelse_or_nl : STD_LOGIC;
  SIGNAL modulo_sub_17_qelse_or_nl : STD_LOGIC;
  SIGNAL modulo_sub_18_qelse_or_nl : STD_LOGIC;
  SIGNAL modulo_sub_19_qelse_or_nl : STD_LOGIC;
  SIGNAL modulo_sub_20_qelse_or_nl : STD_LOGIC;
  SIGNAL modulo_sub_21_qelse_or_nl : STD_LOGIC;
  SIGNAL modulo_sub_22_qelse_or_nl : STD_LOGIC;
  SIGNAL modulo_sub_23_qelse_or_nl : STD_LOGIC;
  SIGNAL modulo_sub_24_qelse_or_nl : STD_LOGIC;
  SIGNAL modulo_sub_25_qelse_or_nl : STD_LOGIC;
  SIGNAL modulo_sub_26_qelse_or_nl : STD_LOGIC;
  SIGNAL modulo_sub_27_qelse_or_nl : STD_LOGIC;
  SIGNAL modulo_sub_28_qelse_or_nl : STD_LOGIC;
  SIGNAL modulo_sub_29_qelse_or_nl : STD_LOGIC;
  SIGNAL modulo_sub_30_qelse_or_nl : STD_LOGIC;
  SIGNAL modulo_sub_31_qelse_or_nl : STD_LOGIC;
  SIGNAL INNER_LOOP1_mux_7_nl : STD_LOGIC;
  SIGNAL butterFly2_f1_butterFly2_f1_nor_nl : STD_LOGIC;
  SIGNAL butterFly2_16_f1_butterFly2_16_f1_nor_nl : STD_LOGIC;
  SIGNAL butterFly2_f1_butterFly2_f1_and_6_nl : STD_LOGIC;
  SIGNAL mult_15_if_acc_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_31_acc_1_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL mult_14_if_acc_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_30_acc_1_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL mult_13_if_acc_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_29_acc_1_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL mult_12_if_acc_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_28_acc_1_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL mult_11_if_acc_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_27_acc_1_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL mult_10_if_acc_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_26_acc_1_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL mult_9_if_acc_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_25_acc_1_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL mult_8_if_acc_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_24_acc_1_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL mult_7_if_acc_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_23_acc_1_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL mult_6_if_acc_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_22_acc_1_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL mult_5_if_acc_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_21_acc_1_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL mult_4_if_acc_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_20_acc_1_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL mult_3_if_acc_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_19_acc_1_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL mult_2_if_acc_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_18_acc_1_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL mult_1_if_acc_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_17_acc_1_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL mult_if_acc_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_16_acc_1_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL nor_62_nl : STD_LOGIC;
  SIGNAL or_325_nl : STD_LOGIC;
  SIGNAL nor_56_nl : STD_LOGIC;
  SIGNAL or_347_nl : STD_LOGIC;
  SIGNAL and_8934_nl : STD_LOGIC;
  SIGNAL mux_44_nl : STD_LOGIC;
  SIGNAL or_409_nl : STD_LOGIC;
  SIGNAL or_408_nl : STD_LOGIC;
  SIGNAL or_419_nl : STD_LOGIC;
  SIGNAL nor_52_nl : STD_LOGIC;
  SIGNAL or_427_nl : STD_LOGIC;
  SIGNAL or_429_nl : STD_LOGIC;
  SIGNAL or_447_nl : STD_LOGIC;
  SIGNAL mux_69_nl : STD_LOGIC;
  SIGNAL or_445_nl : STD_LOGIC;
  SIGNAL or_457_nl : STD_LOGIC;
  SIGNAL mux_4_nl : STD_LOGIC;
  SIGNAL mux_3_nl : STD_LOGIC;
  SIGNAL or_332_nl : STD_LOGIC;
  SIGNAL or_331_nl : STD_LOGIC;
  SIGNAL mux_15_nl : STD_LOGIC;
  SIGNAL or_359_nl : STD_LOGIC;
  SIGNAL mux_14_nl : STD_LOGIC;
  SIGNAL or_357_nl : STD_LOGIC;
  SIGNAL nor_3_nl : STD_LOGIC;
  SIGNAL mux_26_nl : STD_LOGIC;
  SIGNAL mux_25_nl : STD_LOGIC;
  SIGNAL nor_7_nl : STD_LOGIC;
  SIGNAL nor_64_nl : STD_LOGIC;
  SIGNAL mux_29_nl : STD_LOGIC;
  SIGNAL and_8944_nl : STD_LOGIC;
  SIGNAL mux_37_nl : STD_LOGIC;
  SIGNAL mux_36_nl : STD_LOGIC;
  SIGNAL mux_35_nl : STD_LOGIC;
  SIGNAL nor_20_nl : STD_LOGIC;
  SIGNAL mux_40_nl : STD_LOGIC;
  SIGNAL and_8943_nl : STD_LOGIC;
  SIGNAL mux_49_nl : STD_LOGIC;
  SIGNAL mux_48_nl : STD_LOGIC;
  SIGNAL or_415_nl : STD_LOGIC;
  SIGNAL or_414_nl : STD_LOGIC;
  SIGNAL mux_62_nl : STD_LOGIC;
  SIGNAL nand_17_nl : STD_LOGIC;
  SIGNAL mux_61_nl : STD_LOGIC;
  SIGNAL or_434_nl : STD_LOGIC;
  SIGNAL mux_74_nl : STD_LOGIC;
  SIGNAL mux_73_nl : STD_LOGIC;
  SIGNAL nor_31_nl : STD_LOGIC;
  SIGNAL nor_63_nl : STD_LOGIC;
  SIGNAL mux_77_nl : STD_LOGIC;
  SIGNAL and_8942_nl : STD_LOGIC;
  SIGNAL mux_86_nl : STD_LOGIC;
  SIGNAL mux_85_nl : STD_LOGIC;
  SIGNAL INNER_LOOP1_tw_and_nl : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL INNER_LOOP2_tw_and_nl : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL butterFly1_and_4_nl : STD_LOGIC;
  SIGNAL butterFly1_mux1h_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL butterFly1_or_nl : STD_LOGIC;
  SIGNAL butterFly1_1_and_4_nl : STD_LOGIC;
  SIGNAL butterFly1_1_mux_nl : STD_LOGIC;
  SIGNAL butterFly1_1_mux1h_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL butterFly1_1_and_1_nl : STD_LOGIC;
  SIGNAL butterFly1_2_and_4_nl : STD_LOGIC;
  SIGNAL butterFly1_2_mux_nl : STD_LOGIC;
  SIGNAL butterFly1_2_mux1h_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL butterFly1_2_and_1_nl : STD_LOGIC;
  SIGNAL butterFly1_3_and_4_nl : STD_LOGIC;
  SIGNAL butterFly1_3_mux_nl : STD_LOGIC;
  SIGNAL butterFly1_3_mux1h_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL butterFly1_3_and_1_nl : STD_LOGIC;
  SIGNAL butterFly1_4_and_4_nl : STD_LOGIC;
  SIGNAL butterFly1_4_mux_nl : STD_LOGIC;
  SIGNAL butterFly1_4_mux1h_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL butterFly1_4_and_1_nl : STD_LOGIC;
  SIGNAL butterFly1_5_and_4_nl : STD_LOGIC;
  SIGNAL butterFly1_5_mux_nl : STD_LOGIC;
  SIGNAL butterFly1_5_mux1h_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL butterFly1_5_and_1_nl : STD_LOGIC;
  SIGNAL butterFly1_6_and_4_nl : STD_LOGIC;
  SIGNAL butterFly1_6_mux_nl : STD_LOGIC;
  SIGNAL butterFly1_6_mux1h_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL butterFly1_6_and_1_nl : STD_LOGIC;
  SIGNAL butterFly1_7_and_4_nl : STD_LOGIC;
  SIGNAL butterFly1_7_mux_nl : STD_LOGIC;
  SIGNAL butterFly1_7_mux1h_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL butterFly1_7_and_1_nl : STD_LOGIC;
  SIGNAL butterFly1_8_and_4_nl : STD_LOGIC;
  SIGNAL butterFly1_8_mux_nl : STD_LOGIC;
  SIGNAL butterFly1_8_mux1h_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL butterFly1_8_and_1_nl : STD_LOGIC;
  SIGNAL butterFly1_9_and_4_nl : STD_LOGIC;
  SIGNAL butterFly1_9_mux_nl : STD_LOGIC;
  SIGNAL butterFly1_9_mux1h_272_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL butterFly1_9_and_1_nl : STD_LOGIC;
  SIGNAL butterFly1_10_and_4_nl : STD_LOGIC;
  SIGNAL butterFly1_10_mux_nl : STD_LOGIC;
  SIGNAL butterFly1_10_mux1h_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL butterFly1_10_and_1_nl : STD_LOGIC;
  SIGNAL butterFly1_11_and_4_nl : STD_LOGIC;
  SIGNAL butterFly1_11_mux_nl : STD_LOGIC;
  SIGNAL butterFly1_11_mux1h_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL butterFly1_11_and_1_nl : STD_LOGIC;
  SIGNAL butterFly1_12_and_4_nl : STD_LOGIC;
  SIGNAL butterFly1_12_mux_nl : STD_LOGIC;
  SIGNAL butterFly1_12_mux1h_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL butterFly1_12_and_1_nl : STD_LOGIC;
  SIGNAL butterFly1_13_and_4_nl : STD_LOGIC;
  SIGNAL butterFly1_13_mux_nl : STD_LOGIC;
  SIGNAL butterFly1_13_mux1h_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL butterFly1_13_and_1_nl : STD_LOGIC;
  SIGNAL butterFly1_14_and_4_nl : STD_LOGIC;
  SIGNAL butterFly1_14_mux_nl : STD_LOGIC;
  SIGNAL butterFly1_14_mux1h_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL butterFly1_14_and_1_nl : STD_LOGIC;
  SIGNAL butterFly1_15_and_5_nl : STD_LOGIC;
  SIGNAL butterFly1_15_mux1h_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL butterFly1_15_or_nl : STD_LOGIC;
  SIGNAL operator_20_false_mux_2_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL operator_20_false_mux1h_2_nl : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL modulo_sub_15_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_31_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_7_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_30_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_39_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_29_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_6_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_28_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_38_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_27_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_5_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_26_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_37_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_25_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_4_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_24_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_36_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_23_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_3_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_22_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_35_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_21_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_2_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_20_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_34_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_19_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_1_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_18_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_33_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_17_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_16_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL acc_50_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL butterFly1_mux1h_18_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_51_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL butterFly1_1_mux1h_18_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_52_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL butterFly1_2_mux1h_18_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_53_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL butterFly1_3_mux1h_18_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_54_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL butterFly1_4_mux1h_18_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_55_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL butterFly1_5_mux1h_18_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_56_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL butterFly1_6_mux1h_18_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_57_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL butterFly1_7_mux1h_18_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_58_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL butterFly1_8_mux1h_18_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_59_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL butterFly1_9_mux1h_274_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_60_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL butterFly1_10_mux1h_18_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_61_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL butterFly1_11_mux1h_18_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_62_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL butterFly1_12_mux1h_18_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_63_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL butterFly1_13_mux1h_18_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_64_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL butterFly1_14_mux1h_18_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_65_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL butterFly1_15_mux1h_79_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_15_mux1h_80_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_14_mux1h_19_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_13_mux1h_19_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_12_mux1h_19_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_11_mux1h_19_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_10_mux1h_19_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_9_mux1h_275_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_8_mux1h_19_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_7_mux1h_19_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_6_mux1h_19_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_5_mux1h_19_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_4_mux1h_19_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_3_mux1h_19_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_2_mux1h_19_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_1_mux1h_19_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_mux1h_19_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_82_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL modulo_add_1_mux1h_3_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_83_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL modulo_add_10_mux1h_3_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_84_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL modulo_add_54_mux1h_3_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_85_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL modulo_add_48_mux1h_3_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_86_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL modulo_add_33_mux1h_3_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_87_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL modulo_add_34_mux1h_3_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_88_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL modulo_add_6_mux1h_3_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_89_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL modulo_add_50_mux1h_3_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_90_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL modulo_add_51_mux1h_3_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_91_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL modulo_add_14_mux1h_3_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_92_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL modulo_add_36_mux1h_3_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_93_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL modulo_add_52_mux1h_3_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_94_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL modulo_add_41_mux1h_3_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_95_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL modulo_add_2_mux1h_3_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_96_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL modulo_add_53_mux1h_3_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_97_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL modulo_add_55_mux1h_3_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL p_rsci_dat : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL p_rsci_idat_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_t_mul_cmp_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_z_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL mult_t_mul_cmp_1_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_1_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_1_z_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL mult_t_mul_cmp_2_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_2_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_2_z_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL mult_t_mul_cmp_3_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_3_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_3_z_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL mult_t_mul_cmp_4_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_4_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_4_z_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL mult_t_mul_cmp_5_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_5_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_5_z_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL mult_t_mul_cmp_6_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_6_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_6_z_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL mult_t_mul_cmp_7_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_7_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_7_z_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL mult_t_mul_cmp_8_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_8_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_8_z_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL mult_t_mul_cmp_9_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_9_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_9_z_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL mult_t_mul_cmp_10_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_10_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_10_z_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL mult_t_mul_cmp_11_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_11_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_11_z_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL mult_t_mul_cmp_12_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_12_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_12_z_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL mult_t_mul_cmp_13_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_13_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_13_z_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL mult_t_mul_cmp_14_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_14_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_14_z_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL mult_t_mul_cmp_15_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_15_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_15_z_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_1_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_1_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_1_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_2_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_2_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_2_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_3_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_3_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_3_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_4_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_4_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_4_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_5_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_5_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_5_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_6_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_6_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_6_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_7_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_7_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_7_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_8_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_8_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_8_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_9_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_9_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_9_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_10_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_10_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_10_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_11_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_11_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_11_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_12_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_12_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_12_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_13_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_13_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_13_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_14_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_14_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_14_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_15_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_15_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_15_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_16_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_16_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_16_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_17_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_17_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_17_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_18_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_18_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_18_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_19_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_19_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_19_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_20_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_20_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_20_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_21_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_21_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_21_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_22_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_22_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_22_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_23_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_23_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_23_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_24_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_24_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_24_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_25_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_25_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_25_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_26_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_26_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_26_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_27_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_27_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_27_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_28_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_28_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_28_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_29_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_29_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_29_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_30_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_30_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_30_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_31_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_31_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_31_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL operator_33_true_3_lshift_rg_a : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL operator_33_true_3_lshift_rg_s : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL operator_33_true_3_lshift_rg_z : STD_LOGIC_VECTOR (1 DOWNTO 0);

  SIGNAL operator_33_true_1_lshift_rg_a : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL operator_33_true_1_lshift_rg_s : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL operator_33_true_1_lshift_rg_z : STD_LOGIC_VECTOR (10 DOWNTO 0);

  COMPONENT peaseNTT_core_wait_dp
    PORT(
      yt_rsc_0_0_cgo_iro : IN STD_LOGIC;
      yt_rsc_0_0_i_clkr_en_d : OUT STD_LOGIC;
      yt_rsc_0_16_cgo_iro : IN STD_LOGIC;
      yt_rsc_0_16_i_clkr_en_d : OUT STD_LOGIC;
      yt_rsc_1_0_cgo_iro : IN STD_LOGIC;
      yt_rsc_1_0_i_clkr_en_d : OUT STD_LOGIC;
      yt_rsc_1_16_cgo_iro : IN STD_LOGIC;
      yt_rsc_1_16_i_clkr_en_d : OUT STD_LOGIC;
      yt_rsc_2_0_cgo_iro : IN STD_LOGIC;
      yt_rsc_2_0_i_clkr_en_d : OUT STD_LOGIC;
      yt_rsc_2_16_cgo_iro : IN STD_LOGIC;
      yt_rsc_2_16_i_clkr_en_d : OUT STD_LOGIC;
      yt_rsc_3_0_cgo_iro : IN STD_LOGIC;
      yt_rsc_3_0_i_clkr_en_d : OUT STD_LOGIC;
      yt_rsc_3_16_cgo_iro : IN STD_LOGIC;
      yt_rsc_3_16_i_clkr_en_d : OUT STD_LOGIC;
      yt_rsc_4_0_cgo_iro : IN STD_LOGIC;
      yt_rsc_4_0_i_clkr_en_d : OUT STD_LOGIC;
      yt_rsc_4_16_cgo_iro : IN STD_LOGIC;
      yt_rsc_4_16_i_clkr_en_d : OUT STD_LOGIC;
      yt_rsc_5_0_cgo_iro : IN STD_LOGIC;
      yt_rsc_5_0_i_clkr_en_d : OUT STD_LOGIC;
      yt_rsc_5_16_cgo_iro : IN STD_LOGIC;
      yt_rsc_5_16_i_clkr_en_d : OUT STD_LOGIC;
      yt_rsc_6_0_cgo_iro : IN STD_LOGIC;
      yt_rsc_6_0_i_clkr_en_d : OUT STD_LOGIC;
      yt_rsc_6_16_cgo_iro : IN STD_LOGIC;
      yt_rsc_6_16_i_clkr_en_d : OUT STD_LOGIC;
      yt_rsc_7_0_cgo_iro : IN STD_LOGIC;
      yt_rsc_7_0_i_clkr_en_d : OUT STD_LOGIC;
      yt_rsc_7_16_cgo_iro : IN STD_LOGIC;
      yt_rsc_7_16_i_clkr_en_d : OUT STD_LOGIC;
      ensig_cgo_iro : IN STD_LOGIC;
      ensig_cgo_iro_17 : IN STD_LOGIC;
      yt_rsc_0_0_cgo : IN STD_LOGIC;
      yt_rsc_0_16_cgo : IN STD_LOGIC;
      yt_rsc_1_0_cgo : IN STD_LOGIC;
      yt_rsc_1_16_cgo : IN STD_LOGIC;
      yt_rsc_2_0_cgo : IN STD_LOGIC;
      yt_rsc_2_16_cgo : IN STD_LOGIC;
      yt_rsc_3_0_cgo : IN STD_LOGIC;
      yt_rsc_3_16_cgo : IN STD_LOGIC;
      yt_rsc_4_0_cgo : IN STD_LOGIC;
      yt_rsc_4_16_cgo : IN STD_LOGIC;
      yt_rsc_5_0_cgo : IN STD_LOGIC;
      yt_rsc_5_16_cgo : IN STD_LOGIC;
      yt_rsc_6_0_cgo : IN STD_LOGIC;
      yt_rsc_6_16_cgo : IN STD_LOGIC;
      yt_rsc_7_0_cgo : IN STD_LOGIC;
      yt_rsc_7_16_cgo : IN STD_LOGIC;
      ensig_cgo : IN STD_LOGIC;
      mult_t_mul_cmp_en : OUT STD_LOGIC;
      ensig_cgo_17 : IN STD_LOGIC;
      mult_z_mul_cmp_1_en : OUT STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_core_fsm
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      fsm_output : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
      INNER_LOOP1_C_0_tr0 : IN STD_LOGIC;
      INNER_LOOP2_C_0_tr0 : IN STD_LOGIC;
      STAGE_LOOP_C_2_tr0 : IN STD_LOGIC;
      INNER_LOOP3_C_0_tr0 : IN STD_LOGIC;
      INNER_LOOP4_C_0_tr0 : IN STD_LOGIC;
      INNER_LOOP4_C_0_tr1 : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_core_fsm_inst_fsm_output : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL peaseNTT_core_core_fsm_inst_INNER_LOOP1_C_0_tr0 : STD_LOGIC;
  SIGNAL peaseNTT_core_core_fsm_inst_INNER_LOOP2_C_0_tr0 : STD_LOGIC;
  SIGNAL peaseNTT_core_core_fsm_inst_STAGE_LOOP_C_2_tr0 : STD_LOGIC;
  SIGNAL peaseNTT_core_core_fsm_inst_INNER_LOOP4_C_0_tr1 : STD_LOGIC;

  FUNCTION CONV_SL_1_1(input_val:BOOLEAN)
  RETURN STD_LOGIC IS
  BEGIN
    IF input_val THEN RETURN '1';ELSE RETURN '0';END IF;
  END;

  FUNCTION MUX1HOT_s_1_3_2(input_2 : STD_LOGIC;
  input_1 : STD_LOGIC;
  input_0 : STD_LOGIC;
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;
    VARIABLE tmp : STD_LOGIC;

    BEGIN
      tmp := sel(0);
      result := input_0 and tmp;
      tmp := sel(1);
      result := result or ( input_1 and tmp);
      tmp := sel(2);
      result := result or ( input_2 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_s_1_4_2(input_3 : STD_LOGIC;
  input_2 : STD_LOGIC;
  input_1 : STD_LOGIC;
  input_0 : STD_LOGIC;
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;
    VARIABLE tmp : STD_LOGIC;

    BEGIN
      tmp := sel(0);
      result := input_0 and tmp;
      tmp := sel(1);
      result := result or ( input_1 and tmp);
      tmp := sel(2);
      result := result or ( input_2 and tmp);
      tmp := sel(3);
      result := result or ( input_3 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_2_3_2(input_2 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(1 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(1 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_2_4_2(input_3 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(1 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(1 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_2_6_2(input_5 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(5 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(1 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(1 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_31_3_2(input_2 : STD_LOGIC_VECTOR(30 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(30 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(30 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(30 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(30 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_31_4_2(input_3 : STD_LOGIC_VECTOR(30 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(30 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(30 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(30 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(30 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(30 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_32_12_2(input_11 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_10 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(11 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
      tmp := (OTHERS=>sel( 9));
      result := result or ( input_9 and tmp);
      tmp := (OTHERS=>sel( 10));
      result := result or ( input_10 and tmp);
      tmp := (OTHERS=>sel( 11));
      result := result or ( input_11 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_32_32_2(input_31 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_30 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_29 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_28 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_27 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_26 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_25 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_24 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_23 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_22 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_21 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_20 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_19 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_18 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_17 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_16 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_15 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_14 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_13 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_12 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_11 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_10 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(31 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
      tmp := (OTHERS=>sel( 9));
      result := result or ( input_9 and tmp);
      tmp := (OTHERS=>sel( 10));
      result := result or ( input_10 and tmp);
      tmp := (OTHERS=>sel( 11));
      result := result or ( input_11 and tmp);
      tmp := (OTHERS=>sel( 12));
      result := result or ( input_12 and tmp);
      tmp := (OTHERS=>sel( 13));
      result := result or ( input_13 and tmp);
      tmp := (OTHERS=>sel( 14));
      result := result or ( input_14 and tmp);
      tmp := (OTHERS=>sel( 15));
      result := result or ( input_15 and tmp);
      tmp := (OTHERS=>sel( 16));
      result := result or ( input_16 and tmp);
      tmp := (OTHERS=>sel( 17));
      result := result or ( input_17 and tmp);
      tmp := (OTHERS=>sel( 18));
      result := result or ( input_18 and tmp);
      tmp := (OTHERS=>sel( 19));
      result := result or ( input_19 and tmp);
      tmp := (OTHERS=>sel( 20));
      result := result or ( input_20 and tmp);
      tmp := (OTHERS=>sel( 21));
      result := result or ( input_21 and tmp);
      tmp := (OTHERS=>sel( 22));
      result := result or ( input_22 and tmp);
      tmp := (OTHERS=>sel( 23));
      result := result or ( input_23 and tmp);
      tmp := (OTHERS=>sel( 24));
      result := result or ( input_24 and tmp);
      tmp := (OTHERS=>sel( 25));
      result := result or ( input_25 and tmp);
      tmp := (OTHERS=>sel( 26));
      result := result or ( input_26 and tmp);
      tmp := (OTHERS=>sel( 27));
      result := result or ( input_27 and tmp);
      tmp := (OTHERS=>sel( 28));
      result := result or ( input_28 and tmp);
      tmp := (OTHERS=>sel( 29));
      result := result or ( input_29 and tmp);
      tmp := (OTHERS=>sel( 30));
      result := result or ( input_30 and tmp);
      tmp := (OTHERS=>sel( 31));
      result := result or ( input_31 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_32_3_2(input_2 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_32_4_2(input_3 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_32_5_2(input_4 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(4 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_32_6_2(input_5 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(5 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_32_8_2(input_7 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(7 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_32_9_2(input_8 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(8 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_3_3_2(input_2 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(2 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(2 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_3_4_2(input_3 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(2 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(2 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_4_3_2(input_2 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(3 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(3 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_4_4_2(input_3 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(3 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(3 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_7_4_2(input_3 : STD_LOGIC_VECTOR(6 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(6 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(6 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(6 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(6 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(6 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
    RETURN result;
  END;

  FUNCTION MUX_s_1_2_2(input_0 : STD_LOGIC;
  input_1 : STD_LOGIC;
  sel : STD_LOGIC)
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_2_2_2(input_0 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(1 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_31_2_2(input_0 : STD_LOGIC_VECTOR(30 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(30 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(30 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_3_2_2(input_0 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(2 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_4_2_2(input_0 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(3 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_7_2_2(input_0 : STD_LOGIC_VECTOR(6 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(6 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(6 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  p_rsci : work.ccs_in_pkg_v1.ccs_in_v1
    GENERIC MAP(
      rscid => 2,
      width => 32
      )
    PORT MAP(
      dat => p_rsci_dat,
      idat => p_rsci_idat_1
    );
  p_rsci_dat <= p_rsc_dat;
  p_rsci_idat <= p_rsci_idat_1;

  xt_rsc_triosy_7_31_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_7_31_lz
    );
  xt_rsc_triosy_7_30_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_7_30_lz
    );
  xt_rsc_triosy_7_29_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_7_29_lz
    );
  xt_rsc_triosy_7_28_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_7_28_lz
    );
  xt_rsc_triosy_7_27_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_7_27_lz
    );
  xt_rsc_triosy_7_26_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_7_26_lz
    );
  xt_rsc_triosy_7_25_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_7_25_lz
    );
  xt_rsc_triosy_7_24_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_7_24_lz
    );
  xt_rsc_triosy_7_23_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_7_23_lz
    );
  xt_rsc_triosy_7_22_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_7_22_lz
    );
  xt_rsc_triosy_7_21_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_7_21_lz
    );
  xt_rsc_triosy_7_20_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_7_20_lz
    );
  xt_rsc_triosy_7_19_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_7_19_lz
    );
  xt_rsc_triosy_7_18_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_7_18_lz
    );
  xt_rsc_triosy_7_17_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_7_17_lz
    );
  xt_rsc_triosy_7_16_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_7_16_lz
    );
  xt_rsc_triosy_7_15_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_7_15_lz
    );
  xt_rsc_triosy_7_14_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_7_14_lz
    );
  xt_rsc_triosy_7_13_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_7_13_lz
    );
  xt_rsc_triosy_7_12_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_7_12_lz
    );
  xt_rsc_triosy_7_11_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_7_11_lz
    );
  xt_rsc_triosy_7_10_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_7_10_lz
    );
  xt_rsc_triosy_7_9_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_7_9_lz
    );
  xt_rsc_triosy_7_8_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_7_8_lz
    );
  xt_rsc_triosy_7_7_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_7_7_lz
    );
  xt_rsc_triosy_7_6_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_7_6_lz
    );
  xt_rsc_triosy_7_5_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_7_5_lz
    );
  xt_rsc_triosy_7_4_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_7_4_lz
    );
  xt_rsc_triosy_7_3_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_7_3_lz
    );
  xt_rsc_triosy_7_2_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_7_2_lz
    );
  xt_rsc_triosy_7_1_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_7_1_lz
    );
  xt_rsc_triosy_7_0_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_7_0_lz
    );
  xt_rsc_triosy_6_31_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_6_31_lz
    );
  xt_rsc_triosy_6_30_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_6_30_lz
    );
  xt_rsc_triosy_6_29_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_6_29_lz
    );
  xt_rsc_triosy_6_28_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_6_28_lz
    );
  xt_rsc_triosy_6_27_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_6_27_lz
    );
  xt_rsc_triosy_6_26_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_6_26_lz
    );
  xt_rsc_triosy_6_25_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_6_25_lz
    );
  xt_rsc_triosy_6_24_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_6_24_lz
    );
  xt_rsc_triosy_6_23_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_6_23_lz
    );
  xt_rsc_triosy_6_22_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_6_22_lz
    );
  xt_rsc_triosy_6_21_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_6_21_lz
    );
  xt_rsc_triosy_6_20_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_6_20_lz
    );
  xt_rsc_triosy_6_19_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_6_19_lz
    );
  xt_rsc_triosy_6_18_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_6_18_lz
    );
  xt_rsc_triosy_6_17_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_6_17_lz
    );
  xt_rsc_triosy_6_16_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_6_16_lz
    );
  xt_rsc_triosy_6_15_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_6_15_lz
    );
  xt_rsc_triosy_6_14_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_6_14_lz
    );
  xt_rsc_triosy_6_13_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_6_13_lz
    );
  xt_rsc_triosy_6_12_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_6_12_lz
    );
  xt_rsc_triosy_6_11_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_6_11_lz
    );
  xt_rsc_triosy_6_10_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_6_10_lz
    );
  xt_rsc_triosy_6_9_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_6_9_lz
    );
  xt_rsc_triosy_6_8_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_6_8_lz
    );
  xt_rsc_triosy_6_7_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_6_7_lz
    );
  xt_rsc_triosy_6_6_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_6_6_lz
    );
  xt_rsc_triosy_6_5_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_6_5_lz
    );
  xt_rsc_triosy_6_4_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_6_4_lz
    );
  xt_rsc_triosy_6_3_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_6_3_lz
    );
  xt_rsc_triosy_6_2_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_6_2_lz
    );
  xt_rsc_triosy_6_1_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_6_1_lz
    );
  xt_rsc_triosy_6_0_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_6_0_lz
    );
  xt_rsc_triosy_5_31_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_5_31_lz
    );
  xt_rsc_triosy_5_30_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_5_30_lz
    );
  xt_rsc_triosy_5_29_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_5_29_lz
    );
  xt_rsc_triosy_5_28_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_5_28_lz
    );
  xt_rsc_triosy_5_27_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_5_27_lz
    );
  xt_rsc_triosy_5_26_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_5_26_lz
    );
  xt_rsc_triosy_5_25_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_5_25_lz
    );
  xt_rsc_triosy_5_24_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_5_24_lz
    );
  xt_rsc_triosy_5_23_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_5_23_lz
    );
  xt_rsc_triosy_5_22_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_5_22_lz
    );
  xt_rsc_triosy_5_21_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_5_21_lz
    );
  xt_rsc_triosy_5_20_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_5_20_lz
    );
  xt_rsc_triosy_5_19_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_5_19_lz
    );
  xt_rsc_triosy_5_18_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_5_18_lz
    );
  xt_rsc_triosy_5_17_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_5_17_lz
    );
  xt_rsc_triosy_5_16_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_5_16_lz
    );
  xt_rsc_triosy_5_15_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_5_15_lz
    );
  xt_rsc_triosy_5_14_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_5_14_lz
    );
  xt_rsc_triosy_5_13_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_5_13_lz
    );
  xt_rsc_triosy_5_12_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_5_12_lz
    );
  xt_rsc_triosy_5_11_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_5_11_lz
    );
  xt_rsc_triosy_5_10_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_5_10_lz
    );
  xt_rsc_triosy_5_9_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_5_9_lz
    );
  xt_rsc_triosy_5_8_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_5_8_lz
    );
  xt_rsc_triosy_5_7_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_5_7_lz
    );
  xt_rsc_triosy_5_6_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_5_6_lz
    );
  xt_rsc_triosy_5_5_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_5_5_lz
    );
  xt_rsc_triosy_5_4_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_5_4_lz
    );
  xt_rsc_triosy_5_3_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_5_3_lz
    );
  xt_rsc_triosy_5_2_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_5_2_lz
    );
  xt_rsc_triosy_5_1_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_5_1_lz
    );
  xt_rsc_triosy_5_0_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_5_0_lz
    );
  xt_rsc_triosy_4_31_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_4_31_lz
    );
  xt_rsc_triosy_4_30_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_4_30_lz
    );
  xt_rsc_triosy_4_29_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_4_29_lz
    );
  xt_rsc_triosy_4_28_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_4_28_lz
    );
  xt_rsc_triosy_4_27_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_4_27_lz
    );
  xt_rsc_triosy_4_26_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_4_26_lz
    );
  xt_rsc_triosy_4_25_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_4_25_lz
    );
  xt_rsc_triosy_4_24_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_4_24_lz
    );
  xt_rsc_triosy_4_23_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_4_23_lz
    );
  xt_rsc_triosy_4_22_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_4_22_lz
    );
  xt_rsc_triosy_4_21_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_4_21_lz
    );
  xt_rsc_triosy_4_20_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_4_20_lz
    );
  xt_rsc_triosy_4_19_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_4_19_lz
    );
  xt_rsc_triosy_4_18_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_4_18_lz
    );
  xt_rsc_triosy_4_17_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_4_17_lz
    );
  xt_rsc_triosy_4_16_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_4_16_lz
    );
  xt_rsc_triosy_4_15_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_4_15_lz
    );
  xt_rsc_triosy_4_14_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_4_14_lz
    );
  xt_rsc_triosy_4_13_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_4_13_lz
    );
  xt_rsc_triosy_4_12_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_4_12_lz
    );
  xt_rsc_triosy_4_11_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_4_11_lz
    );
  xt_rsc_triosy_4_10_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_4_10_lz
    );
  xt_rsc_triosy_4_9_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_4_9_lz
    );
  xt_rsc_triosy_4_8_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_4_8_lz
    );
  xt_rsc_triosy_4_7_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_4_7_lz
    );
  xt_rsc_triosy_4_6_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_4_6_lz
    );
  xt_rsc_triosy_4_5_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_4_5_lz
    );
  xt_rsc_triosy_4_4_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_4_4_lz
    );
  xt_rsc_triosy_4_3_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_4_3_lz
    );
  xt_rsc_triosy_4_2_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_4_2_lz
    );
  xt_rsc_triosy_4_1_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_4_1_lz
    );
  xt_rsc_triosy_4_0_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_4_0_lz
    );
  xt_rsc_triosy_3_31_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_3_31_lz
    );
  xt_rsc_triosy_3_30_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_3_30_lz
    );
  xt_rsc_triosy_3_29_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_3_29_lz
    );
  xt_rsc_triosy_3_28_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_3_28_lz
    );
  xt_rsc_triosy_3_27_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_3_27_lz
    );
  xt_rsc_triosy_3_26_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_3_26_lz
    );
  xt_rsc_triosy_3_25_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_3_25_lz
    );
  xt_rsc_triosy_3_24_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_3_24_lz
    );
  xt_rsc_triosy_3_23_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_3_23_lz
    );
  xt_rsc_triosy_3_22_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_3_22_lz
    );
  xt_rsc_triosy_3_21_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_3_21_lz
    );
  xt_rsc_triosy_3_20_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_3_20_lz
    );
  xt_rsc_triosy_3_19_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_3_19_lz
    );
  xt_rsc_triosy_3_18_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_3_18_lz
    );
  xt_rsc_triosy_3_17_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_3_17_lz
    );
  xt_rsc_triosy_3_16_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_3_16_lz
    );
  xt_rsc_triosy_3_15_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_3_15_lz
    );
  xt_rsc_triosy_3_14_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_3_14_lz
    );
  xt_rsc_triosy_3_13_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_3_13_lz
    );
  xt_rsc_triosy_3_12_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_3_12_lz
    );
  xt_rsc_triosy_3_11_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_3_11_lz
    );
  xt_rsc_triosy_3_10_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_3_10_lz
    );
  xt_rsc_triosy_3_9_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_3_9_lz
    );
  xt_rsc_triosy_3_8_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_3_8_lz
    );
  xt_rsc_triosy_3_7_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_3_7_lz
    );
  xt_rsc_triosy_3_6_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_3_6_lz
    );
  xt_rsc_triosy_3_5_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_3_5_lz
    );
  xt_rsc_triosy_3_4_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_3_4_lz
    );
  xt_rsc_triosy_3_3_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_3_3_lz
    );
  xt_rsc_triosy_3_2_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_3_2_lz
    );
  xt_rsc_triosy_3_1_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_3_1_lz
    );
  xt_rsc_triosy_3_0_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_3_0_lz
    );
  xt_rsc_triosy_2_31_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_2_31_lz
    );
  xt_rsc_triosy_2_30_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_2_30_lz
    );
  xt_rsc_triosy_2_29_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_2_29_lz
    );
  xt_rsc_triosy_2_28_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_2_28_lz
    );
  xt_rsc_triosy_2_27_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_2_27_lz
    );
  xt_rsc_triosy_2_26_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_2_26_lz
    );
  xt_rsc_triosy_2_25_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_2_25_lz
    );
  xt_rsc_triosy_2_24_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_2_24_lz
    );
  xt_rsc_triosy_2_23_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_2_23_lz
    );
  xt_rsc_triosy_2_22_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_2_22_lz
    );
  xt_rsc_triosy_2_21_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_2_21_lz
    );
  xt_rsc_triosy_2_20_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_2_20_lz
    );
  xt_rsc_triosy_2_19_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_2_19_lz
    );
  xt_rsc_triosy_2_18_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_2_18_lz
    );
  xt_rsc_triosy_2_17_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_2_17_lz
    );
  xt_rsc_triosy_2_16_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_2_16_lz
    );
  xt_rsc_triosy_2_15_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_2_15_lz
    );
  xt_rsc_triosy_2_14_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_2_14_lz
    );
  xt_rsc_triosy_2_13_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_2_13_lz
    );
  xt_rsc_triosy_2_12_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_2_12_lz
    );
  xt_rsc_triosy_2_11_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_2_11_lz
    );
  xt_rsc_triosy_2_10_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_2_10_lz
    );
  xt_rsc_triosy_2_9_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_2_9_lz
    );
  xt_rsc_triosy_2_8_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_2_8_lz
    );
  xt_rsc_triosy_2_7_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_2_7_lz
    );
  xt_rsc_triosy_2_6_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_2_6_lz
    );
  xt_rsc_triosy_2_5_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_2_5_lz
    );
  xt_rsc_triosy_2_4_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_2_4_lz
    );
  xt_rsc_triosy_2_3_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_2_3_lz
    );
  xt_rsc_triosy_2_2_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_2_2_lz
    );
  xt_rsc_triosy_2_1_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_2_1_lz
    );
  xt_rsc_triosy_2_0_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_2_0_lz
    );
  xt_rsc_triosy_1_31_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_1_31_lz
    );
  xt_rsc_triosy_1_30_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_1_30_lz
    );
  xt_rsc_triosy_1_29_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_1_29_lz
    );
  xt_rsc_triosy_1_28_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_1_28_lz
    );
  xt_rsc_triosy_1_27_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_1_27_lz
    );
  xt_rsc_triosy_1_26_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_1_26_lz
    );
  xt_rsc_triosy_1_25_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_1_25_lz
    );
  xt_rsc_triosy_1_24_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_1_24_lz
    );
  xt_rsc_triosy_1_23_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_1_23_lz
    );
  xt_rsc_triosy_1_22_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_1_22_lz
    );
  xt_rsc_triosy_1_21_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_1_21_lz
    );
  xt_rsc_triosy_1_20_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_1_20_lz
    );
  xt_rsc_triosy_1_19_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_1_19_lz
    );
  xt_rsc_triosy_1_18_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_1_18_lz
    );
  xt_rsc_triosy_1_17_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_1_17_lz
    );
  xt_rsc_triosy_1_16_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_1_16_lz
    );
  xt_rsc_triosy_1_15_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_1_15_lz
    );
  xt_rsc_triosy_1_14_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_1_14_lz
    );
  xt_rsc_triosy_1_13_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_1_13_lz
    );
  xt_rsc_triosy_1_12_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_1_12_lz
    );
  xt_rsc_triosy_1_11_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_1_11_lz
    );
  xt_rsc_triosy_1_10_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_1_10_lz
    );
  xt_rsc_triosy_1_9_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_1_9_lz
    );
  xt_rsc_triosy_1_8_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_1_8_lz
    );
  xt_rsc_triosy_1_7_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_1_7_lz
    );
  xt_rsc_triosy_1_6_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_1_6_lz
    );
  xt_rsc_triosy_1_5_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_1_5_lz
    );
  xt_rsc_triosy_1_4_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_1_4_lz
    );
  xt_rsc_triosy_1_3_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_1_3_lz
    );
  xt_rsc_triosy_1_2_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_1_2_lz
    );
  xt_rsc_triosy_1_1_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_1_1_lz
    );
  xt_rsc_triosy_1_0_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_1_0_lz
    );
  xt_rsc_triosy_0_31_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_0_31_lz
    );
  xt_rsc_triosy_0_30_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_0_30_lz
    );
  xt_rsc_triosy_0_29_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_0_29_lz
    );
  xt_rsc_triosy_0_28_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_0_28_lz
    );
  xt_rsc_triosy_0_27_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_0_27_lz
    );
  xt_rsc_triosy_0_26_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_0_26_lz
    );
  xt_rsc_triosy_0_25_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_0_25_lz
    );
  xt_rsc_triosy_0_24_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_0_24_lz
    );
  xt_rsc_triosy_0_23_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_0_23_lz
    );
  xt_rsc_triosy_0_22_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_0_22_lz
    );
  xt_rsc_triosy_0_21_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_0_21_lz
    );
  xt_rsc_triosy_0_20_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_0_20_lz
    );
  xt_rsc_triosy_0_19_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_0_19_lz
    );
  xt_rsc_triosy_0_18_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_0_18_lz
    );
  xt_rsc_triosy_0_17_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_0_17_lz
    );
  xt_rsc_triosy_0_16_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_0_16_lz
    );
  xt_rsc_triosy_0_15_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_0_15_lz
    );
  xt_rsc_triosy_0_14_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_0_14_lz
    );
  xt_rsc_triosy_0_13_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_0_13_lz
    );
  xt_rsc_triosy_0_12_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_0_12_lz
    );
  xt_rsc_triosy_0_11_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_0_11_lz
    );
  xt_rsc_triosy_0_10_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_0_10_lz
    );
  xt_rsc_triosy_0_9_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_0_9_lz
    );
  xt_rsc_triosy_0_8_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_0_8_lz
    );
  xt_rsc_triosy_0_7_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_0_7_lz
    );
  xt_rsc_triosy_0_6_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_0_6_lz
    );
  xt_rsc_triosy_0_5_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_0_5_lz
    );
  xt_rsc_triosy_0_4_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_0_4_lz
    );
  xt_rsc_triosy_0_3_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_0_3_lz
    );
  xt_rsc_triosy_0_2_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_0_2_lz
    );
  xt_rsc_triosy_0_1_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_0_1_lz
    );
  xt_rsc_triosy_0_0_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => xt_rsc_triosy_0_0_lz
    );
  p_rsc_triosy_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => p_rsc_triosy_lz
    );
  r_rsc_triosy_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => r_rsc_triosy_lz
    );
  twiddle_rsc_triosy_0_15_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_15_lz
    );
  twiddle_rsc_triosy_0_14_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_14_lz
    );
  twiddle_rsc_triosy_0_13_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_13_lz
    );
  twiddle_rsc_triosy_0_12_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_12_lz
    );
  twiddle_rsc_triosy_0_11_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_11_lz
    );
  twiddle_rsc_triosy_0_10_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_10_lz
    );
  twiddle_rsc_triosy_0_9_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_9_lz
    );
  twiddle_rsc_triosy_0_8_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_8_lz
    );
  twiddle_rsc_triosy_0_7_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_7_lz
    );
  twiddle_rsc_triosy_0_6_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_6_lz
    );
  twiddle_rsc_triosy_0_5_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_5_lz
    );
  twiddle_rsc_triosy_0_4_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_4_lz
    );
  twiddle_rsc_triosy_0_3_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_3_lz
    );
  twiddle_rsc_triosy_0_2_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_2_lz
    );
  twiddle_rsc_triosy_0_1_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_1_lz
    );
  twiddle_rsc_triosy_0_0_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_0_lz
    );
  twiddle_h_rsc_triosy_0_15_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => twiddle_h_rsc_triosy_0_15_lz
    );
  twiddle_h_rsc_triosy_0_14_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => twiddle_h_rsc_triosy_0_14_lz
    );
  twiddle_h_rsc_triosy_0_13_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => twiddle_h_rsc_triosy_0_13_lz
    );
  twiddle_h_rsc_triosy_0_12_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => twiddle_h_rsc_triosy_0_12_lz
    );
  twiddle_h_rsc_triosy_0_11_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => twiddle_h_rsc_triosy_0_11_lz
    );
  twiddle_h_rsc_triosy_0_10_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => twiddle_h_rsc_triosy_0_10_lz
    );
  twiddle_h_rsc_triosy_0_9_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => twiddle_h_rsc_triosy_0_9_lz
    );
  twiddle_h_rsc_triosy_0_8_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => twiddle_h_rsc_triosy_0_8_lz
    );
  twiddle_h_rsc_triosy_0_7_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => twiddle_h_rsc_triosy_0_7_lz
    );
  twiddle_h_rsc_triosy_0_6_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => twiddle_h_rsc_triosy_0_6_lz
    );
  twiddle_h_rsc_triosy_0_5_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => twiddle_h_rsc_triosy_0_5_lz
    );
  twiddle_h_rsc_triosy_0_4_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => twiddle_h_rsc_triosy_0_4_lz
    );
  twiddle_h_rsc_triosy_0_3_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => twiddle_h_rsc_triosy_0_3_lz
    );
  twiddle_h_rsc_triosy_0_2_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => twiddle_h_rsc_triosy_0_2_lz
    );
  twiddle_h_rsc_triosy_0_1_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => twiddle_h_rsc_triosy_0_1_lz
    );
  twiddle_h_rsc_triosy_0_0_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_7_31_obj_ld_cse,
      lz => twiddle_h_rsc_triosy_0_0_lz
    );
  mult_t_mul_cmp : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 64,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_t_mul_cmp_a,
      b => mult_t_mul_cmp_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_t_mul_cmp_z_1
    );
  mult_t_mul_cmp_a <= MUX1HOT_v_32_4_2(z_out_43, z_out_59, z_out_49, z_out_35, STD_LOGIC_VECTOR'(
      (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  mult_t_mul_cmp_b <= MUX1HOT_v_32_9_2((twiddle_h_rsc_0_0_i_qa_d(31 DOWNTO 0)), (twiddle_h_rsc_0_8_i_qa_d(31
      DOWNTO 0)), (twiddle_h_rsc_0_9_i_qa_d(31 DOWNTO 0)), (twiddle_h_rsc_0_10_i_qa_d(31
      DOWNTO 0)), (twiddle_h_rsc_0_11_i_qa_d(31 DOWNTO 0)), (twiddle_h_rsc_0_12_i_qa_d(31
      DOWNTO 0)), (twiddle_h_rsc_0_13_i_qa_d(31 DOWNTO 0)), (twiddle_h_rsc_0_14_i_qa_d(31
      DOWNTO 0)), (twiddle_h_rsc_0_15_i_qa_d(31 DOWNTO 0)), STD_LOGIC_VECTOR'( modulo_add_1_qelse_or_m1c
      & mult_15_t_and_44_cse & mult_15_t_and_45_cse & mult_15_t_and_46_cse & mult_15_t_and_47_cse
      & mult_15_t_or_9_cse & mult_15_t_or_10_cse & mult_15_t_or_11_cse & mult_15_t_or_12_cse));
  mult_t_mul_cmp_z <= mult_t_mul_cmp_z_1;

  mult_t_mul_cmp_1 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 64,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_t_mul_cmp_1_a,
      b => mult_t_mul_cmp_1_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_t_mul_cmp_1_z_1
    );
  mult_t_mul_cmp_1_a <= MUX1HOT_v_32_4_2(z_out_49, z_out_35, z_out_42, z_out_59,
      STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  mult_t_mul_cmp_1_b <= MUX1HOT_v_32_5_2((twiddle_h_rsc_0_0_i_qa_d(31 DOWNTO 0)),
      (twiddle_h_rsc_0_8_i_qa_d(31 DOWNTO 0)), (twiddle_h_rsc_0_10_i_qa_d(31 DOWNTO
      0)), (twiddle_h_rsc_0_12_i_qa_d(31 DOWNTO 0)), (twiddle_h_rsc_0_14_i_qa_d(31
      DOWNTO 0)), STD_LOGIC_VECTOR'( or_tmp_3231 & mult_15_t_and_40_cse & mult_15_t_and_41_cse
      & mult_15_t_and_42_cse & mult_15_t_and_43_cse));
  mult_t_mul_cmp_1_z <= mult_t_mul_cmp_1_z_1;

  mult_t_mul_cmp_2 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 64,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_t_mul_cmp_2_a,
      b => mult_t_mul_cmp_2_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_t_mul_cmp_2_z_1
    );
  mult_t_mul_cmp_2_a <= MUX1HOT_v_32_4_2(z_out_42, z_out_50, z_out_41, z_out_32,
      STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  mult_t_mul_cmp_2_b <= MUX1HOT_v_32_6_2((twiddle_h_rsc_0_0_i_qa_d(31 DOWNTO 0)),
      (twiddle_h_rsc_0_8_i_qa_d(31 DOWNTO 0)), (twiddle_h_rsc_0_9_i_qa_d(31 DOWNTO
      0)), (twiddle_h_rsc_0_12_i_qa_d(31 DOWNTO 0)), (twiddle_h_rsc_0_13_i_qa_d(31
      DOWNTO 0)), (twiddle_h_rsc_0_1_i_qa_d(31 DOWNTO 0)), STD_LOGIC_VECTOR'( or_tmp_3239
      & mult_15_t_and_36_cse & mult_15_t_and_37_cse & mult_15_t_and_38_cse & mult_15_t_and_39_cse
      & or_tmp_3242));
  mult_t_mul_cmp_2_z <= mult_t_mul_cmp_2_z_1;

  mult_t_mul_cmp_3 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 64,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_t_mul_cmp_3_a,
      b => mult_t_mul_cmp_3_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_t_mul_cmp_3_z_1
    );
  mult_t_mul_cmp_3_a <= MUX1HOT_v_32_4_2(z_out_41, z_out_51, z_out_40, z_out_33,
      STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  mult_t_mul_cmp_3_b <= MUX1HOT_v_32_4_2((twiddle_h_rsc_0_0_i_qa_d(31 DOWNTO 0)),
      (twiddle_h_rsc_0_12_i_qa_d(31 DOWNTO 0)), (twiddle_h_rsc_0_8_i_qa_d(31 DOWNTO
      0)), (twiddle_h_rsc_0_2_i_qa_d(31 DOWNTO 0)), STD_LOGIC_VECTOR'( (and_7109_cse
      OR modulo_add_1_qelse_or_m1c) & or_tmp_3250 & and_7115_cse & or_tmp_3252));
  mult_t_mul_cmp_3_z <= mult_t_mul_cmp_3_z_1;

  mult_t_mul_cmp_4 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 64,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_t_mul_cmp_4_a,
      b => mult_t_mul_cmp_4_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_t_mul_cmp_4_z_1
    );
  mult_t_mul_cmp_4_a <= MUX1HOT_v_32_4_2(z_out_40, z_out_52, z_out_39, z_out_34,
      STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  mult_t_mul_cmp_4_b <= MUX1HOT_v_32_8_2((twiddle_h_rsc_0_0_i_qa_d(31 DOWNTO 0)),
      (twiddle_h_rsc_0_8_i_qa_d(31 DOWNTO 0)), (twiddle_h_rsc_0_9_i_qa_d(31 DOWNTO
      0)), (twiddle_h_rsc_0_10_i_qa_d(31 DOWNTO 0)), (twiddle_h_rsc_0_11_i_qa_d(31
      DOWNTO 0)), (twiddle_h_rsc_0_1_i_qa_d(31 DOWNTO 0)), (twiddle_h_rsc_0_2_i_qa_d(31
      DOWNTO 0)), (twiddle_h_rsc_0_3_i_qa_d(31 DOWNTO 0)), STD_LOGIC_VECTOR'( (modulo_add_1_qelse_or_m1c
      OR mult_15_t_and_49_cse) & mult_15_t_and_29_cse & mult_15_t_and_30_cse & mult_15_t_and_31_cse
      & mult_15_t_and_32_cse & mult_15_t_and_51_cse & mult_15_t_and_53_cse & mult_15_t_and_55_cse));
  mult_t_mul_cmp_4_z <= mult_t_mul_cmp_4_z_1;

  mult_t_mul_cmp_5 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 64,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_t_mul_cmp_5_a,
      b => mult_t_mul_cmp_5_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_t_mul_cmp_5_z_1
    );
  mult_t_mul_cmp_5_a <= MUX1HOT_v_32_4_2(z_out_39, mult_t_mul_cmp_5_a_mx0w1, z_out_38,
      mult_t_mul_cmp_5_a_mx0w4, STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4))
      & (fsm_output(7)) & (fsm_output(9))));
  mult_t_mul_cmp_5_b <= MUX1HOT_v_32_4_2((twiddle_h_rsc_0_0_i_qa_d(31 DOWNTO 0)),
      (twiddle_h_rsc_0_10_i_qa_d(31 DOWNTO 0)), (twiddle_h_rsc_0_8_i_qa_d(31 DOWNTO
      0)), (twiddle_h_rsc_0_4_i_qa_d(31 DOWNTO 0)), STD_LOGIC_VECTOR'( modulo_add_1_qelse_or_m1c
      & or_tmp_3269 & and_7153_cse & (fsm_output(9))));
  mult_t_mul_cmp_5_z <= mult_t_mul_cmp_5_z_1;

  mult_t_mul_cmp_6 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 64,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_t_mul_cmp_6_a,
      b => mult_t_mul_cmp_6_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_t_mul_cmp_6_z_1
    );
  mult_t_mul_cmp_6_a <= MUX1HOT_v_32_4_2(z_out_38, z_out_53, z_out_37, z_out_54,
      STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  mult_t_mul_cmp_6_b <= MUX1HOT_v_32_5_2((twiddle_h_rsc_0_0_i_qa_d(31 DOWNTO 0)),
      (twiddle_h_rsc_0_9_i_qa_d(31 DOWNTO 0)), (twiddle_h_rsc_0_8_i_qa_d(31 DOWNTO
      0)), (twiddle_h_rsc_0_5_i_qa_d(31 DOWNTO 0)), (twiddle_h_rsc_0_4_i_qa_d(31
      DOWNTO 0)), STD_LOGIC_VECTOR'( modulo_add_1_qelse_or_m1c & or_tmp_3279 & and_7173_cse
      & or_tmp_3242 & and_7090_cse));
  mult_t_mul_cmp_6_z <= mult_t_mul_cmp_6_z_1;

  mult_t_mul_cmp_7 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 64,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_t_mul_cmp_7_a,
      b => mult_t_mul_cmp_7_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_t_mul_cmp_7_z_1
    );
  mult_t_mul_cmp_7_a <= MUX1HOT_v_32_4_2(z_out_37, z_out_55, z_out_48, z_out_56,
      STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  mult_t_mul_cmp_7_b <= MUX1HOT_v_32_4_2((twiddle_h_rsc_0_0_i_qa_d(31 DOWNTO 0)),
      (twiddle_h_rsc_0_8_i_qa_d(31 DOWNTO 0)), (twiddle_h_rsc_0_6_i_qa_d(31 DOWNTO
      0)), (twiddle_h_rsc_0_4_i_qa_d(31 DOWNTO 0)), STD_LOGIC_VECTOR'( modulo_add_1_qelse_or_m1c
      & (fsm_output(7)) & or_tmp_3252 & and_7109_cse));
  mult_t_mul_cmp_7_z <= mult_t_mul_cmp_7_z_1;

  mult_t_mul_cmp_8 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 64,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_t_mul_cmp_8_a,
      b => mult_t_mul_cmp_8_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_t_mul_cmp_8_z_1
    );
  mult_t_mul_cmp_8_a <= MUX1HOT_v_32_4_2(z_out_48, z_out_57, z_out_47, z_out_58,
      STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  mult_t_mul_cmp_8_b <= MUX1HOT_v_32_8_2((twiddle_h_rsc_0_0_i_qa_d(31 DOWNTO 0)),
      (twiddle_h_rsc_0_1_i_qa_d(31 DOWNTO 0)), (twiddle_h_rsc_0_2_i_qa_d(31 DOWNTO
      0)), (twiddle_h_rsc_0_3_i_qa_d(31 DOWNTO 0)), (twiddle_h_rsc_0_4_i_qa_d(31
      DOWNTO 0)), (twiddle_h_rsc_0_5_i_qa_d(31 DOWNTO 0)), (twiddle_h_rsc_0_6_i_qa_d(31
      DOWNTO 0)), (twiddle_h_rsc_0_7_i_qa_d(31 DOWNTO 0)), STD_LOGIC_VECTOR'( mult_15_t_or_3_cse
      & mult_15_t_and_45_cse & mult_15_t_and_46_cse & mult_15_t_and_47_cse & mult_15_t_or_9_cse
      & mult_15_t_or_10_cse & mult_15_t_or_11_cse & mult_15_t_or_12_cse));
  mult_t_mul_cmp_8_z <= mult_t_mul_cmp_8_z_1;

  mult_t_mul_cmp_9 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 64,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_t_mul_cmp_9_a,
      b => mult_t_mul_cmp_9_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_t_mul_cmp_9_z_1
    );
  mult_t_mul_cmp_9_a <= MUX1HOT_v_32_4_2(z_out_47, z_out_58, z_out_46, z_out_57,
      STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  mult_t_mul_cmp_9_b <= MUX1HOT_v_32_5_2((twiddle_h_rsc_0_0_i_qa_d(31 DOWNTO 0)),
      (twiddle_h_rsc_0_2_i_qa_d(31 DOWNTO 0)), (twiddle_h_rsc_0_4_i_qa_d(31 DOWNTO
      0)), (twiddle_h_rsc_0_6_i_qa_d(31 DOWNTO 0)), (twiddle_h_rsc_0_8_i_qa_d(31
      DOWNTO 0)), STD_LOGIC_VECTOR'( (modulo_add_1_qelse_or_m1c OR mult_15_t_and_40_cse)
      & mult_15_t_and_41_cse & mult_15_t_and_42_cse & mult_15_t_and_43_cse & (fsm_output(9))));
  mult_t_mul_cmp_9_z <= mult_t_mul_cmp_9_z_1;

  mult_t_mul_cmp_10 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 64,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_t_mul_cmp_10_a,
      b => mult_t_mul_cmp_10_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_t_mul_cmp_10_z_1
    );
  mult_t_mul_cmp_10_a <= MUX1HOT_v_32_4_2(z_out_46, z_out_56, z_out_36, z_out_55,
      STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  mult_t_mul_cmp_10_b <= MUX1HOT_v_32_6_2((twiddle_h_rsc_0_0_i_qa_d(31 DOWNTO 0)),
      (twiddle_h_rsc_0_1_i_qa_d(31 DOWNTO 0)), (twiddle_h_rsc_0_4_i_qa_d(31 DOWNTO
      0)), (twiddle_h_rsc_0_5_i_qa_d(31 DOWNTO 0)), (twiddle_h_rsc_0_9_i_qa_d(31
      DOWNTO 0)), (twiddle_h_rsc_0_8_i_qa_d(31 DOWNTO 0)), STD_LOGIC_VECTOR'( mult_15_t_or_1_cse
      & mult_15_t_and_37_cse & mult_15_t_and_38_cse & mult_15_t_and_39_cse & or_tmp_3242
      & and_7090_cse));
  mult_t_mul_cmp_10_z <= mult_t_mul_cmp_10_z_1;

  mult_t_mul_cmp_11 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 64,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_t_mul_cmp_11_a,
      b => mult_t_mul_cmp_11_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_t_mul_cmp_11_z_1
    );
  mult_t_mul_cmp_11_a <= MUX1HOT_v_32_4_2(z_out_36, z_out_54, mult_t_mul_cmp_11_a_mx0w3,
      z_out_53, STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7))
      & (fsm_output(9))));
  mult_t_mul_cmp_11_b <= MUX1HOT_v_32_4_2((twiddle_h_rsc_0_0_i_qa_d(31 DOWNTO 0)),
      (twiddle_h_rsc_0_4_i_qa_d(31 DOWNTO 0)), (twiddle_h_rsc_0_10_i_qa_d(31 DOWNTO
      0)), (twiddle_h_rsc_0_8_i_qa_d(31 DOWNTO 0)), STD_LOGIC_VECTOR'( (and_7115_cse
      OR modulo_add_1_qelse_or_m1c) & or_tmp_3250 & or_tmp_3252 & and_7109_cse));
  mult_t_mul_cmp_11_z <= mult_t_mul_cmp_11_z_1;

  mult_t_mul_cmp_12 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 64,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_t_mul_cmp_12_a,
      b => mult_t_mul_cmp_12_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_t_mul_cmp_12_z_1
    );
  mult_t_mul_cmp_12_a <= mult_4_t_mux1h_1_rmff;
  mult_t_mul_cmp_12_b <= MUX1HOT_v_32_8_2((twiddle_h_rsc_0_0_i_qa_d(31 DOWNTO 0)),
      (twiddle_h_rsc_0_1_i_qa_d(31 DOWNTO 0)), (twiddle_h_rsc_0_2_i_qa_d(31 DOWNTO
      0)), (twiddle_h_rsc_0_3_i_qa_d(31 DOWNTO 0)), (twiddle_h_rsc_0_8_i_qa_d(31
      DOWNTO 0)), (twiddle_h_rsc_0_9_i_qa_d(31 DOWNTO 0)), (twiddle_h_rsc_0_10_i_qa_d(31
      DOWNTO 0)), (twiddle_h_rsc_0_11_i_qa_d(31 DOWNTO 0)), STD_LOGIC_VECTOR'( mult_15_t_or_cse
      & mult_15_t_and_30_cse & mult_15_t_and_31_cse & mult_15_t_and_32_cse & mult_15_t_and_49_cse
      & mult_15_t_and_51_cse & mult_15_t_and_53_cse & mult_15_t_and_55_cse));
  mult_t_mul_cmp_12_z <= mult_t_mul_cmp_12_z_1;

  mult_t_mul_cmp_13 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 64,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_t_mul_cmp_13_a,
      b => mult_t_mul_cmp_13_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_t_mul_cmp_13_z_1
    );
  mult_t_mul_cmp_13_a <= MUX1HOT_v_32_4_2(tmp_71_lpi_3_dfm_1, z_out_34, z_out_45,
      z_out_52, STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7))
      & (fsm_output(9))));
  mult_t_mul_cmp_13_b <= MUX1HOT_v_32_3_2((twiddle_h_rsc_0_0_i_qa_d(31 DOWNTO 0)),
      (twiddle_h_rsc_0_2_i_qa_d(31 DOWNTO 0)), (twiddle_h_rsc_0_12_i_qa_d(31 DOWNTO
      0)), STD_LOGIC_VECTOR'( or_tmp_3345 & or_tmp_3269 & (fsm_output(9))));
  mult_t_mul_cmp_13_z <= mult_t_mul_cmp_13_z_1;

  mult_t_mul_cmp_14 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 64,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_t_mul_cmp_14_a,
      b => mult_t_mul_cmp_14_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_t_mul_cmp_14_z_1
    );
  mult_t_mul_cmp_14_a <= MUX1HOT_v_32_4_2(z_out_45, z_out_33, z_out_44, z_out_51,
      STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  mult_t_mul_cmp_14_b <= MUX1HOT_v_32_4_2((twiddle_h_rsc_0_0_i_qa_d(31 DOWNTO 0)),
      (twiddle_h_rsc_0_1_i_qa_d(31 DOWNTO 0)), (twiddle_h_rsc_0_13_i_qa_d(31 DOWNTO
      0)), (twiddle_h_rsc_0_12_i_qa_d(31 DOWNTO 0)), STD_LOGIC_VECTOR'( or_tmp_3354
      & or_tmp_3279 & or_tmp_3242 & and_7090_cse));
  mult_t_mul_cmp_14_z <= mult_t_mul_cmp_14_z_1;

  mult_t_mul_cmp_15 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 64,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_t_mul_cmp_15_a,
      b => mult_t_mul_cmp_15_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_t_mul_cmp_15_z_1
    );
  mult_t_mul_cmp_15_a <= MUX1HOT_v_32_4_2(z_out_44, z_out_32, z_out_43, z_out_50,
      STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  mult_t_mul_cmp_15_b <= MUX1HOT_v_32_3_2((twiddle_h_rsc_0_0_i_qa_d(31 DOWNTO 0)),
      (twiddle_h_rsc_0_14_i_qa_d(31 DOWNTO 0)), (twiddle_h_rsc_0_12_i_qa_d(31 DOWNTO
      0)), STD_LOGIC_VECTOR'( (modulo_add_1_qelse_or_m1c OR (fsm_output(7))) & or_tmp_3252
      & and_7109_cse));
  mult_t_mul_cmp_15_z <= mult_t_mul_cmp_15_z_1;

  mult_z_mul_cmp : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_z_mul_cmp_a,
      b => mult_z_mul_cmp_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_z_1
    );
  mult_z_mul_cmp_a <= MUX1HOT_v_32_3_2(z_out_43, z_out_59, z_out_49, STD_LOGIC_VECTOR'(
      (fsm_output(2)) & ((fsm_output(4)) OR (fsm_output(9))) & (fsm_output(7))));
  mult_z_mul_cmp_b <= MUX1HOT_v_32_9_2((twiddle_rsc_0_0_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_8_i_qa_d(31
      DOWNTO 0)), (twiddle_rsc_0_9_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_10_i_qa_d(31
      DOWNTO 0)), (twiddle_rsc_0_11_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_12_i_qa_d(31
      DOWNTO 0)), (twiddle_rsc_0_13_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_14_i_qa_d(31
      DOWNTO 0)), (twiddle_rsc_0_15_i_qa_d(31 DOWNTO 0)), STD_LOGIC_VECTOR'( or_tmp_3231
      & mult_15_t_and_44_cse & mult_15_t_and_45_cse & mult_15_t_and_46_cse & mult_15_t_and_47_cse
      & mult_15_t_and_48_cse & mult_15_t_and_50_cse & mult_15_t_and_52_cse & mult_15_t_and_54_cse));
  mult_z_mul_cmp_z <= mult_z_mul_cmp_z_1;

  mult_z_mul_cmp_1 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_z_mul_cmp_1_a,
      b => mult_z_mul_cmp_1_b,
      clk => clk,
      en => mult_z_mul_cmp_1_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_1_z_1
    );
  mult_z_mul_cmp_1_a <= MUX1HOT_v_32_3_2((mult_t_mul_cmp_1_z(63 DOWNTO 32)), (mult_t_mul_cmp_11_z(63
      DOWNTO 32)), (mult_t_mul_cmp_12_z(63 DOWNTO 32)), STD_LOGIC_VECTOR'( modulo_add_1_qelse_or_m1c
      & (fsm_output(7)) & (fsm_output(9))));
  mult_z_mul_cmp_1_b <= p_sva;
  mult_z_mul_cmp_1_z <= mult_z_mul_cmp_1_z_1;

  mult_z_mul_cmp_2 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_z_mul_cmp_2_a,
      b => mult_z_mul_cmp_2_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_2_z_1
    );
  mult_z_mul_cmp_2_a <= MUX1HOT_v_32_4_2(z_out_49, z_out_35, z_out_43, z_out_57,
      STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  mult_z_mul_cmp_2_b <= MUX_v_32_2_2((twiddle_rsc_0_0_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_8_i_qa_d(31
      DOWNTO 0)), fsm_output(9));
  mult_z_mul_cmp_2_z <= mult_z_mul_cmp_2_z_1;

  mult_z_mul_cmp_3 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_z_mul_cmp_3_a,
      b => mult_z_mul_cmp_3_b,
      clk => clk,
      en => mult_z_mul_cmp_1_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_3_z_1
    );
  mult_z_mul_cmp_3_a <= MUX1HOT_v_32_3_2((mult_t_mul_cmp_2_z(63 DOWNTO 32)), (mult_t_mul_cmp_5_z(63
      DOWNTO 32)), (mult_t_mul_cmp_6_z(63 DOWNTO 32)), STD_LOGIC_VECTOR'( modulo_add_1_qelse_or_m1c
      & (fsm_output(7)) & (fsm_output(9))));
  mult_z_mul_cmp_3_b <= p_sva;
  mult_z_mul_cmp_3_z <= mult_z_mul_cmp_3_z_1;

  mult_z_mul_cmp_4 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_z_mul_cmp_4_a,
      b => mult_z_mul_cmp_4_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_4_z_1
    );
  mult_z_mul_cmp_4_a <= MUX1HOT_v_32_3_2(z_out_42, z_out_50, mult_t_mul_cmp_5_a_mx0w4,
      STD_LOGIC_VECTOR'( ((fsm_output(2)) OR (fsm_output(7))) & (fsm_output(4)) &
      (fsm_output(9))));
  mult_z_mul_cmp_4_b <= MUX1HOT_v_32_6_2((twiddle_rsc_0_0_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_8_i_qa_d(31
      DOWNTO 0)), (twiddle_rsc_0_10_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_12_i_qa_d(31
      DOWNTO 0)), (twiddle_rsc_0_14_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_4_i_qa_d(31
      DOWNTO 0)), STD_LOGIC_VECTOR'( modulo_add_1_qelse_or_m1c & mult_15_t_and_40_cse
      & mult_15_t_and_41_cse & mult_15_t_and_42_cse & mult_15_t_and_43_cse & (fsm_output(9))));
  mult_z_mul_cmp_4_z <= mult_z_mul_cmp_4_z_1;

  mult_z_mul_cmp_5 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_z_mul_cmp_5_a,
      b => mult_z_mul_cmp_5_b,
      clk => clk,
      en => mult_z_mul_cmp_1_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_5_z_1
    );
  mult_z_mul_cmp_5_a <= MUX1HOT_v_32_3_2((mult_t_mul_cmp_3_z(63 DOWNTO 32)), (mult_t_mul_cmp_12_z(63
      DOWNTO 32)), (mult_t_mul_cmp_13_z(63 DOWNTO 32)), STD_LOGIC_VECTOR'( modulo_add_1_qelse_or_m1c
      & (fsm_output(7)) & (fsm_output(9))));
  mult_z_mul_cmp_5_b <= p_sva;
  mult_z_mul_cmp_5_z <= mult_z_mul_cmp_5_z_1;

  mult_z_mul_cmp_6 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_z_mul_cmp_6_a,
      b => mult_z_mul_cmp_6_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_6_z_1
    );
  mult_z_mul_cmp_6_a <= MUX1HOT_v_32_4_2(z_out_41, z_out_51, z_out_47, z_out_35,
      STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  mult_z_mul_cmp_6_b <= MUX1HOT_v_32_12_2((twiddle_rsc_0_0_i_qa_d(31 DOWNTO 0)),
      (twiddle_rsc_0_1_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_2_i_qa_d(31 DOWNTO 0)),
      (twiddle_rsc_0_3_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_4_i_qa_d(31 DOWNTO 0)),
      (twiddle_rsc_0_5_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_6_i_qa_d(31 DOWNTO 0)),
      (twiddle_rsc_0_7_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_12_i_qa_d(31 DOWNTO 0)),
      (twiddle_rsc_0_13_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_14_i_qa_d(31 DOWNTO
      0)), (twiddle_rsc_0_15_i_qa_d(31 DOWNTO 0)), STD_LOGIC_VECTOR'( mult_15_t_or_3_cse
      & mult_15_t_and_45_cse & mult_15_t_and_46_cse & mult_15_t_and_47_cse & mult_15_t_and_48_cse
      & mult_15_t_and_50_cse & mult_15_t_and_52_cse & mult_15_t_and_54_cse & mult_15_t_and_49_cse
      & mult_15_t_and_51_cse & mult_15_t_and_53_cse & mult_15_t_and_55_cse));
  mult_z_mul_cmp_6_z <= mult_z_mul_cmp_6_z_1;

  mult_z_mul_cmp_7 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_z_mul_cmp_7_a,
      b => mult_z_mul_cmp_7_b,
      clk => clk,
      en => mult_z_mul_cmp_1_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_7_z_1
    );
  mult_z_mul_cmp_7_a <= MUX1HOT_v_32_3_2((mult_t_mul_cmp_4_z(63 DOWNTO 32)), (mult_t_mul_cmp_2_z(63
      DOWNTO 32)), (mult_t_mul_cmp_3_z(63 DOWNTO 32)), STD_LOGIC_VECTOR'( modulo_add_1_qelse_or_m1c
      & (fsm_output(7)) & (fsm_output(9))));
  mult_z_mul_cmp_7_b <= p_sva;
  mult_z_mul_cmp_7_z <= mult_z_mul_cmp_7_z_1;

  mult_z_mul_cmp_8 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_z_mul_cmp_8_a,
      b => mult_z_mul_cmp_8_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_8_z_1
    );
  mult_z_mul_cmp_8_a <= MUX1HOT_v_32_4_2(z_out_40, z_out_52, z_out_44, z_out_55,
      STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  mult_z_mul_cmp_8_b <= MUX1HOT_v_32_4_2((twiddle_rsc_0_0_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_1_i_qa_d(31
      DOWNTO 0)), (twiddle_rsc_0_9_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_8_i_qa_d(31
      DOWNTO 0)), STD_LOGIC_VECTOR'( or_tmp_3354 & or_tmp_3279 & or_tmp_3242 & and_7090_cse));
  mult_z_mul_cmp_8_z <= mult_z_mul_cmp_8_z_1;

  mult_z_mul_cmp_9 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_z_mul_cmp_9_a,
      b => mult_z_mul_cmp_9_b,
      clk => clk,
      en => mult_z_mul_cmp_1_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_9_z_1
    );
  mult_z_mul_cmp_9_a <= MUX1HOT_v_32_3_2((mult_t_mul_cmp_5_z(63 DOWNTO 32)), (mult_t_mul_cmp_10_z(63
      DOWNTO 32)), (mult_t_mul_cmp_11_z(63 DOWNTO 32)), STD_LOGIC_VECTOR'( modulo_add_1_qelse_or_m1c
      & (fsm_output(7)) & (fsm_output(9))));
  mult_z_mul_cmp_9_b <= p_sva;
  mult_z_mul_cmp_9_z <= mult_z_mul_cmp_9_z_1;

  mult_z_mul_cmp_10 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_z_mul_cmp_10_a,
      b => mult_z_mul_cmp_10_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_10_z_1
    );
  mult_z_mul_cmp_10_a <= MUX1HOT_v_32_4_2(z_out_39, mult_t_mul_cmp_5_a_mx0w1, z_out_48,
      z_out_58, STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7))
      & (fsm_output(9))));
  mult_z_mul_cmp_10_b <= MUX1HOT_v_32_6_2((twiddle_rsc_0_0_i_qa_d(31 DOWNTO 0)),
      (twiddle_rsc_0_8_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_4_i_qa_d(31 DOWNTO 0)),
      (twiddle_rsc_0_5_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_6_i_qa_d(31 DOWNTO 0)),
      (twiddle_rsc_0_7_i_qa_d(31 DOWNTO 0)), STD_LOGIC_VECTOR'( modulo_add_1_qelse_or_m1c
      & (fsm_output(7)) & mult_15_t_and_49_cse & mult_15_t_and_51_cse & mult_15_t_and_53_cse
      & mult_15_t_and_55_cse));
  mult_z_mul_cmp_10_z <= mult_z_mul_cmp_10_z_1;

  mult_z_mul_cmp_11 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_z_mul_cmp_11_a,
      b => mult_z_mul_cmp_11_b,
      clk => clk,
      en => mult_z_mul_cmp_1_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_11_z_1
    );
  mult_z_mul_cmp_11_a <= MUX_v_32_2_2((mult_t_mul_cmp_6_z(63 DOWNTO 32)), (mult_t_mul_cmp_7_z(63
      DOWNTO 32)), fsm_output(9));
  mult_z_mul_cmp_11_b <= p_sva;
  mult_z_mul_cmp_11_z <= mult_z_mul_cmp_11_z_1;

  mult_z_mul_cmp_12 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_z_mul_cmp_12_a,
      b => mult_z_mul_cmp_12_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_12_z_1
    );
  mult_z_mul_cmp_12_a <= MUX1HOT_v_32_4_2(z_out_38, z_out_53, z_out_45, z_out_34,
      STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  mult_z_mul_cmp_12_b <= MUX1HOT_v_32_4_2((twiddle_rsc_0_0_i_qa_d(31 DOWNTO 0)),
      (twiddle_rsc_0_2_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_1_i_qa_d(31 DOWNTO 0)),
      (twiddle_rsc_0_3_i_qa_d(31 DOWNTO 0)), STD_LOGIC_VECTOR'( (or_tmp_3345 OR mult_15_t_and_49_cse)
      & (or_tmp_3269 OR mult_15_t_and_53_cse) & mult_15_t_and_51_cse & mult_15_t_and_55_cse));
  mult_z_mul_cmp_12_z <= mult_z_mul_cmp_12_z_1;

  mult_z_mul_cmp_13 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_z_mul_cmp_13_a,
      b => mult_z_mul_cmp_13_b,
      clk => clk,
      en => mult_z_mul_cmp_1_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_13_z_1
    );
  mult_z_mul_cmp_13_a <= MUX1HOT_v_32_3_2((mult_t_mul_cmp_7_z(63 DOWNTO 32)), (mult_t_mul_cmp_1_z(63
      DOWNTO 32)), (mult_t_mul_cmp_2_z(63 DOWNTO 32)), STD_LOGIC_VECTOR'( modulo_add_1_qelse_or_m1c
      & (fsm_output(7)) & (fsm_output(9))));
  mult_z_mul_cmp_13_b <= p_sva;
  mult_z_mul_cmp_13_z <= mult_z_mul_cmp_13_z_1;

  mult_z_mul_cmp_14 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_z_mul_cmp_14_a,
      b => mult_z_mul_cmp_14_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_14_z_1
    );
  mult_z_mul_cmp_14_a <= MUX1HOT_v_32_4_2(z_out_37, z_out_55, z_out_41, z_out_50,
      STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  mult_z_mul_cmp_14_b <= MUX1HOT_v_32_6_2((twiddle_rsc_0_0_i_qa_d(31 DOWNTO 0)),
      (twiddle_rsc_0_8_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_9_i_qa_d(31 DOWNTO 0)),
      (twiddle_rsc_0_12_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_13_i_qa_d(31 DOWNTO
      0)), (twiddle_rsc_0_14_i_qa_d(31 DOWNTO 0)), STD_LOGIC_VECTOR'( modulo_add_1_qelse_or_m1c
      & mult_15_t_and_36_cse & mult_15_t_and_37_cse & (mult_15_t_and_38_cse OR and_7109_cse)
      & mult_15_t_and_39_cse & or_tmp_3252));
  mult_z_mul_cmp_14_z <= mult_z_mul_cmp_14_z_1;

  mult_z_mul_cmp_15 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_z_mul_cmp_15_a,
      b => mult_z_mul_cmp_15_b,
      clk => clk,
      en => mult_z_mul_cmp_1_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_15_z_1
    );
  mult_z_mul_cmp_15_a <= MUX1HOT_v_32_3_2((mult_t_mul_cmp_8_z(63 DOWNTO 32)), (mult_t_mul_cmp_13_z(63
      DOWNTO 32)), (mult_t_mul_cmp_14_z(63 DOWNTO 32)), STD_LOGIC_VECTOR'( modulo_add_1_qelse_or_m1c
      & (fsm_output(7)) & (fsm_output(9))));
  mult_z_mul_cmp_15_b <= p_sva;
  mult_z_mul_cmp_15_z <= mult_z_mul_cmp_15_z_1;

  mult_z_mul_cmp_16 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_z_mul_cmp_16_a,
      b => mult_z_mul_cmp_16_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_16_z_1
    );
  mult_z_mul_cmp_16_a <= MUX1HOT_v_32_4_2(z_out_48, z_out_57, z_out_46, z_out_32,
      STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  mult_z_mul_cmp_16_b <= MUX1HOT_v_32_5_2((twiddle_rsc_0_0_i_qa_d(31 DOWNTO 0)),
      (twiddle_rsc_0_2_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_4_i_qa_d(31 DOWNTO 0)),
      (twiddle_rsc_0_6_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_1_i_qa_d(31 DOWNTO 0)),
      STD_LOGIC_VECTOR'( (or_tmp_3239 OR mult_15_t_and_40_cse) & mult_15_t_and_41_cse
      & mult_15_t_and_42_cse & mult_15_t_and_43_cse & or_tmp_3242));
  mult_z_mul_cmp_16_z <= mult_z_mul_cmp_16_z_1;

  mult_z_mul_cmp_17 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_z_mul_cmp_17_a,
      b => mult_z_mul_cmp_17_b,
      clk => clk,
      en => mult_z_mul_cmp_1_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_17_z_1
    );
  mult_z_mul_cmp_17_a <= MUX_v_32_2_2((mult_t_mul_cmp_9_z(63 DOWNTO 32)), (mult_t_mul_cmp_10_z(63
      DOWNTO 32)), fsm_output(9));
  mult_z_mul_cmp_17_b <= p_sva;
  mult_z_mul_cmp_17_z <= mult_z_mul_cmp_17_z_1;

  mult_z_mul_cmp_18 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_z_mul_cmp_18_a,
      b => mult_z_mul_cmp_18_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_18_z_1
    );
  mult_z_mul_cmp_18_a <= MUX1HOT_v_32_4_2(z_out_47, z_out_58, z_out_37, z_out_53,
      STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  mult_z_mul_cmp_18_b <= MUX1HOT_v_32_4_2((twiddle_rsc_0_0_i_qa_d(31 DOWNTO 0)),
      (twiddle_rsc_0_9_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_8_i_qa_d(31 DOWNTO 0)),
      (twiddle_rsc_0_10_i_qa_d(31 DOWNTO 0)), STD_LOGIC_VECTOR'( modulo_add_1_qelse_or_m1c
      & or_tmp_3279 & (and_7173_cse OR and_7109_cse) & or_tmp_3252));
  mult_z_mul_cmp_18_z <= mult_z_mul_cmp_18_z_1;

  mult_z_mul_cmp_19 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_z_mul_cmp_19_a,
      b => mult_z_mul_cmp_19_b,
      clk => clk,
      en => mult_z_mul_cmp_1_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_19_z_1
    );
  mult_z_mul_cmp_19_a <= MUX1HOT_v_32_3_2((mult_t_mul_cmp_10_z(63 DOWNTO 32)), (mult_t_mul_cmp_4_z(63
      DOWNTO 32)), (mult_t_mul_cmp_5_z(63 DOWNTO 32)), STD_LOGIC_VECTOR'( modulo_add_1_qelse_or_m1c
      & (fsm_output(7)) & (fsm_output(9))));
  mult_z_mul_cmp_19_b <= p_sva;
  mult_z_mul_cmp_19_z <= mult_z_mul_cmp_19_z_1;

  mult_z_mul_cmp_20 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_z_mul_cmp_20_a,
      b => mult_z_mul_cmp_20_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_20_z_1
    );
  mult_z_mul_cmp_20_a <= MUX1HOT_v_32_4_2(z_out_46, z_out_56, z_out_40, z_out_54,
      STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  mult_z_mul_cmp_20_b <= MUX1HOT_v_32_5_2((twiddle_rsc_0_0_i_qa_d(31 DOWNTO 0)),
      (twiddle_rsc_0_12_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_8_i_qa_d(31 DOWNTO 0)),
      (twiddle_rsc_0_5_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_4_i_qa_d(31 DOWNTO 0)),
      STD_LOGIC_VECTOR'( modulo_add_1_qelse_or_m1c & or_tmp_3250 & and_7115_cse &
      or_tmp_3242 & and_7090_cse));
  mult_z_mul_cmp_20_z <= mult_z_mul_cmp_20_z_1;

  mult_z_mul_cmp_21 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_z_mul_cmp_21_a,
      b => mult_z_mul_cmp_21_b,
      clk => clk,
      en => mult_z_mul_cmp_1_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_21_z_1
    );
  mult_z_mul_cmp_21_a <= MUX1HOT_v_32_3_2((mult_t_mul_cmp_11_z(63 DOWNTO 32)), (mult_t_mul_cmp_14_z(63
      DOWNTO 32)), (mult_t_mul_cmp_15_z(63 DOWNTO 32)), STD_LOGIC_VECTOR'( modulo_add_1_qelse_or_m1c
      & (fsm_output(7)) & (fsm_output(9))));
  mult_z_mul_cmp_21_b <= p_sva;
  mult_z_mul_cmp_21_z <= mult_z_mul_cmp_21_z_1;

  mult_z_mul_cmp_22 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_z_mul_cmp_22_a,
      b => mult_z_mul_cmp_22_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_22_z_1
    );
  mult_z_mul_cmp_22_a <= MUX1HOT_v_32_3_2(z_out_36, z_out_54, z_out_51, STD_LOGIC_VECTOR'(
      ((fsm_output(2)) OR (fsm_output(7))) & (fsm_output(4)) & (fsm_output(9))));
  mult_z_mul_cmp_22_b <= MUX1HOT_v_32_6_2((twiddle_rsc_0_0_i_qa_d(31 DOWNTO 0)),
      (twiddle_rsc_0_1_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_4_i_qa_d(31 DOWNTO 0)),
      (twiddle_rsc_0_5_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_13_i_qa_d(31 DOWNTO 0)),
      (twiddle_rsc_0_12_i_qa_d(31 DOWNTO 0)), STD_LOGIC_VECTOR'( mult_15_t_or_1_cse
      & mult_15_t_and_37_cse & mult_15_t_and_38_cse & mult_15_t_and_39_cse & or_tmp_3242
      & and_7090_cse));
  mult_z_mul_cmp_22_z <= mult_z_mul_cmp_22_z_1;

  mult_z_mul_cmp_23 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_z_mul_cmp_23_a,
      b => mult_z_mul_cmp_23_b,
      clk => clk,
      en => mult_z_mul_cmp_1_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_23_z_1
    );
  mult_z_mul_cmp_23_a <= MUX1HOT_v_32_3_2((mult_t_mul_cmp_12_z(63 DOWNTO 32)), (mult_t_mul_cmp_3_z(63
      DOWNTO 32)), (mult_t_mul_cmp_4_z(63 DOWNTO 32)), STD_LOGIC_VECTOR'( modulo_add_1_qelse_or_m1c
      & (fsm_output(7)) & (fsm_output(9))));
  mult_z_mul_cmp_23_b <= p_sva;
  mult_z_mul_cmp_23_z <= mult_z_mul_cmp_23_z_1;

  mult_z_mul_cmp_24 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_z_mul_cmp_24_a,
      b => mult_z_mul_cmp_24_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_24_z_1
    );
  mult_z_mul_cmp_24_a <= mult_4_t_mux1h_1_rmff;
  mult_z_mul_cmp_24_b <= MUX1HOT_v_32_8_2((twiddle_rsc_0_0_i_qa_d(31 DOWNTO 0)),
      (twiddle_rsc_0_1_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_2_i_qa_d(31 DOWNTO 0)),
      (twiddle_rsc_0_3_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_8_i_qa_d(31 DOWNTO 0)),
      (twiddle_rsc_0_9_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_10_i_qa_d(31 DOWNTO 0)),
      (twiddle_rsc_0_11_i_qa_d(31 DOWNTO 0)), STD_LOGIC_VECTOR'( mult_15_t_or_cse
      & mult_15_t_and_30_cse & mult_15_t_and_31_cse & mult_15_t_and_32_cse & mult_15_t_and_49_cse
      & mult_15_t_and_51_cse & mult_15_t_and_53_cse & mult_15_t_and_55_cse));
  mult_z_mul_cmp_24_z <= mult_z_mul_cmp_24_z_1;

  mult_z_mul_cmp_25 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_z_mul_cmp_25_a,
      b => mult_z_mul_cmp_25_b,
      clk => clk,
      en => mult_z_mul_cmp_1_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_25_z_1
    );
  mult_z_mul_cmp_25_a <= MUX1HOT_v_32_3_2((mult_t_mul_cmp_13_z(63 DOWNTO 32)), (mult_t_mul_cmp_8_z(63
      DOWNTO 32)), (mult_t_mul_cmp_9_z(63 DOWNTO 32)), STD_LOGIC_VECTOR'( modulo_add_1_qelse_or_m1c
      & (fsm_output(7)) & (fsm_output(9))));
  mult_z_mul_cmp_25_b <= p_sva;
  mult_z_mul_cmp_25_z <= mult_z_mul_cmp_25_z_1;

  mult_z_mul_cmp_26 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_z_mul_cmp_26_a,
      b => mult_z_mul_cmp_26_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_26_z_1
    );
  mult_z_mul_cmp_26_a <= MUX1HOT_v_32_4_2(tmp_71_lpi_3_dfm_1, z_out_34, z_out_38,
      z_out_56, STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7))
      & (fsm_output(9))));
  mult_z_mul_cmp_26_b <= MUX1HOT_v_32_5_2((twiddle_rsc_0_0_i_qa_d(31 DOWNTO 0)),
      (twiddle_rsc_0_10_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_8_i_qa_d(31 DOWNTO 0)),
      (twiddle_rsc_0_6_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_4_i_qa_d(31 DOWNTO 0)),
      STD_LOGIC_VECTOR'( modulo_add_1_qelse_or_m1c & or_tmp_3269 & and_7153_cse &
      or_tmp_3252 & and_7109_cse));
  mult_z_mul_cmp_26_z <= mult_z_mul_cmp_26_z_1;

  mult_z_mul_cmp_27 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_z_mul_cmp_27_a,
      b => mult_z_mul_cmp_27_b,
      clk => clk,
      en => mult_z_mul_cmp_1_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_27_z_1
    );
  mult_z_mul_cmp_27_a <= MUX1HOT_v_32_3_2((mult_t_mul_cmp_14_z(63 DOWNTO 32)), (mult_t_mul_cmp_7_z(63
      DOWNTO 32)), (mult_t_mul_cmp_8_z(63 DOWNTO 32)), STD_LOGIC_VECTOR'( modulo_add_1_qelse_or_m1c
      & (fsm_output(7)) & (fsm_output(9))));
  mult_z_mul_cmp_27_b <= p_sva;
  mult_z_mul_cmp_27_z <= mult_z_mul_cmp_27_z_1;

  mult_z_mul_cmp_28 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_z_mul_cmp_28_a,
      b => mult_z_mul_cmp_28_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_28_z_1
    );
  mult_z_mul_cmp_28_a <= MUX1HOT_v_32_3_2(z_out_45, z_out_33, mult_t_mul_cmp_11_a_mx0w3,
      STD_LOGIC_VECTOR'( (fsm_output(2)) & ((fsm_output(4)) OR (fsm_output(9))) &
      (fsm_output(7))));
  mult_z_mul_cmp_28_b <= MUX1HOT_v_32_3_2((twiddle_rsc_0_0_i_qa_d(31 DOWNTO 0)),
      (twiddle_rsc_0_4_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_2_i_qa_d(31 DOWNTO 0)),
      STD_LOGIC_VECTOR'( (and_7115_cse OR and_7109_cse OR modulo_add_1_qelse_or_m1c)
      & or_tmp_3250 & or_tmp_3252));
  mult_z_mul_cmp_28_z <= mult_z_mul_cmp_28_z_1;

  mult_z_mul_cmp_29 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_z_mul_cmp_29_a,
      b => mult_z_mul_cmp_29_b,
      clk => clk,
      en => mult_z_mul_cmp_1_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_29_z_1
    );
  mult_z_mul_cmp_29_a <= MUX1HOT_v_32_3_2((mult_t_mul_cmp_15_z(63 DOWNTO 32)), (mult_t_mul_cmp_z(63
      DOWNTO 32)), (mult_t_mul_cmp_1_z(63 DOWNTO 32)), STD_LOGIC_VECTOR'( modulo_add_1_qelse_or_m1c
      & (fsm_output(7)) & (fsm_output(9))));
  mult_z_mul_cmp_29_b <= p_sva;
  mult_z_mul_cmp_29_z <= mult_z_mul_cmp_29_z_1;

  mult_z_mul_cmp_30 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_z_mul_cmp_30_a,
      b => mult_z_mul_cmp_30_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_30_z_1
    );
  mult_z_mul_cmp_30_a <= MUX1HOT_v_32_4_2(z_out_44, z_out_32, z_out_39, z_out_52,
      STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  mult_z_mul_cmp_30_b <= MUX1HOT_v_32_6_2((twiddle_rsc_0_0_i_qa_d(31 DOWNTO 0)),
      (twiddle_rsc_0_8_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_9_i_qa_d(31 DOWNTO 0)),
      (twiddle_rsc_0_10_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_11_i_qa_d(31 DOWNTO
      0)), (twiddle_rsc_0_12_i_qa_d(31 DOWNTO 0)), STD_LOGIC_VECTOR'( modulo_add_1_qelse_or_m1c
      & mult_15_t_and_29_cse & mult_15_t_and_30_cse & mult_15_t_and_31_cse & mult_15_t_and_32_cse
      & (fsm_output(9))));
  mult_z_mul_cmp_30_z <= mult_z_mul_cmp_30_z_1;

  mult_z_mul_cmp_31 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_z_mul_cmp_31_a,
      b => mult_z_mul_cmp_31_b,
      clk => clk,
      en => mult_z_mul_cmp_1_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_31_z_1
    );
  mult_z_mul_cmp_31_a <= MUX_v_32_2_2((mult_t_mul_cmp_z(63 DOWNTO 32)), (mult_t_mul_cmp_15_z(63
      DOWNTO 32)), fsm_output(7));
  mult_z_mul_cmp_31_b <= p_sva;
  mult_z_mul_cmp_31_z <= mult_z_mul_cmp_31_z_1;

  operator_33_true_3_lshift_rg : work.mgc_shift_comps_v5.mgc_shift_bl_v5
    GENERIC MAP(
      width_a => 1,
      signd_a => 1,
      width_s => 3,
      width_z => 2
      )
    PORT MAP(
      a => operator_33_true_3_lshift_rg_a,
      s => operator_33_true_3_lshift_rg_s,
      z => operator_33_true_3_lshift_rg_z
    );
  operator_33_true_3_lshift_rg_a(0) <= '1';
  operator_33_true_3_lshift_rg_s <= STD_LOGIC_VECTOR'( '0' & (NOT c_1_sva) & '0');
  operator_33_true_3_lshift_psp_1_0_sva_mx0w5 <= operator_33_true_3_lshift_rg_z;

  operator_33_true_1_lshift_rg : work.mgc_shift_comps_v5.mgc_shift_l_v5
    GENERIC MAP(
      width_a => 1,
      signd_a => 1,
      width_s => 4,
      width_z => 11
      )
    PORT MAP(
      a => operator_33_true_1_lshift_rg_a,
      s => operator_33_true_1_lshift_rg_s,
      z => operator_33_true_1_lshift_rg_z
    );
  operator_33_true_1_lshift_rg_a(0) <= '1';
  operator_33_true_1_lshift_rg_s <= (MUX1HOT_v_3_3_2(z_out_61, operator_20_false_acc_cse_sva,
      (STD_LOGIC_VECTOR'( "00") & (NOT c_1_sva)), STD_LOGIC_VECTOR'( (fsm_output(1))
      & (fsm_output(3)) & (fsm_output(6))))) & ((NOT (fsm_output(3))) OR (fsm_output(1))
      OR (fsm_output(6)));
  z_out_60 <= operator_33_true_1_lshift_rg_z;

  peaseNTT_core_wait_dp_inst : peaseNTT_core_wait_dp
    PORT MAP(
      yt_rsc_0_0_cgo_iro => or_553_rmff,
      yt_rsc_0_0_i_clkr_en_d => yt_rsc_0_0_i_clkr_en_d,
      yt_rsc_0_16_cgo_iro => or_652_rmff,
      yt_rsc_0_16_i_clkr_en_d => yt_rsc_0_16_i_clkr_en_d,
      yt_rsc_1_0_cgo_iro => or_718_rmff,
      yt_rsc_1_0_i_clkr_en_d => yt_rsc_1_0_i_clkr_en_d,
      yt_rsc_1_16_cgo_iro => or_785_rmff,
      yt_rsc_1_16_i_clkr_en_d => yt_rsc_1_16_i_clkr_en_d,
      yt_rsc_2_0_cgo_iro => or_851_rmff,
      yt_rsc_2_0_i_clkr_en_d => yt_rsc_2_0_i_clkr_en_d,
      yt_rsc_2_16_cgo_iro => or_918_rmff,
      yt_rsc_2_16_i_clkr_en_d => yt_rsc_2_16_i_clkr_en_d,
      yt_rsc_3_0_cgo_iro => or_984_rmff,
      yt_rsc_3_0_i_clkr_en_d => yt_rsc_3_0_i_clkr_en_d,
      yt_rsc_3_16_cgo_iro => or_1051_rmff,
      yt_rsc_3_16_i_clkr_en_d => yt_rsc_3_16_i_clkr_en_d,
      yt_rsc_4_0_cgo_iro => or_1117_rmff,
      yt_rsc_4_0_i_clkr_en_d => yt_rsc_4_0_i_clkr_en_d,
      yt_rsc_4_16_cgo_iro => or_1216_rmff,
      yt_rsc_4_16_i_clkr_en_d => yt_rsc_4_16_i_clkr_en_d,
      yt_rsc_5_0_cgo_iro => or_1282_rmff,
      yt_rsc_5_0_i_clkr_en_d => yt_rsc_5_0_i_clkr_en_d,
      yt_rsc_5_16_cgo_iro => or_1349_rmff,
      yt_rsc_5_16_i_clkr_en_d => yt_rsc_5_16_i_clkr_en_d,
      yt_rsc_6_0_cgo_iro => or_1415_rmff,
      yt_rsc_6_0_i_clkr_en_d => yt_rsc_6_0_i_clkr_en_d,
      yt_rsc_6_16_cgo_iro => or_1482_rmff,
      yt_rsc_6_16_i_clkr_en_d => yt_rsc_6_16_i_clkr_en_d,
      yt_rsc_7_0_cgo_iro => or_1548_rmff,
      yt_rsc_7_0_i_clkr_en_d => yt_rsc_7_0_i_clkr_en_d,
      yt_rsc_7_16_cgo_iro => or_1615_rmff,
      yt_rsc_7_16_i_clkr_en_d => yt_rsc_7_16_i_clkr_en_d,
      ensig_cgo_iro => or_3599_rmff,
      ensig_cgo_iro_17 => or_3759_rmff,
      yt_rsc_0_0_cgo => reg_yt_rsc_0_0_cgo_cse,
      yt_rsc_0_16_cgo => reg_yt_rsc_0_16_cgo_cse,
      yt_rsc_1_0_cgo => reg_yt_rsc_1_0_cgo_cse,
      yt_rsc_1_16_cgo => reg_yt_rsc_1_16_cgo_cse,
      yt_rsc_2_0_cgo => reg_yt_rsc_2_0_cgo_cse,
      yt_rsc_2_16_cgo => reg_yt_rsc_2_16_cgo_cse,
      yt_rsc_3_0_cgo => reg_yt_rsc_3_0_cgo_cse,
      yt_rsc_3_16_cgo => reg_yt_rsc_3_16_cgo_cse,
      yt_rsc_4_0_cgo => reg_yt_rsc_4_0_cgo_cse,
      yt_rsc_4_16_cgo => reg_yt_rsc_4_16_cgo_cse,
      yt_rsc_5_0_cgo => reg_yt_rsc_5_0_cgo_cse,
      yt_rsc_5_16_cgo => reg_yt_rsc_5_16_cgo_cse,
      yt_rsc_6_0_cgo => reg_yt_rsc_6_0_cgo_cse,
      yt_rsc_6_16_cgo => reg_yt_rsc_6_16_cgo_cse,
      yt_rsc_7_0_cgo => reg_yt_rsc_7_0_cgo_cse,
      yt_rsc_7_16_cgo => reg_yt_rsc_7_16_cgo_cse,
      ensig_cgo => reg_ensig_cgo_cse,
      mult_t_mul_cmp_en => mult_t_mul_cmp_en,
      ensig_cgo_17 => reg_ensig_cgo_17_cse,
      mult_z_mul_cmp_1_en => mult_z_mul_cmp_1_en
    );
  peaseNTT_core_core_fsm_inst : peaseNTT_core_core_fsm
    PORT MAP(
      clk => clk,
      rst => rst,
      fsm_output => peaseNTT_core_core_fsm_inst_fsm_output,
      INNER_LOOP1_C_0_tr0 => peaseNTT_core_core_fsm_inst_INNER_LOOP1_C_0_tr0,
      INNER_LOOP2_C_0_tr0 => peaseNTT_core_core_fsm_inst_INNER_LOOP2_C_0_tr0,
      STAGE_LOOP_C_2_tr0 => peaseNTT_core_core_fsm_inst_STAGE_LOOP_C_2_tr0,
      INNER_LOOP3_C_0_tr0 => INNER_LOOP4_nor_tmp,
      INNER_LOOP4_C_0_tr0 => and_dcpl_62,
      INNER_LOOP4_C_0_tr1 => peaseNTT_core_core_fsm_inst_INNER_LOOP4_C_0_tr1
    );
  fsm_output <= peaseNTT_core_core_fsm_inst_fsm_output;
  peaseNTT_core_core_fsm_inst_INNER_LOOP1_C_0_tr0 <= NOT(INNER_LOOP1_stage_0 OR INNER_LOOP1_stage_0_2
      OR INNER_LOOP1_stage_0_3 OR butterFly2_15_conc_2_itm_0 OR butterFly2_15_conc_2_itm_1_0
      OR butterFly2_15_conc_2_itm_2_0 OR butterFly2_15_conc_2_itm_3_0 OR butterFly2_15_conc_2_itm_4_0
      OR butterFly2_15_conc_2_itm_5_0 OR INNER_LOOP1_stage_0_10);
  peaseNTT_core_core_fsm_inst_INNER_LOOP2_C_0_tr0 <= NOT(INNER_LOOP1_stage_0 OR butterFly2_15_conc_2_itm_7_0
      OR butterFly2_15_conc_2_itm_8_0 OR butterFly2_15_conc_2_itm_0 OR butterFly2_15_conc_2_itm_1_0
      OR butterFly2_15_conc_2_itm_2_0 OR butterFly2_15_conc_2_itm_3_0 OR butterFly2_15_conc_2_itm_4_0
      OR butterFly2_15_conc_2_itm_5_0 OR INNER_LOOP2_stage_0_10);
  peaseNTT_core_core_fsm_inst_STAGE_LOOP_C_2_tr0 <= z_out_61(2);
  peaseNTT_core_core_fsm_inst_INNER_LOOP4_C_0_tr1 <= NOT INNER_LOOP4_nor_tmp;

  or_4976_cse <= (fsm_output(10)) OR (fsm_output(0));
  mux_1_nl <= MUX_s_1_2_2(mux_tmp, or_tmp_26, butterFly2_15_conc_2_itm_9_2_1(0));
  or_322_nl <= CONV_SL_1_1(butterFly2_15_conc_2_itm_9_2_1/=STD_LOGIC_VECTOR'("00"))
      OR butterFly1_15_f1_equal_tmp_1_1 OR (NOT butterFly1_15_conc_2_itm_0);
  mux_2_nl <= MUX_s_1_2_2(mux_1_nl, or_322_nl, butterFly2_15_conc_itm_10_2_1(0));
  or_337_nl <= (butterFly1_15_conc_2_itm_9_2_1(0)) OR butterFly1_15_conc_2_itm_9_0
      OR (butterFly1_15_conc_2_itm_9_2_1(1));
  mux_5_nl <= MUX_s_1_2_2(not_tmp_29, or_tmp_40, or_337_nl);
  mux_6_nl <= MUX_s_1_2_2(mux_5_nl, or_tmp_38, butterFly2_15_conc_2_itm_6_2_1(0));
  or_553_rmff <= ((NOT mux_2_nl) AND (fsm_output(7))) OR and_344_cse OR ((NOT mux_6_nl)
      AND (fsm_output(2))) OR and_346_cse;
  mux_8_nl <= MUX_s_1_2_2(mux_tmp_7, or_tmp_48, butterFly2_15_conc_2_itm_9_2_1(0));
  or_344_nl <= CONV_SL_1_1(butterFly2_15_conc_2_itm_9_2_1/=STD_LOGIC_VECTOR'("00"))
      OR (NOT nor_tmp_1);
  mux_9_nl <= MUX_s_1_2_2(mux_8_nl, or_344_nl, butterFly2_15_conc_itm_10_2_1(0));
  or_352_nl <= (butterFly1_15_conc_2_itm_9_2_1(0)) OR (NOT butterFly1_15_conc_2_itm_9_0)
      OR (butterFly1_15_conc_2_itm_9_2_1(1));
  mux_10_nl <= MUX_s_1_2_2(not_tmp_50, or_tmp_55, or_352_nl);
  mux_11_nl <= MUX_s_1_2_2(mux_10_nl, or_tmp_53, butterFly2_15_conc_2_itm_6_2_1(0));
  or_652_rmff <= ((NOT mux_9_nl) AND (fsm_output(7))) OR and_344_cse OR ((NOT mux_11_nl)
      AND (fsm_output(2))) OR and_346_cse;
  or_356_nl <= CONV_SL_1_1(butterFly2_15_conc_2_itm_9_2_1/=STD_LOGIC_VECTOR'("01"))
      OR butterFly1_15_f1_equal_tmp_1_1 OR (NOT butterFly1_15_conc_2_itm_0);
  mux_12_nl <= MUX_s_1_2_2(or_tmp_26, mux_tmp, butterFly2_15_conc_2_itm_9_2_1(0));
  mux_13_nl <= MUX_s_1_2_2(or_356_nl, mux_12_nl, butterFly2_15_conc_itm_10_2_1(0));
  or_360_nl <= (NOT (butterFly1_15_conc_2_itm_9_2_1(0))) OR butterFly1_15_conc_2_itm_9_0
      OR (butterFly1_15_conc_2_itm_9_2_1(1));
  mux_16_nl <= MUX_s_1_2_2(not_tmp_29, or_tmp_40, or_360_nl);
  mux_17_nl <= MUX_s_1_2_2(or_tmp_64, mux_16_nl, butterFly2_15_conc_2_itm_6_2_1(0));
  or_718_rmff <= ((NOT mux_13_nl) AND (fsm_output(7))) OR and_715_cse OR ((NOT mux_17_nl)
      AND (fsm_output(2))) OR and_717_cse;
  or_367_nl <= CONV_SL_1_1(butterFly2_15_conc_2_itm_9_2_1/=STD_LOGIC_VECTOR'("01"))
      OR (NOT nor_tmp_1);
  mux_18_nl <= MUX_s_1_2_2(or_tmp_48, mux_tmp_7, butterFly2_15_conc_2_itm_9_2_1(0));
  mux_19_nl <= MUX_s_1_2_2(or_367_nl, mux_18_nl, butterFly2_15_conc_itm_10_2_1(0));
  or_368_nl <= (NOT (butterFly1_15_conc_2_itm_9_2_1(0))) OR (NOT butterFly1_15_conc_2_itm_9_0)
      OR (butterFly1_15_conc_2_itm_9_2_1(1));
  mux_20_nl <= MUX_s_1_2_2(not_tmp_50, or_tmp_55, or_368_nl);
  mux_21_nl <= MUX_s_1_2_2(or_tmp_72, mux_20_nl, butterFly2_15_conc_2_itm_6_2_1(0));
  or_785_rmff <= ((NOT mux_19_nl) AND (fsm_output(7))) OR and_715_cse OR ((NOT mux_21_nl)
      AND (fsm_output(2))) OR and_717_cse;
  mux_23_nl <= MUX_s_1_2_2(mux_tmp_22, or_tmp_75, butterFly2_15_conc_2_itm_9_2_1(0));
  or_372_nl <= CONV_SL_1_1(butterFly2_15_conc_2_itm_9_2_1/=STD_LOGIC_VECTOR'("10"))
      OR butterFly1_15_f1_equal_tmp_1_1 OR (NOT butterFly1_15_conc_2_itm_0);
  mux_24_nl <= MUX_s_1_2_2(mux_23_nl, or_372_nl, butterFly2_15_conc_itm_10_2_1(0));
  mux_27_nl <= MUX_s_1_2_2(not_tmp_67, or_tmp_86, or_383_cse);
  mux_28_nl <= MUX_s_1_2_2(mux_27_nl, or_tmp_84, butterFly2_15_conc_2_itm_6_2_1(0));
  or_851_rmff <= ((NOT mux_24_nl) AND (fsm_output(7))) OR and_1022_cse OR ((NOT mux_28_nl)
      AND (fsm_output(2))) OR and_1024_cse;
  mux_30_nl <= MUX_s_1_2_2(or_tmp_93, nor_tmp_15, butterFly2_15_conc_2_itm_9_2_1(0));
  nor_49_nl <= NOT((butterFly2_15_conc_2_itm_9_2_1(0)) OR (NOT nor_tmp_14));
  mux_31_nl <= MUX_s_1_2_2(mux_30_nl, nor_49_nl, butterFly2_15_conc_itm_10_2_1(0));
  nor_50_nl <= NOT(((NOT (butterFly1_15_conc_2_itm_9_2_1(0))) AND butterFly1_15_conc_2_itm_9_0
      AND (butterFly1_15_conc_2_itm_9_2_1(1)) AND INNER_LOOP1_stage_0_10) OR nor_tmp_19);
  mux_32_nl <= MUX_s_1_2_2(nor_50_nl, or_tmp_94, butterFly2_15_conc_2_itm_6_2_1(0));
  or_918_rmff <= (mux_31_nl AND (fsm_output(7))) OR and_1022_cse OR ((NOT mux_32_nl)
      AND (fsm_output(2))) OR and_1024_cse;
  nand_1_nl <= NOT(CONV_SL_1_1(butterFly2_15_conc_2_itm_9_2_1=STD_LOGIC_VECTOR'("11"))
      AND (NOT butterFly1_15_f1_equal_tmp_1_1) AND butterFly1_15_conc_2_itm_0);
  mux_33_nl <= MUX_s_1_2_2(or_tmp_75, mux_tmp_22, butterFly2_15_conc_2_itm_9_2_1(0));
  mux_34_nl <= MUX_s_1_2_2(nand_1_nl, mux_33_nl, butterFly2_15_conc_itm_10_2_1(0));
  mux_38_nl <= MUX_s_1_2_2(not_tmp_67, or_tmp_86, or_398_cse);
  mux_39_nl <= MUX_s_1_2_2(or_tmp_102, mux_38_nl, butterFly2_15_conc_2_itm_6_2_1(0));
  or_984_rmff <= ((NOT mux_34_nl) AND (fsm_output(7))) OR and_1329_cse OR ((NOT mux_39_nl)
      AND (fsm_output(2))) OR and_1331_cse;
  mux_41_nl <= MUX_s_1_2_2(nor_tmp_15, or_tmp_93, butterFly2_15_conc_2_itm_9_2_1(0));
  mux_42_nl <= MUX_s_1_2_2(nor_tmp_22, mux_41_nl, butterFly2_15_conc_itm_10_2_1(0));
  or_404_nl <= and_8913_cse OR nor_tmp_19;
  mux_43_nl <= MUX_s_1_2_2(and_8913_cse, or_404_nl, butterFly2_15_conc_2_itm_6_2_1(0));
  or_1051_rmff <= (mux_42_nl AND (fsm_output(7))) OR and_1329_cse OR (mux_43_nl AND
      (fsm_output(2))) OR and_1331_cse;
  mux_46_nl <= MUX_s_1_2_2(mux_tmp_45, or_tmp_29, butterFly2_15_conc_2_itm_8_2_1(0));
  or_406_nl <= CONV_SL_1_1(butterFly2_15_conc_2_itm_8_2_1/=STD_LOGIC_VECTOR'("00"))
      OR butterFly2_15_conc_2_itm_8_0 OR (NOT butterFly1_15_conc_2_itm_9_0);
  mux_47_nl <= MUX_s_1_2_2(mux_46_nl, or_406_nl, butterFly2_15_conc_2_itm_9_2_1(0));
  mux_51_nl <= MUX_s_1_2_2(mux_tmp_50, or_tmp_120, or_383_cse);
  mux_52_nl <= MUX_s_1_2_2(mux_51_nl, or_tmp_38, butterFly1_15_conc_2_itm_8_2_1(0));
  or_1117_rmff <= ((NOT mux_47_nl) AND (fsm_output(7))) OR and_1636_cse OR ((NOT
      mux_52_nl) AND (fsm_output(2))) OR and_1638_cse;
  mux_54_nl <= MUX_s_1_2_2(mux_tmp_53, or_tmp_50, butterFly2_15_conc_2_itm_8_2_1(0));
  or_426_nl <= CONV_SL_1_1(butterFly2_15_conc_2_itm_8_2_1/=STD_LOGIC_VECTOR'("00"))
      OR (NOT nor_tmp_25);
  mux_55_nl <= MUX_s_1_2_2(mux_54_nl, or_426_nl, butterFly2_15_conc_2_itm_9_2_1(0));
  mux_57_nl <= MUX_s_1_2_2(or_tmp_133, mux_tmp_56, nor_27_cse);
  mux_58_nl <= MUX_s_1_2_2(mux_57_nl, or_tmp_53, butterFly1_15_conc_2_itm_8_2_1(0));
  or_1216_rmff <= ((NOT mux_55_nl) AND (fsm_output(7))) OR and_1636_cse OR ((NOT
      mux_58_nl) AND (fsm_output(2))) OR and_1638_cse;
  or_433_nl <= CONV_SL_1_1(butterFly2_15_conc_2_itm_8_2_1/=STD_LOGIC_VECTOR'("01"))
      OR butterFly2_15_conc_2_itm_8_0 OR (NOT butterFly1_15_conc_2_itm_9_0);
  mux_59_nl <= MUX_s_1_2_2(or_tmp_29, mux_tmp_45, butterFly2_15_conc_2_itm_8_2_1(0));
  mux_60_nl <= MUX_s_1_2_2(or_433_nl, mux_59_nl, butterFly2_15_conc_2_itm_9_2_1(0));
  mux_63_nl <= MUX_s_1_2_2(mux_tmp_50, or_tmp_120, or_398_cse);
  mux_64_nl <= MUX_s_1_2_2(or_tmp_64, mux_63_nl, butterFly1_15_conc_2_itm_8_2_1(0));
  or_1282_rmff <= ((NOT mux_60_nl) AND (fsm_output(7))) OR and_2007_cse OR ((NOT
      mux_64_nl) AND (fsm_output(2))) OR and_2009_cse;
  or_442_nl <= CONV_SL_1_1(butterFly2_15_conc_2_itm_8_2_1/=STD_LOGIC_VECTOR'("01"))
      OR (NOT nor_tmp_25);
  mux_65_nl <= MUX_s_1_2_2(or_tmp_50, mux_tmp_53, butterFly2_15_conc_2_itm_8_2_1(0));
  mux_66_nl <= MUX_s_1_2_2(or_442_nl, mux_65_nl, butterFly2_15_conc_2_itm_9_2_1(0));
  mux_67_nl <= MUX_s_1_2_2(or_tmp_133, mux_tmp_56, and_8912_cse);
  mux_68_nl <= MUX_s_1_2_2(or_tmp_72, mux_67_nl, butterFly1_15_conc_2_itm_8_2_1(0));
  or_1349_rmff <= ((NOT mux_66_nl) AND (fsm_output(7))) OR and_2007_cse OR ((NOT
      mux_68_nl) AND (fsm_output(2))) OR and_2009_cse;
  mux_71_nl <= MUX_s_1_2_2(mux_tmp_70, or_tmp_77, butterFly2_15_conc_2_itm_8_2_1(0));
  or_444_nl <= CONV_SL_1_1(butterFly2_15_conc_2_itm_8_2_1/=STD_LOGIC_VECTOR'("10"))
      OR butterFly2_15_conc_2_itm_8_0 OR (NOT butterFly1_15_conc_2_itm_9_0);
  mux_72_nl <= MUX_s_1_2_2(mux_71_nl, or_444_nl, butterFly2_15_conc_2_itm_9_2_1(0));
  mux_75_nl <= MUX_s_1_2_2(not_tmp_115, or_tmp_153, or_383_cse);
  mux_76_nl <= MUX_s_1_2_2(mux_75_nl, or_tmp_84, butterFly1_15_conc_2_itm_8_2_1(0));
  or_1415_rmff <= ((NOT mux_72_nl) AND (fsm_output(7))) OR and_2314_cse OR ((NOT
      mux_76_nl) AND (fsm_output(2))) OR and_2316_cse;
  mux_79_nl <= MUX_s_1_2_2(mux_tmp_78, nor_tmp_14, butterFly2_15_conc_2_itm_8_2_1(0));
  nor_48_nl <= NOT((butterFly2_15_conc_2_itm_8_2_1(0)) OR (NOT nor_tmp_36));
  mux_80_nl <= MUX_s_1_2_2(mux_79_nl, nor_48_nl, butterFly2_15_conc_2_itm_9_2_1(0));
  mux_81_nl <= MUX_s_1_2_2(and_8919_cse, or_tmp_160, nor_27_cse);
  mux_82_nl <= MUX_s_1_2_2(mux_81_nl, (NOT or_tmp_94), butterFly1_15_conc_2_itm_8_2_1(0));
  or_1482_rmff <= (mux_80_nl AND (fsm_output(7))) OR and_2314_cse OR (mux_82_nl AND
      (fsm_output(2))) OR and_2316_cse;
  nand_nl <= NOT(CONV_SL_1_1(butterFly2_15_conc_2_itm_8_2_1=STD_LOGIC_VECTOR'("11"))
      AND (NOT butterFly2_15_conc_2_itm_8_0) AND butterFly1_15_conc_2_itm_9_0);
  mux_83_nl <= MUX_s_1_2_2(or_tmp_77, mux_tmp_70, butterFly2_15_conc_2_itm_8_2_1(0));
  mux_84_nl <= MUX_s_1_2_2(nand_nl, mux_83_nl, butterFly2_15_conc_2_itm_9_2_1(0));
  mux_87_nl <= MUX_s_1_2_2(not_tmp_115, or_tmp_153, or_398_cse);
  mux_88_nl <= MUX_s_1_2_2(or_tmp_102, mux_87_nl, butterFly1_15_conc_2_itm_8_2_1(0));
  or_1548_rmff <= ((NOT mux_84_nl) AND (fsm_output(7))) OR and_2621_cse OR ((NOT
      mux_88_nl) AND (fsm_output(2))) OR and_2623_cse;
  mux_89_nl <= MUX_s_1_2_2(nor_tmp_14, mux_tmp_78, butterFly2_15_conc_2_itm_8_2_1(0));
  mux_90_nl <= MUX_s_1_2_2(nor_tmp_46, mux_89_nl, butterFly2_15_conc_2_itm_9_2_1(0));
  mux_91_nl <= MUX_s_1_2_2(and_8919_cse, or_tmp_160, and_8912_cse);
  mux_92_nl <= MUX_s_1_2_2(and_8913_cse, mux_91_nl, butterFly1_15_conc_2_itm_8_2_1(0));
  or_1615_rmff <= (mux_90_nl AND (fsm_output(7))) OR and_2621_cse OR (mux_92_nl AND
      (fsm_output(2))) OR and_2623_cse;
  and_6824_rmff <= INNER_LOOP1_stage_0 AND or_dcpl_300;
  butterFly2_1_tw_butterFly2_1_tw_mux_rmff <= MUX_v_7_2_2(INNER_LOOP3_r_11_4_sva_6_0,
      INNER_LOOP4_r_11_4_sva_6_0, fsm_output(9));
  or_3498_rmff <= (and_dcpl_173 AND (fsm_output(7))) OR and_6834_cse;
  or_3502_rmff <= (and_dcpl_175 AND (fsm_output(7))) OR and_6843_cse;
  or_3506_rmff <= (and_dcpl_175 AND (operator_20_false_acc_cse_sva(0)) AND (fsm_output(7)))
      OR and_6852_cse;
  or_3510_rmff <= (INNER_LOOP1_stage_0 AND (operator_20_false_acc_cse_sva(2)) AND
      (fsm_output(7))) OR (INNER_LOOP1_stage_0 AND (fsm_output(9)));
  or_3514_rmff <= (and_dcpl_173 AND (operator_20_false_acc_cse_sva(2)) AND (fsm_output(7)))
      OR and_6834_cse;
  or_3518_rmff <= (and_dcpl_175 AND (operator_20_false_acc_cse_sva(2)) AND (fsm_output(7)))
      OR and_6843_cse;
  or_3522_rmff <= (and_dcpl_175 AND (operator_20_false_acc_cse_sva(0)) AND (operator_20_false_acc_cse_sva(2))
      AND (fsm_output(7))) OR and_6852_cse;
  and_6895_rmff <= INNER_LOOP1_stage_0 AND or_dcpl_298;
  or_3599_rmff <= ((butterFly1_15_conc_2_itm_2_0 OR butterFly1_15_conc_2_itm_4_0
      OR butterFly1_15_conc_2_itm_3_0) AND or_dcpl_298) OR ((INNER_LOOP1_stage_0_3
      OR INNER_LOOP1_stage_0_2 OR butterFly2_15_conc_2_itm_0) AND (fsm_output(2)))
      OR ((butterFly2_15_conc_2_itm_0 OR butterFly2_15_conc_2_itm_8_0 OR butterFly2_15_conc_2_itm_7_0)
      AND (fsm_output(4)));
  mult_15_t_and_49_cse <= CONV_SL_1_1(operator_33_true_3_lshift_psp_1_0_sva=STD_LOGIC_VECTOR'("00"))
      AND (fsm_output(9));
  mult_15_t_and_51_cse <= CONV_SL_1_1(operator_33_true_3_lshift_psp_1_0_sva=STD_LOGIC_VECTOR'("01"))
      AND (fsm_output(9));
  mult_15_t_and_53_cse <= CONV_SL_1_1(operator_33_true_3_lshift_psp_1_0_sva=STD_LOGIC_VECTOR'("10"))
      AND (fsm_output(9));
  mult_15_t_and_55_cse <= CONV_SL_1_1(operator_33_true_3_lshift_psp_1_0_sva=STD_LOGIC_VECTOR'("11"))
      AND (fsm_output(9));
  mult_15_t_and_44_cse <= butterFly2_15_tw_equal_tmp_1 AND (fsm_output(7));
  butterFly2_7_tw_nor_cse <= NOT(CONV_SL_1_1(operator_20_false_acc_cse_sva(2 DOWNTO
      1)/=STD_LOGIC_VECTOR'("00")));
  mult_15_t_and_45_cse <= (operator_20_false_acc_cse_sva(0)) AND butterFly2_7_tw_nor_cse
      AND (fsm_output(7));
  butterFly2_7_tw_nor_1_cse <= NOT((operator_20_false_acc_cse_sva(2)) OR (operator_20_false_acc_cse_sva(0)));
  mult_15_t_and_46_cse <= (operator_20_false_acc_cse_sva(1)) AND butterFly2_7_tw_nor_1_cse
      AND (fsm_output(7));
  mult_15_t_and_47_cse <= butterFly2_15_tw_equal_tmp_3_1 AND (fsm_output(7));
  butterFly2_7_tw_nor_2_cse <= NOT(CONV_SL_1_1(operator_20_false_acc_cse_sva(1 DOWNTO
      0)/=STD_LOGIC_VECTOR'("00")));
  mult_15_t_and_48_cse <= (operator_20_false_acc_cse_sva(2)) AND butterFly2_7_tw_nor_2_cse
      AND (fsm_output(7));
  mult_15_t_and_50_cse <= butterFly2_15_tw_equal_tmp_5_1 AND (fsm_output(7));
  mult_15_t_and_52_cse <= butterFly2_15_tw_equal_tmp_6_1 AND (fsm_output(7));
  mult_15_t_and_54_cse <= butterFly2_15_tw_equal_tmp_7_1 AND (fsm_output(7));
  mult_15_t_or_9_cse <= mult_15_t_and_48_cse OR mult_15_t_and_49_cse;
  mult_15_t_or_10_cse <= mult_15_t_and_50_cse OR mult_15_t_and_51_cse;
  mult_15_t_or_11_cse <= mult_15_t_and_52_cse OR mult_15_t_and_53_cse;
  mult_15_t_or_12_cse <= mult_15_t_and_54_cse OR mult_15_t_and_55_cse;
  mult_15_t_and_41_cse <= CONV_SL_1_1(operator_20_false_acc_cse_sva(2 DOWNTO 1)=STD_LOGIC_VECTOR'("01"))
      AND (fsm_output(7));
  mult_15_t_and_42_cse <= CONV_SL_1_1(operator_20_false_acc_cse_sva(2 DOWNTO 1)=STD_LOGIC_VECTOR'("10"))
      AND (fsm_output(7));
  mult_15_t_and_43_cse <= CONV_SL_1_1(operator_20_false_acc_cse_sva(2 DOWNTO 1)=STD_LOGIC_VECTOR'("11"))
      AND (fsm_output(7));
  mult_15_t_and_40_cse <= butterFly2_7_tw_nor_cse AND (fsm_output(7));
  mult_15_t_and_37_cse <= (operator_20_false_acc_cse_sva(0)) AND (NOT (operator_20_false_acc_cse_sva(2)))
      AND (fsm_output(7));
  mult_15_t_and_38_cse <= (operator_20_false_acc_cse_sva(2)) AND (NOT (operator_20_false_acc_cse_sva(0)))
      AND (fsm_output(7));
  mult_15_t_and_39_cse <= (operator_20_false_acc_cse_sva(2)) AND (operator_20_false_acc_cse_sva(0))
      AND (fsm_output(7));
  mult_15_t_and_36_cse <= butterFly2_7_tw_nor_1_cse AND (fsm_output(7));
  mult_15_t_and_30_cse <= CONV_SL_1_1(operator_20_false_acc_cse_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("01"))
      AND (fsm_output(7));
  mult_15_t_and_31_cse <= CONV_SL_1_1(operator_20_false_acc_cse_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("10"))
      AND (fsm_output(7));
  mult_15_t_and_32_cse <= CONV_SL_1_1(operator_20_false_acc_cse_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND (fsm_output(7));
  mult_15_t_and_29_cse <= butterFly2_7_tw_nor_2_cse AND (fsm_output(7));
  mult_15_t_or_3_cse <= modulo_add_1_qelse_or_m1c OR mult_15_t_and_44_cse;
  mult_15_t_or_1_cse <= modulo_add_1_qelse_or_m1c OR mult_15_t_and_36_cse;
  mult_4_t_and_nl <= butterFly1_15_f1_equal_tmp_1 AND (fsm_output(2));
  mult_4_t_and_1_nl <= butterFly1_15_f1_equal_tmp_1_1 AND (fsm_output(2));
  mult_4_t_and_2_nl <= butterFly1_15_f1_equal_tmp_2_1 AND (fsm_output(2));
  mult_4_t_and_3_nl <= butterFly1_15_f1_equal_tmp_3_1 AND (fsm_output(2));
  mult_4_t_and_4_nl <= butterFly1_15_f1_equal_tmp_4_1 AND (fsm_output(2));
  mult_4_t_and_5_nl <= butterFly1_15_f1_equal_tmp_5_1 AND (fsm_output(2));
  mult_4_t_and_6_nl <= butterFly1_15_f1_equal_tmp_6_1 AND (fsm_output(2));
  mult_4_t_and_7_nl <= butterFly1_15_f1_equal_tmp_7_1 AND (fsm_output(2));
  mult_4_t_and_8_nl <= butterFly1_15_f1_equal_tmp_1 AND (fsm_output(4));
  mult_4_t_and_9_nl <= butterFly1_15_f1_equal_tmp_1_1 AND (fsm_output(4));
  mult_4_t_and_10_nl <= butterFly1_15_f1_equal_tmp_2_1 AND (fsm_output(4));
  mult_4_t_and_11_nl <= butterFly1_15_f1_equal_tmp_3_1 AND (fsm_output(4));
  mult_4_t_and_12_nl <= butterFly1_15_f1_equal_tmp_4_1 AND (fsm_output(4));
  mult_4_t_and_13_nl <= butterFly1_15_f1_equal_tmp_5_1 AND (fsm_output(4));
  mult_4_t_and_14_nl <= butterFly1_15_f1_equal_tmp_6_1 AND (fsm_output(4));
  mult_4_t_and_15_nl <= butterFly1_15_f1_equal_tmp_7_1 AND (fsm_output(4));
  mult_4_t_and_16_nl <= butterFly2_15_f1_equal_tmp_1 AND (fsm_output(7));
  mult_4_t_and_17_nl <= butterFly1_15_f1_equal_tmp_3_1 AND (fsm_output(7));
  mult_4_t_and_18_nl <= butterFly1_15_f1_equal_tmp_4_1 AND (fsm_output(7));
  mult_4_t_and_19_nl <= butterFly1_15_f1_equal_tmp_5_1 AND (fsm_output(7));
  mult_4_t_and_20_nl <= butterFly1_15_f1_equal_tmp_6_1 AND (fsm_output(7));
  mult_4_t_and_21_nl <= butterFly1_15_f1_equal_tmp_7_1 AND (fsm_output(7));
  mult_4_t_and_22_nl <= butterFly1_15_f1_equal_tmp_1 AND (fsm_output(7));
  mult_4_t_and_23_nl <= butterFly2_15_f1_equal_tmp_7_1 AND (fsm_output(7));
  mult_4_t_and_24_nl <= butterFly2_15_f1_equal_tmp_1 AND (fsm_output(9));
  mult_4_t_and_25_nl <= butterFly1_15_f1_equal_tmp_3_1 AND (fsm_output(9));
  mult_4_t_and_26_nl <= butterFly1_15_f1_equal_tmp_4_1 AND (fsm_output(9));
  mult_4_t_and_27_nl <= butterFly1_15_f1_equal_tmp_5_1 AND (fsm_output(9));
  mult_4_t_and_28_nl <= butterFly1_15_f1_equal_tmp_6_1 AND (fsm_output(9));
  mult_4_t_and_29_nl <= butterFly1_15_f1_equal_tmp_7_1 AND (fsm_output(9));
  mult_4_t_and_30_nl <= butterFly1_15_f1_equal_tmp_1 AND (fsm_output(9));
  mult_4_t_and_31_nl <= butterFly2_15_f1_equal_tmp_7_1 AND (fsm_output(9));
  mult_4_t_mux1h_1_rmff <= MUX1HOT_v_32_32_2(xt_rsc_0_9_i_qa_d, xt_rsc_1_9_i_qa_d,
      xt_rsc_2_9_i_qa_d, xt_rsc_3_9_i_qa_d, xt_rsc_4_9_i_qa_d, xt_rsc_5_9_i_qa_d,
      xt_rsc_6_9_i_qa_d, xt_rsc_7_9_i_qa_d, yt_rsc_0_9_i_q_d, yt_rsc_1_9_i_q_d, yt_rsc_2_9_i_q_d,
      yt_rsc_3_9_i_q_d, yt_rsc_4_9_i_q_d, yt_rsc_5_9_i_q_d, yt_rsc_6_9_i_q_d, yt_rsc_7_9_i_q_d,
      xt_rsc_0_7_i_qa_d, xt_rsc_1_7_i_qa_d, xt_rsc_2_7_i_qa_d, xt_rsc_3_7_i_qa_d,
      xt_rsc_4_7_i_qa_d, xt_rsc_5_7_i_qa_d, xt_rsc_6_7_i_qa_d, xt_rsc_7_7_i_qa_d,
      yt_rsc_0_23_i_q_d, yt_rsc_1_23_i_q_d, yt_rsc_2_23_i_q_d, yt_rsc_3_23_i_q_d,
      yt_rsc_4_23_i_q_d, yt_rsc_5_23_i_q_d, yt_rsc_6_23_i_q_d, yt_rsc_7_23_i_q_d,
      STD_LOGIC_VECTOR'( mult_4_t_and_nl & mult_4_t_and_1_nl & mult_4_t_and_2_nl
      & mult_4_t_and_3_nl & mult_4_t_and_4_nl & mult_4_t_and_5_nl & mult_4_t_and_6_nl
      & mult_4_t_and_7_nl & mult_4_t_and_8_nl & mult_4_t_and_9_nl & mult_4_t_and_10_nl
      & mult_4_t_and_11_nl & mult_4_t_and_12_nl & mult_4_t_and_13_nl & mult_4_t_and_14_nl
      & mult_4_t_and_15_nl & mult_4_t_and_16_nl & mult_4_t_and_17_nl & mult_4_t_and_18_nl
      & mult_4_t_and_19_nl & mult_4_t_and_20_nl & mult_4_t_and_21_nl & mult_4_t_and_22_nl
      & mult_4_t_and_23_nl & mult_4_t_and_24_nl & mult_4_t_and_25_nl & mult_4_t_and_26_nl
      & mult_4_t_and_27_nl & mult_4_t_and_28_nl & mult_4_t_and_29_nl & mult_4_t_and_30_nl
      & mult_4_t_and_31_nl));
  mult_15_t_or_cse <= modulo_add_1_qelse_or_m1c OR mult_15_t_and_29_cse;
  or_3759_rmff <= ((butterFly1_15_conc_2_itm_7_0 OR butterFly1_15_conc_2_itm_6_0
      OR butterFly1_15_conc_2_itm_5_0) AND or_dcpl_298) OR ((butterFly2_15_conc_2_itm_1_0
      OR butterFly2_15_conc_2_itm_2_0 OR butterFly2_15_conc_2_itm_3_0) AND modulo_add_1_qelse_or_m1c);
  modulo_add_1_qelse_or_m1c <= (fsm_output(2)) OR (fsm_output(4));
  butterFly1_f1_nor_cse <= NOT(CONV_SL_1_1(INNER_LOOP1_r_11_4_sva_6_0(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("00")));
  butterFly2_f1_nor_cse <= NOT(CONV_SL_1_1(INNER_LOOP3_r_11_4_sva_6_0(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("00")));
  butterFly2_16_f1_nor_1_cse <= NOT((INNER_LOOP4_r_11_4_sva_6_0(6)) OR (INNER_LOOP4_r_11_4_sva_6_0(4)));
  INNER_LOOP1_r_INNER_LOOP1_r_and_cse <= MUX_v_7_2_2(STD_LOGIC_VECTOR'("0000000"),
      (z_out_62(6 DOWNTO 0)), (fsm_output(2)));
  modulo_sub_16_qelse_and_ssc <= NOT((z_out_126(31)) OR (fsm_output(9)));
  modulo_sub_16_qelse_and_ssc_1 <= (NOT (z_out_111(31))) AND (fsm_output(9));
  modulo_sub_17_qelse_and_ssc <= NOT((z_out_116(31)) OR (fsm_output(9)));
  modulo_sub_17_qelse_and_ssc_1 <= (NOT (z_out_112(31))) AND (fsm_output(9));
  modulo_sub_18_qelse_and_ssc <= NOT((z_out_123(31)) OR (fsm_output(9)));
  modulo_sub_18_qelse_and_ssc_1 <= (NOT (z_out_113(31))) AND (fsm_output(9));
  modulo_sub_19_qelse_and_ssc <= NOT((z_out_124(31)) OR (fsm_output(9)));
  modulo_sub_19_qelse_and_ssc_1 <= (NOT (z_out_114(31))) AND (fsm_output(9));
  modulo_sub_20_qelse_and_ssc <= NOT((z_out_125(31)) OR (fsm_output(9)));
  modulo_sub_20_qelse_and_ssc_1 <= (NOT (z_out_115(31))) AND (fsm_output(9));
  modulo_sub_21_qelse_and_ssc <= NOT((z_out_111(31)) OR (fsm_output(9)));
  modulo_sub_21_qelse_and_ssc_1 <= (NOT (z_out_116(31))) AND (fsm_output(9));
  modulo_sub_22_qelse_and_ssc <= NOT((z_out_112(31)) OR (fsm_output(9)));
  modulo_sub_22_qelse_and_ssc_1 <= (NOT (z_out_117(31))) AND (fsm_output(9));
  modulo_sub_23_qelse_and_ssc <= NOT((z_out_113(31)) OR (fsm_output(9)));
  modulo_sub_23_qelse_and_ssc_1 <= (NOT (z_out_118(31))) AND (fsm_output(9));
  modulo_sub_24_qelse_and_ssc <= NOT((z_out_114(31)) OR (fsm_output(9)));
  modulo_sub_24_qelse_and_ssc_1 <= (NOT (z_out_119(31))) AND (fsm_output(9));
  modulo_sub_25_qelse_and_ssc <= NOT((z_out_115(31)) OR (fsm_output(9)));
  modulo_sub_25_qelse_and_ssc_1 <= (NOT (z_out_120(31))) AND (fsm_output(9));
  modulo_sub_26_qelse_and_ssc <= NOT((z_out_117(31)) OR (fsm_output(9)));
  modulo_sub_26_qelse_and_ssc_1 <= (NOT (z_out_121(31))) AND (fsm_output(9));
  modulo_sub_27_qelse_and_ssc <= NOT((z_out_118(31)) OR (fsm_output(9)));
  modulo_sub_27_qelse_and_ssc_1 <= (NOT (z_out_122(31))) AND (fsm_output(9));
  modulo_sub_28_qelse_and_ssc <= NOT((z_out_119(31)) OR (fsm_output(9)));
  modulo_sub_28_qelse_and_ssc_1 <= (NOT (z_out_123(31))) AND (fsm_output(9));
  modulo_sub_29_qelse_and_ssc <= NOT((z_out_120(31)) OR (fsm_output(9)));
  modulo_sub_29_qelse_and_ssc_1 <= (NOT (z_out_124(31))) AND (fsm_output(9));
  modulo_sub_30_qelse_and_ssc <= NOT((z_out_121(31)) OR (fsm_output(9)));
  modulo_sub_30_qelse_and_ssc_1 <= (NOT (z_out_125(31))) AND (fsm_output(9));
  modulo_sub_31_qelse_and_ssc <= NOT((z_out_122(31)) OR (fsm_output(9)));
  modulo_sub_31_qelse_and_ssc_1 <= (NOT (z_out_126(31))) AND (fsm_output(9));
  butterFly2_16_f1_butterFly2_16_f1_and_6_cse <= CONV_SL_1_1(INNER_LOOP4_r_11_4_sva_6_0(6
      DOWNTO 4)=STD_LOGIC_VECTOR'("111"));
  INNER_LOOP1_r_INNER_LOOP1_r_and_3_cse <= MUX_v_7_2_2(STD_LOGIC_VECTOR'("0000000"),
      (z_out_62(6 DOWNTO 0)), (fsm_output(7)));
  INNER_LOOP1_r_INNER_LOOP1_r_and_5_cse <= MUX_v_7_2_2(STD_LOGIC_VECTOR'("0000000"),
      (z_out_62(6 DOWNTO 0)), (fsm_output(9)));
  or_383_cse <= (butterFly1_15_conc_2_itm_9_2_1(0)) OR butterFly1_15_conc_2_itm_9_0;
  or_398_cse <= (NOT (butterFly1_15_conc_2_itm_9_2_1(0))) OR butterFly1_15_conc_2_itm_9_0;
  and_8913_cse <= (butterFly1_15_conc_2_itm_9_2_1(0)) AND butterFly1_15_conc_2_itm_9_0
      AND (butterFly1_15_conc_2_itm_9_2_1(1)) AND INNER_LOOP1_stage_0_10;
  nor_27_cse <= NOT((butterFly1_15_conc_2_itm_9_2_1(0)) OR (NOT butterFly1_15_conc_2_itm_9_0));
  and_8912_cse <= (butterFly1_15_conc_2_itm_9_2_1(0)) AND butterFly1_15_conc_2_itm_9_0;
  mult_t_mul_cmp_5_a_mx0w1 <= MUX1HOT_v_32_8_2(yt_rsc_0_23_i_q_d, yt_rsc_1_23_i_q_d,
      yt_rsc_2_23_i_q_d, yt_rsc_3_23_i_q_d, yt_rsc_4_23_i_q_d, yt_rsc_5_23_i_q_d,
      yt_rsc_6_23_i_q_d, yt_rsc_7_23_i_q_d, STD_LOGIC_VECTOR'( butterFly1_15_f1_equal_tmp_1
      & butterFly1_15_f1_equal_tmp_1_1 & butterFly1_15_f1_equal_tmp_2_1 & butterFly1_15_f1_equal_tmp_3_1
      & butterFly1_15_f1_equal_tmp_4_1 & butterFly1_15_f1_equal_tmp_5_1 & butterFly1_15_f1_equal_tmp_6_1
      & butterFly1_15_f1_equal_tmp_7_1));
  mult_t_mul_cmp_5_a_mx0w4 <= MUX1HOT_v_32_8_2(yt_rsc_0_9_i_q_d, yt_rsc_1_9_i_q_d,
      yt_rsc_2_9_i_q_d, yt_rsc_3_9_i_q_d, yt_rsc_4_9_i_q_d, yt_rsc_5_9_i_q_d, yt_rsc_6_9_i_q_d,
      yt_rsc_7_9_i_q_d, STD_LOGIC_VECTOR'( butterFly2_15_f1_equal_tmp_1 & butterFly1_15_f1_equal_tmp_3_1
      & butterFly1_15_f1_equal_tmp_4_1 & butterFly1_15_f1_equal_tmp_5_1 & butterFly1_15_f1_equal_tmp_6_1
      & butterFly1_15_f1_equal_tmp_7_1 & butterFly1_15_f1_equal_tmp_1 & butterFly2_15_f1_equal_tmp_7_1));
  mult_t_mul_cmp_11_a_mx0w3 <= MUX1HOT_v_32_8_2(xt_rsc_0_9_i_qa_d, xt_rsc_1_9_i_qa_d,
      xt_rsc_2_9_i_qa_d, xt_rsc_3_9_i_qa_d, xt_rsc_4_9_i_qa_d, xt_rsc_5_9_i_qa_d,
      xt_rsc_6_9_i_qa_d, xt_rsc_7_9_i_qa_d, STD_LOGIC_VECTOR'( butterFly2_15_f1_equal_tmp_1
      & butterFly1_15_f1_equal_tmp_3_1 & butterFly1_15_f1_equal_tmp_4_1 & butterFly1_15_f1_equal_tmp_5_1
      & butterFly1_15_f1_equal_tmp_6_1 & butterFly1_15_f1_equal_tmp_7_1 & butterFly1_15_f1_equal_tmp_1
      & butterFly2_15_f1_equal_tmp_7_1));
  mult_15_if_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_15_res_sva_1)
      - UNSIGNED(p_sva), 32));
  mult_31_acc_1_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & mult_15_res_sva_1)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(NOT p_sva), 32), 33) + UNSIGNED'( "000000000000000000000000000000001"),
      33));
  mult_15_res_lpi_3_dfm_1_mx0 <= MUX_v_32_2_2(STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_15_if_acc_nl),
      32)), mult_15_res_sva_1, mult_31_acc_1_nl(32));
  mult_14_if_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_14_res_sva_1)
      - UNSIGNED(p_sva), 32));
  mult_30_acc_1_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & mult_14_res_sva_1)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(NOT p_sva), 32), 33) + UNSIGNED'( "000000000000000000000000000000001"),
      33));
  mult_14_res_lpi_3_dfm_1_mx0 <= MUX_v_32_2_2(STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_14_if_acc_nl),
      32)), mult_14_res_sva_1, mult_30_acc_1_nl(32));
  mult_13_if_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_13_res_sva_1)
      - UNSIGNED(p_sva), 32));
  mult_29_acc_1_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & mult_13_res_sva_1)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(NOT p_sva), 32), 33) + UNSIGNED'( "000000000000000000000000000000001"),
      33));
  mult_13_res_lpi_3_dfm_1_mx0 <= MUX_v_32_2_2(STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_13_if_acc_nl),
      32)), mult_13_res_sva_1, mult_29_acc_1_nl(32));
  mult_12_if_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_12_res_sva_1)
      - UNSIGNED(p_sva), 32));
  mult_28_acc_1_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & mult_12_res_sva_1)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(NOT p_sva), 32), 33) + UNSIGNED'( "000000000000000000000000000000001"),
      33));
  mult_12_res_lpi_3_dfm_1_mx0 <= MUX_v_32_2_2(STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_12_if_acc_nl),
      32)), mult_12_res_sva_1, mult_28_acc_1_nl(32));
  mult_11_if_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_11_res_sva_1)
      - UNSIGNED(p_sva), 32));
  mult_27_acc_1_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & mult_11_res_sva_1)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(NOT p_sva), 32), 33) + UNSIGNED'( "000000000000000000000000000000001"),
      33));
  mult_11_res_lpi_3_dfm_1_mx0 <= MUX_v_32_2_2(STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_11_if_acc_nl),
      32)), mult_11_res_sva_1, mult_27_acc_1_nl(32));
  mult_10_if_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_10_res_sva_1)
      - UNSIGNED(p_sva), 32));
  mult_26_acc_1_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & mult_10_res_sva_1)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(NOT p_sva), 32), 33) + UNSIGNED'( "000000000000000000000000000000001"),
      33));
  mult_10_res_lpi_3_dfm_1_mx0 <= MUX_v_32_2_2(STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_10_if_acc_nl),
      32)), mult_10_res_sva_1, mult_26_acc_1_nl(32));
  mult_9_if_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_9_res_sva_1) -
      UNSIGNED(p_sva), 32));
  mult_25_acc_1_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & mult_9_res_sva_1)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(NOT p_sva), 32), 33) + UNSIGNED'( "000000000000000000000000000000001"),
      33));
  mult_9_res_lpi_3_dfm_1_mx0 <= MUX_v_32_2_2(STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_9_if_acc_nl),
      32)), mult_9_res_sva_1, mult_25_acc_1_nl(32));
  mult_8_if_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_8_res_sva_1) -
      UNSIGNED(p_sva), 32));
  mult_24_acc_1_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & mult_8_res_sva_1)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(NOT p_sva), 32), 33) + UNSIGNED'( "000000000000000000000000000000001"),
      33));
  mult_8_res_lpi_3_dfm_1_mx0 <= MUX_v_32_2_2(STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_8_if_acc_nl),
      32)), mult_8_res_sva_1, mult_24_acc_1_nl(32));
  mult_7_if_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_7_res_sva_1) -
      UNSIGNED(p_sva), 32));
  mult_23_acc_1_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & mult_7_res_sva_1)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(NOT p_sva), 32), 33) + UNSIGNED'( "000000000000000000000000000000001"),
      33));
  mult_7_res_lpi_3_dfm_1_mx0 <= MUX_v_32_2_2(STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_7_if_acc_nl),
      32)), mult_7_res_sva_1, mult_23_acc_1_nl(32));
  mult_6_if_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_6_res_sva_1) -
      UNSIGNED(p_sva), 32));
  mult_22_acc_1_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & mult_6_res_sva_1)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(NOT p_sva), 32), 33) + UNSIGNED'( "000000000000000000000000000000001"),
      33));
  mult_6_res_lpi_3_dfm_1_mx0 <= MUX_v_32_2_2(STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_6_if_acc_nl),
      32)), mult_6_res_sva_1, mult_22_acc_1_nl(32));
  mult_5_if_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_5_res_sva_1) -
      UNSIGNED(p_sva), 32));
  mult_21_acc_1_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & mult_5_res_sva_1)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(NOT p_sva), 32), 33) + UNSIGNED'( "000000000000000000000000000000001"),
      33));
  mult_5_res_lpi_3_dfm_1_mx0 <= MUX_v_32_2_2(STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_5_if_acc_nl),
      32)), mult_5_res_sva_1, mult_21_acc_1_nl(32));
  mult_4_if_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_4_res_sva_1) -
      UNSIGNED(p_sva), 32));
  mult_20_acc_1_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & mult_4_res_sva_1)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(NOT p_sva), 32), 33) + UNSIGNED'( "000000000000000000000000000000001"),
      33));
  mult_4_res_lpi_3_dfm_1_mx0 <= MUX_v_32_2_2(STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_4_if_acc_nl),
      32)), mult_4_res_sva_1, mult_20_acc_1_nl(32));
  mult_3_if_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_3_res_sva_1) -
      UNSIGNED(p_sva), 32));
  mult_19_acc_1_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & mult_3_res_sva_1)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(NOT p_sva), 32), 33) + UNSIGNED'( "000000000000000000000000000000001"),
      33));
  mult_3_res_lpi_3_dfm_1_mx0 <= MUX_v_32_2_2(STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_3_if_acc_nl),
      32)), mult_3_res_sva_1, mult_19_acc_1_nl(32));
  mult_2_if_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_2_res_sva_1) -
      UNSIGNED(p_sva), 32));
  mult_18_acc_1_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & mult_2_res_sva_1)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(NOT p_sva), 32), 33) + UNSIGNED'( "000000000000000000000000000000001"),
      33));
  mult_2_res_lpi_3_dfm_1_mx0 <= MUX_v_32_2_2(STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_2_if_acc_nl),
      32)), mult_2_res_sva_1, mult_18_acc_1_nl(32));
  mult_1_if_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_1_res_sva_1) -
      UNSIGNED(p_sva), 32));
  mult_17_acc_1_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & mult_1_res_sva_1)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(NOT p_sva), 32), 33) + UNSIGNED'( "000000000000000000000000000000001"),
      33));
  mult_1_res_lpi_3_dfm_1_mx0 <= MUX_v_32_2_2(STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_1_if_acc_nl),
      32)), mult_1_res_sva_1, mult_17_acc_1_nl(32));
  mult_if_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_res_sva_1) - UNSIGNED(p_sva),
      32));
  mult_16_acc_1_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & mult_res_sva_1)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(NOT p_sva), 32), 33) + UNSIGNED'( "000000000000000000000000000000001"),
      33));
  mult_res_lpi_3_dfm_1_mx0 <= MUX_v_32_2_2(STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_if_acc_nl),
      32)), mult_res_sva_1, mult_16_acc_1_nl(32));
  INNER_LOOP2_r_11_4_sva_6_0_mx1 <= MUX_v_7_2_2(STD_LOGIC_VECTOR'("0000000"), (z_out_62(6
      DOWNTO 0)), (fsm_output(4)));
  mult_15_res_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_15_z_asn_itm_3)
      - UNSIGNED(mult_z_mul_cmp_1_z), 32));
  mult_14_res_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_14_z_asn_itm_3)
      - UNSIGNED(mult_z_mul_cmp_3_z), 32));
  mult_13_res_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_13_z_asn_itm_3)
      - UNSIGNED(mult_z_mul_cmp_5_z), 32));
  mult_12_res_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_12_z_asn_itm_3)
      - UNSIGNED(mult_z_mul_cmp_7_z), 32));
  mult_11_res_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_11_z_asn_itm_3)
      - UNSIGNED(mult_z_mul_cmp_9_z), 32));
  mult_10_res_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_10_z_asn_itm_3)
      - UNSIGNED(mult_z_mul_cmp_11_z), 32));
  mult_9_res_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_25_z_asn_itm_3)
      - UNSIGNED(mult_z_mul_cmp_13_z), 32));
  mult_8_res_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_24_z_asn_itm_3)
      - UNSIGNED(mult_z_mul_cmp_15_z), 32));
  mult_7_res_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_23_z_asn_itm_3)
      - UNSIGNED(mult_z_mul_cmp_17_z), 32));
  mult_6_res_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_22_z_asn_itm_3)
      - UNSIGNED(mult_z_mul_cmp_19_z), 32));
  mult_5_res_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_21_z_asn_itm_3)
      - UNSIGNED(mult_z_mul_cmp_21_z), 32));
  mult_4_res_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_20_z_asn_itm_3)
      - UNSIGNED(mult_z_mul_cmp_23_z), 32));
  mult_3_res_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_19_z_asn_itm_3)
      - UNSIGNED(mult_z_mul_cmp_25_z), 32));
  mult_2_res_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_18_z_asn_itm_3)
      - UNSIGNED(mult_z_mul_cmp_27_z), 32));
  mult_1_res_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_17_z_asn_itm_3)
      - UNSIGNED(mult_z_mul_cmp_29_z), 32));
  mult_res_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_16_z_asn_itm_3)
      - UNSIGNED(mult_z_mul_cmp_31_z), 32));
  tmp_71_lpi_3_dfm_1 <= MUX1HOT_v_32_8_2(xt_rsc_0_7_i_qa_d, xt_rsc_1_7_i_qa_d, xt_rsc_2_7_i_qa_d,
      xt_rsc_3_7_i_qa_d, xt_rsc_4_7_i_qa_d, xt_rsc_5_7_i_qa_d, xt_rsc_6_7_i_qa_d,
      xt_rsc_7_7_i_qa_d, STD_LOGIC_VECTOR'( butterFly1_15_f1_equal_tmp_1 & butterFly1_15_f1_equal_tmp_1_1
      & butterFly1_15_f1_equal_tmp_2_1 & butterFly1_15_f1_equal_tmp_3_1 & butterFly1_15_f1_equal_tmp_4_1
      & butterFly1_15_f1_equal_tmp_5_1 & butterFly1_15_f1_equal_tmp_6_1 & butterFly1_15_f1_equal_tmp_7_1));
  operator_33_true_2_lshift_psp_2_0_sva_mx0 <= MUX_v_3_2_2((z_out_60(2 DOWNTO 0)),
      operator_20_false_acc_cse_sva, fsm_output(7));
  INNER_LOOP4_nor_tmp <= NOT(INNER_LOOP1_stage_0 OR butterFly1_15_conc_2_itm_2_0
      OR butterFly1_15_conc_2_itm_3_0 OR butterFly1_15_conc_2_itm_4_0 OR butterFly1_15_conc_2_itm_5_0
      OR butterFly1_15_conc_2_itm_6_0 OR butterFly1_15_conc_2_itm_7_0 OR butterFly1_15_conc_2_itm_8_0
      OR butterFly1_15_conc_2_itm_9_0 OR butterFly1_15_conc_2_itm_0);
  or_dcpl <= butterFly1_15_conc_2_itm_5_0 OR butterFly2_15_conc_2_itm_1_0;
  or_dcpl_2 <= butterFly1_15_conc_2_itm_4_0 OR butterFly2_15_conc_2_itm_0;
  or_dcpl_8 <= butterFly1_15_conc_2_itm_8_0 OR butterFly2_15_conc_2_itm_4_0;
  or_dcpl_10 <= butterFly1_15_conc_2_itm_7_0 OR butterFly2_15_conc_2_itm_3_0;
  or_dcpl_12 <= butterFly1_15_conc_2_itm_6_0 OR butterFly2_15_conc_2_itm_2_0;
  or_dcpl_19 <= butterFly2_15_conc_2_itm_4_0 OR butterFly2_15_conc_2_itm_0;
  or_dcpl_22 <= butterFly2_15_conc_2_itm_4_0 OR butterFly2_15_conc_2_itm_8_0;
  or_dcpl_25 <= butterFly2_15_conc_2_itm_4_0 OR butterFly2_15_conc_2_itm_7_0;
  or_dcpl_30 <= butterFly2_15_conc_2_itm_4_0 OR butterFly2_15_conc_2_itm_3_0;
  or_dcpl_33 <= butterFly2_15_conc_2_itm_4_0 OR butterFly2_15_conc_2_itm_2_0;
  or_dcpl_36 <= butterFly2_15_conc_2_itm_4_0 OR butterFly2_15_conc_2_itm_1_0;
  or_dcpl_63 <= butterFly1_15_conc_2_itm_7_0 OR butterFly1_15_conc_2_itm_8_0;
  or_dcpl_70 <= butterFly1_15_conc_2_itm_8_0 OR butterFly1_15_conc_2_itm_9_0;
  or_dcpl_72 <= butterFly2_15_conc_2_itm_3_0 OR butterFly2_15_conc_2_itm_5_0;
  or_dcpl_76 <= butterFly1_15_conc_2_itm_2_0 OR butterFly1_15_conc_2_itm_8_0;
  or_dcpl_78 <= butterFly2_15_conc_2_itm_3_0 OR butterFly2_15_conc_2_itm_7_0;
  or_dcpl_80 <= butterFly1_15_conc_2_itm_3_0 OR butterFly1_15_conc_2_itm_8_0;
  or_dcpl_82 <= butterFly2_15_conc_2_itm_3_0 OR butterFly2_15_conc_2_itm_8_0;
  or_dcpl_88 <= butterFly2_15_conc_2_itm_2_0 OR butterFly2_15_conc_2_itm_8_0;
  or_dcpl_89 <= butterFly1_15_conc_2_itm_7_0 OR butterFly1_15_conc_2_itm_3_0;
  or_dcpl_94 <= butterFly1_15_conc_2_itm_7_0 OR butterFly2_15_conc_2_itm_2_0;
  or_dcpl_105 <= butterFly1_15_conc_2_itm_7_0 OR butterFly1_15_conc_2_itm_9_0;
  or_dcpl_107 <= butterFly2_15_conc_2_itm_2_0 OR butterFly2_15_conc_2_itm_5_0;
  or_dcpl_109 <= butterFly1_15_conc_2_itm_2_0 OR butterFly1_15_conc_2_itm_7_0;
  or_dcpl_111 <= butterFly2_15_conc_2_itm_2_0 OR butterFly2_15_conc_2_itm_7_0;
  or_dcpl_116 <= butterFly2_15_conc_2_itm_1_0 OR butterFly2_15_conc_2_itm_7_0;
  or_dcpl_117 <= butterFly1_15_conc_2_itm_2_0 OR butterFly1_15_conc_2_itm_6_0;
  or_dcpl_119 <= butterFly1_15_conc_2_itm_6_0 OR butterFly1_15_conc_2_itm_3_0;
  or_dcpl_121 <= butterFly2_15_conc_2_itm_1_0 OR butterFly2_15_conc_2_itm_8_0;
  or_dcpl_125 <= butterFly1_15_conc_2_itm_6_0 OR butterFly2_15_conc_2_itm_1_0;
  or_dcpl_133 <= butterFly1_15_conc_2_itm_7_0 OR butterFly1_15_conc_2_itm_6_0;
  or_dcpl_135 <= butterFly2_15_conc_2_itm_1_0 OR butterFly2_15_conc_2_itm_3_0;
  or_dcpl_139 <= butterFly1_15_conc_2_itm_6_0 OR butterFly1_15_conc_2_itm_9_0;
  or_dcpl_141 <= butterFly2_15_conc_2_itm_1_0 OR butterFly2_15_conc_2_itm_5_0;
  or_dcpl_146 <= butterFly1_15_conc_2_itm_2_0 OR butterFly1_15_conc_2_itm_5_0;
  or_dcpl_148 <= butterFly2_15_conc_2_itm_0 OR butterFly2_15_conc_2_itm_7_0;
  or_dcpl_150 <= butterFly1_15_conc_2_itm_5_0 OR butterFly1_15_conc_2_itm_3_0;
  or_dcpl_152 <= butterFly2_15_conc_2_itm_0 OR butterFly2_15_conc_2_itm_8_0;
  or_dcpl_161 <= butterFly1_15_conc_2_itm_6_0 OR butterFly1_15_conc_2_itm_5_0;
  or_dcpl_163 <= butterFly2_15_conc_2_itm_0 OR butterFly2_15_conc_2_itm_2_0;
  or_dcpl_165 <= butterFly1_15_conc_2_itm_7_0 OR butterFly1_15_conc_2_itm_5_0;
  or_dcpl_167 <= butterFly2_15_conc_2_itm_0 OR butterFly2_15_conc_2_itm_3_0;
  or_dcpl_171 <= butterFly1_15_conc_2_itm_5_0 OR butterFly1_15_conc_2_itm_9_0;
  or_dcpl_173 <= butterFly2_15_conc_2_itm_0 OR butterFly2_15_conc_2_itm_5_0;
  or_dcpl_180 <= INNER_LOOP1_stage_0_3 OR butterFly2_15_conc_2_itm_5_0;
  or_dcpl_181 <= butterFly1_15_conc_2_itm_4_0 OR butterFly1_15_conc_2_itm_9_0;
  or_dcpl_185 <= butterFly1_15_conc_2_itm_2_0 OR butterFly1_15_conc_2_itm_4_0;
  or_dcpl_187 <= INNER_LOOP1_stage_0_3 OR butterFly2_15_conc_2_itm_7_0;
  or_dcpl_189 <= butterFly1_15_conc_2_itm_4_0 OR butterFly1_15_conc_2_itm_3_0;
  or_dcpl_197 <= butterFly1_15_conc_2_itm_5_0 OR butterFly1_15_conc_2_itm_4_0;
  or_dcpl_199 <= INNER_LOOP1_stage_0_3 OR butterFly2_15_conc_2_itm_1_0;
  or_dcpl_201 <= butterFly1_15_conc_2_itm_6_0 OR butterFly1_15_conc_2_itm_4_0;
  or_dcpl_203 <= INNER_LOOP1_stage_0_3 OR butterFly2_15_conc_2_itm_2_0;
  or_dcpl_205 <= butterFly1_15_conc_2_itm_7_0 OR butterFly1_15_conc_2_itm_4_0;
  or_dcpl_207 <= INNER_LOOP1_stage_0_3 OR butterFly2_15_conc_2_itm_3_0;
  or_dcpl_210 <= INNER_LOOP1_stage_0_3 OR butterFly2_15_conc_2_itm_4_0;
  or_dcpl_215 <= INNER_LOOP1_stage_0_2 OR butterFly2_15_conc_2_itm_4_0;
  or_dcpl_218 <= butterFly1_15_conc_2_itm_3_0 OR butterFly1_15_conc_2_itm_9_0;
  or_dcpl_220 <= INNER_LOOP1_stage_0_2 OR butterFly2_15_conc_2_itm_5_0;
  or_dcpl_224 <= butterFly1_15_conc_2_itm_2_0 OR butterFly1_15_conc_2_itm_3_0;
  or_dcpl_234 <= INNER_LOOP1_stage_0_2 OR butterFly2_15_conc_2_itm_0;
  or_dcpl_238 <= INNER_LOOP1_stage_0_2 OR butterFly2_15_conc_2_itm_1_0;
  or_dcpl_242 <= INNER_LOOP1_stage_0_2 OR butterFly2_15_conc_2_itm_2_0;
  or_dcpl_246 <= INNER_LOOP1_stage_0_2 OR butterFly2_15_conc_2_itm_3_0;
  or_dcpl_274 <= butterFly1_15_conc_2_itm_9_0 OR butterFly2_15_conc_2_itm_5_0;
  and_dcpl_62 <= INNER_LOOP4_nor_tmp AND c_1_sva;
  or_tmp_26 <= butterFly1_15_f1_equal_tmp_2_1 OR (butterFly2_15_conc_itm_10_2_1(1))
      OR (NOT butterFly1_15_conc_2_itm_1_0);
  or_tmp_29 <= (butterFly2_15_conc_2_itm_9_2_1(1)) OR butterFly1_15_f1_equal_tmp_1_1
      OR (NOT butterFly1_15_conc_2_itm_0);
  nor_62_nl <= NOT(butterFly1_15_conc_2_itm_1_0 OR (NOT or_tmp_29));
  or_325_nl <= butterFly1_15_f1_equal_tmp_2_1 OR (butterFly2_15_conc_itm_10_2_1(1));
  mux_tmp <= MUX_s_1_2_2(nor_62_nl, or_tmp_29, or_325_nl);
  or_tmp_35 <= (butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1(1)) OR (NOT butterFly1_15_conc_2_itm_2_0);
  not_tmp_25 <= NOT((NOT((butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1(1)) OR
      (NOT butterFly1_15_conc_2_itm_2_0))) OR INNER_LOOP1_stage_0);
  or_tmp_38 <= (butterFly1_15_conc_2_itm_9_2_1(0)) OR butterFly1_15_conc_2_itm_9_0
      OR (butterFly1_15_conc_2_itm_9_2_1(1)) OR (NOT INNER_LOOP1_stage_0_10);
  or_tmp_40 <= (butterFly2_15_conc_2_itm_6_2_1(1)) OR (NOT INNER_LOOP1_stage_0_11)
      OR INNER_LOOP2_stage_0_10;
  not_tmp_29 <= NOT(INNER_LOOP1_stage_0_10 OR (NOT or_tmp_40));
  and_dcpl_66 <= NOT(CONV_SL_1_1(butterFly2_15_conc_2_itm_9_2_1/=STD_LOGIC_VECTOR'("00")));
  and_dcpl_67 <= butterFly1_15_conc_2_itm_0 AND (NOT butterFly1_15_f1_equal_tmp_1_1);
  and_dcpl_68 <= and_dcpl_67 AND and_dcpl_66;
  and_dcpl_69 <= NOT(butterFly1_15_conc_2_itm_9_0 OR (butterFly1_15_conc_2_itm_9_2_1(0)));
  and_dcpl_70 <= INNER_LOOP1_stage_0_10 AND (NOT (butterFly1_15_conc_2_itm_9_2_1(1)));
  and_dcpl_73 <= INNER_LOOP1_stage_0 AND (NOT (INNER_LOOP4_r_11_4_sva_6_0(5)));
  and_dcpl_76 <= INNER_LOOP1_stage_0 AND (NOT (INNER_LOOP2_r_11_4_sva_6_0(5)));
  nor_tmp_1 <= butterFly1_15_f1_equal_tmp_1_1 AND butterFly1_15_conc_2_itm_0;
  or_tmp_48 <= (NOT butterFly1_15_f1_equal_tmp_2_1) OR (butterFly2_15_conc_itm_10_2_1(1))
      OR (NOT butterFly1_15_conc_2_itm_1_0);
  or_tmp_50 <= (butterFly2_15_conc_2_itm_9_2_1(1)) OR (NOT nor_tmp_1);
  nor_56_nl <= NOT(butterFly1_15_conc_2_itm_1_0 OR (NOT or_tmp_50));
  or_347_nl <= (NOT butterFly1_15_f1_equal_tmp_2_1) OR (butterFly2_15_conc_itm_10_2_1(1));
  mux_tmp_7 <= MUX_s_1_2_2(nor_56_nl, or_tmp_50, or_347_nl);
  or_tmp_53 <= (butterFly1_15_conc_2_itm_9_2_1(0)) OR (NOT butterFly1_15_conc_2_itm_9_0)
      OR (butterFly1_15_conc_2_itm_9_2_1(1)) OR (NOT INNER_LOOP1_stage_0_10);
  or_tmp_55 <= (butterFly2_15_conc_2_itm_6_2_1(1)) OR (NOT(INNER_LOOP1_stage_0_11
      AND INNER_LOOP2_stage_0_10));
  not_tmp_50 <= NOT(INNER_LOOP1_stage_0_10 OR (NOT or_tmp_55));
  and_dcpl_78 <= nor_tmp_1 AND and_dcpl_66;
  and_dcpl_79 <= butterFly1_15_conc_2_itm_9_0 AND (NOT (butterFly1_15_conc_2_itm_9_2_1(0)));
  or_tmp_64 <= (NOT (butterFly1_15_conc_2_itm_9_2_1(0))) OR butterFly1_15_conc_2_itm_9_0
      OR (butterFly1_15_conc_2_itm_9_2_1(1)) OR (NOT INNER_LOOP1_stage_0_10);
  and_dcpl_81 <= CONV_SL_1_1(butterFly2_15_conc_2_itm_9_2_1=STD_LOGIC_VECTOR'("01"));
  and_dcpl_82 <= and_dcpl_67 AND and_dcpl_81;
  and_dcpl_83 <= (NOT butterFly1_15_conc_2_itm_9_0) AND (butterFly1_15_conc_2_itm_9_2_1(0));
  or_tmp_72 <= NOT((butterFly1_15_conc_2_itm_9_2_1(0)) AND butterFly1_15_conc_2_itm_9_0
      AND (NOT (butterFly1_15_conc_2_itm_9_2_1(1))) AND INNER_LOOP1_stage_0_10);
  and_dcpl_89 <= nor_tmp_1 AND and_dcpl_81;
  nand_7_cse <= NOT((butterFly2_15_conc_itm_10_2_1(1)) AND butterFly1_15_conc_2_itm_1_0);
  or_tmp_75 <= butterFly1_15_f1_equal_tmp_2_1 OR nand_7_cse;
  or_tmp_77 <= (NOT (butterFly2_15_conc_2_itm_9_2_1(1))) OR butterFly1_15_f1_equal_tmp_1_1
      OR (NOT butterFly1_15_conc_2_itm_0);
  and_8934_nl <= nand_7_cse AND or_tmp_77;
  mux_tmp_22 <= MUX_s_1_2_2(and_8934_nl, or_tmp_77, butterFly1_15_f1_equal_tmp_2_1);
  nor_tmp_6 <= (INNER_LOOP4_r_11_4_sva_6_0(5)) AND INNER_LOOP1_stage_0;
  and_8932_cse <= (butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1(1)) AND butterFly1_15_conc_2_itm_2_0;
  or_tmp_82 <= and_8932_cse OR INNER_LOOP1_stage_0;
  nor_tmp_10 <= (butterFly1_15_conc_2_itm_9_2_1(1)) AND INNER_LOOP1_stage_0_10;
  or_tmp_84 <= (butterFly1_15_conc_2_itm_9_2_1(0)) OR butterFly1_15_conc_2_itm_9_0
      OR (NOT nor_tmp_10);
  or_tmp_86 <= (NOT (butterFly2_15_conc_2_itm_6_2_1(1))) OR (NOT INNER_LOOP1_stage_0_11)
      OR INNER_LOOP2_stage_0_10;
  not_tmp_67 <= (NOT((butterFly1_15_conc_2_itm_9_2_1(1)) AND INNER_LOOP1_stage_0_10))
      AND or_tmp_86;
  not_tmp_69 <= NOT((INNER_LOOP2_r_11_4_sva_6_0(5)) AND INNER_LOOP1_stage_0);
  or_tmp_90 <= (INNER_LOOP2_r_11_4_sva_6_0(4)) OR (INNER_LOOP2_r_11_4_sva_6_0(6))
      OR not_tmp_69;
  and_dcpl_92 <= CONV_SL_1_1(butterFly2_15_conc_2_itm_9_2_1=STD_LOGIC_VECTOR'("10"));
  and_dcpl_93 <= and_dcpl_67 AND and_dcpl_92;
  nor_tmp_14 <= (butterFly2_15_conc_2_itm_9_2_1(1)) AND butterFly1_15_f1_equal_tmp_1_1
      AND butterFly1_15_conc_2_itm_0;
  nor_tmp_15 <= butterFly1_15_f1_equal_tmp_2_1 AND (butterFly2_15_conc_itm_10_2_1(1))
      AND butterFly1_15_conc_2_itm_1_0;
  or_tmp_93 <= nor_tmp_15 OR nor_tmp_14;
  or_tmp_94 <= (butterFly1_15_conc_2_itm_9_2_1(0)) OR (NOT(butterFly1_15_conc_2_itm_9_0
      AND (butterFly1_15_conc_2_itm_9_2_1(1)) AND INNER_LOOP1_stage_0_10));
  nor_tmp_19 <= (butterFly2_15_conc_2_itm_6_2_1(1)) AND INNER_LOOP1_stage_0_11 AND
      INNER_LOOP2_stage_0_10;
  and_dcpl_96 <= nor_tmp_1 AND and_dcpl_92;
  or_tmp_99 <= (NOT (INNER_LOOP4_r_11_4_sva_6_0(4))) OR (INNER_LOOP4_r_11_4_sva_6_0(6))
      OR (NOT nor_tmp_6);
  or_tmp_102 <= (NOT (butterFly1_15_conc_2_itm_9_2_1(0))) OR butterFly1_15_conc_2_itm_9_0
      OR (NOT nor_tmp_10);
  or_tmp_104 <= (NOT (INNER_LOOP2_r_11_4_sva_6_0(4))) OR (INNER_LOOP2_r_11_4_sva_6_0(6))
      OR not_tmp_69;
  and_dcpl_99 <= and_dcpl_67 AND CONV_SL_1_1(butterFly2_15_conc_2_itm_9_2_1=STD_LOGIC_VECTOR'("11"));
  nor_tmp_22 <= CONV_SL_1_1(butterFly2_15_conc_2_itm_9_2_1=STD_LOGIC_VECTOR'("11"))
      AND butterFly1_15_f1_equal_tmp_1_1 AND butterFly1_15_conc_2_itm_0;
  or_tmp_112 <= butterFly1_15_f1_equal_tmp_1_1 OR (NOT butterFly1_15_conc_2_itm_0);
  not_tmp_87 <= NOT(butterFly1_15_conc_2_itm_9_0 OR and_dcpl_67);
  or_409_nl <= (butterFly2_15_conc_2_itm_8_2_1(1)) OR butterFly2_15_conc_2_itm_8_0;
  mux_44_nl <= MUX_s_1_2_2(not_tmp_87, or_tmp_112, or_409_nl);
  or_408_nl <= (butterFly2_15_conc_2_itm_8_2_1(1)) OR butterFly2_15_conc_2_itm_8_0
      OR (NOT butterFly1_15_conc_2_itm_9_0);
  mux_tmp_45 <= MUX_s_1_2_2(mux_44_nl, or_408_nl, butterFly2_15_conc_2_itm_9_2_1(1));
  or_tmp_120 <= butterFly1_15_conc_2_itm_8_0 OR (butterFly1_15_conc_2_itm_8_2_1(1))
      OR (NOT butterFly2_15_conc_2_itm_5_0);
  or_tmp_122 <= (butterFly1_15_conc_2_itm_9_2_1(1)) OR (NOT INNER_LOOP1_stage_0_10);
  not_tmp_91 <= NOT(butterFly2_15_conc_2_itm_5_0 OR and_dcpl_70);
  or_419_nl <= butterFly1_15_conc_2_itm_8_0 OR (butterFly1_15_conc_2_itm_8_2_1(1));
  mux_tmp_50 <= MUX_s_1_2_2(not_tmp_91, or_tmp_122, or_419_nl);
  and_dcpl_101 <= NOT(CONV_SL_1_1(butterFly2_15_conc_2_itm_8_2_1/=STD_LOGIC_VECTOR'("00")));
  and_dcpl_102 <= butterFly1_15_conc_2_itm_9_0 AND (NOT butterFly2_15_conc_2_itm_8_0);
  and_dcpl_104 <= NOT(butterFly1_15_conc_2_itm_8_0 OR (butterFly1_15_conc_2_itm_8_2_1(0)));
  and_dcpl_105 <= butterFly2_15_conc_2_itm_5_0 AND (NOT (butterFly1_15_conc_2_itm_8_2_1(1)));
  and_dcpl_107 <= (INNER_LOOP4_r_11_4_sva_6_0(6)) AND (NOT (INNER_LOOP4_r_11_4_sva_6_0(4)));
  nor_tmp_25 <= butterFly2_15_conc_2_itm_8_0 AND butterFly1_15_conc_2_itm_9_0;
  nor_52_nl <= NOT((NOT((butterFly2_15_conc_2_itm_8_2_1(1)) OR (NOT butterFly2_15_conc_2_itm_8_0)
      OR (NOT butterFly1_15_conc_2_itm_9_0))) OR nor_tmp_1);
  or_427_nl <= (butterFly2_15_conc_2_itm_8_2_1(1)) OR (NOT nor_tmp_25);
  mux_tmp_53 <= MUX_s_1_2_2(nor_52_nl, or_427_nl, butterFly2_15_conc_2_itm_9_2_1(1));
  or_429_nl <= (NOT butterFly1_15_conc_2_itm_8_0) OR (butterFly1_15_conc_2_itm_8_2_1(1));
  mux_tmp_56 <= MUX_s_1_2_2(not_tmp_91, or_tmp_122, or_429_nl);
  or_tmp_133 <= (NOT butterFly1_15_conc_2_itm_8_0) OR (butterFly1_15_conc_2_itm_8_2_1(1))
      OR (NOT butterFly2_15_conc_2_itm_5_0);
  and_dcpl_112 <= butterFly1_15_conc_2_itm_8_0 AND (NOT (butterFly1_15_conc_2_itm_8_2_1(0)));
  and_dcpl_114 <= CONV_SL_1_1(butterFly2_15_conc_2_itm_8_2_1=STD_LOGIC_VECTOR'("01"));
  and_dcpl_116 <= (NOT butterFly1_15_conc_2_itm_8_0) AND (butterFly1_15_conc_2_itm_8_2_1(0));
  and_dcpl_123 <= butterFly1_15_conc_2_itm_8_0 AND (butterFly1_15_conc_2_itm_8_2_1(0));
  or_447_nl <= (NOT (butterFly2_15_conc_2_itm_8_2_1(1))) OR butterFly2_15_conc_2_itm_8_0
      OR (NOT butterFly1_15_conc_2_itm_9_0);
  or_445_nl <= (NOT (butterFly2_15_conc_2_itm_8_2_1(1))) OR butterFly2_15_conc_2_itm_8_0;
  mux_69_nl <= MUX_s_1_2_2(not_tmp_87, or_tmp_112, or_445_nl);
  mux_tmp_70 <= MUX_s_1_2_2(or_447_nl, mux_69_nl, butterFly2_15_conc_2_itm_9_2_1(1));
  nor_tmp_32 <= (butterFly1_15_conc_2_itm_8_2_1(1)) AND butterFly2_15_conc_2_itm_5_0;
  or_tmp_153 <= butterFly1_15_conc_2_itm_8_0 OR (NOT nor_tmp_32);
  not_tmp_115 <= NOT((NOT(butterFly1_15_conc_2_itm_8_0 OR (NOT (butterFly1_15_conc_2_itm_8_2_1(1)))
      OR (NOT butterFly2_15_conc_2_itm_5_0))) OR nor_tmp_10);
  or_tmp_156 <= (INNER_LOOP2_r_11_4_sva_6_0(4)) OR (NOT(CONV_SL_1_1(INNER_LOOP2_r_11_4_sva_6_0(6
      DOWNTO 5)=STD_LOGIC_VECTOR'("11")) AND INNER_LOOP1_stage_0));
  and_dcpl_125 <= CONV_SL_1_1(butterFly2_15_conc_2_itm_8_2_1=STD_LOGIC_VECTOR'("10"));
  nor_tmp_36 <= (butterFly2_15_conc_2_itm_8_2_1(1)) AND butterFly2_15_conc_2_itm_8_0
      AND butterFly1_15_conc_2_itm_9_0;
  or_457_nl <= nor_tmp_36 OR nor_tmp_1;
  mux_tmp_78 <= MUX_s_1_2_2(nor_tmp_36, or_457_nl, butterFly2_15_conc_2_itm_9_2_1(1));
  and_8919_cse <= butterFly1_15_conc_2_itm_8_0 AND (butterFly1_15_conc_2_itm_8_2_1(1))
      AND butterFly2_15_conc_2_itm_5_0;
  or_tmp_160 <= and_8919_cse OR nor_tmp_10;
  nor_tmp_43 <= CONV_SL_1_1(INNER_LOOP4_r_11_4_sva_6_0(6 DOWNTO 4)=STD_LOGIC_VECTOR'("111"))
      AND INNER_LOOP1_stage_0;
  nor_tmp_45 <= CONV_SL_1_1(INNER_LOOP2_r_11_4_sva_6_0(6 DOWNTO 4)=STD_LOGIC_VECTOR'("111"))
      AND INNER_LOOP1_stage_0;
  nor_tmp_46 <= CONV_SL_1_1(butterFly2_15_conc_2_itm_8_2_1=STD_LOGIC_VECTOR'("11"))
      AND butterFly2_15_conc_2_itm_8_0 AND butterFly1_15_conc_2_itm_9_0;
  and_dcpl_135 <= INNER_LOOP2_stage_0_10 AND (NOT (butterFly1_15_conc_2_itm_9_2_1(1)));
  and_dcpl_138 <= INNER_LOOP1_stage_0 AND (NOT (INNER_LOOP3_r_11_4_sva_6_0(4)));
  and_dcpl_141 <= INNER_LOOP1_stage_0 AND (NOT (INNER_LOOP1_r_11_4_sva_6_0(4)));
  and_dcpl_145 <= INNER_LOOP1_stage_0 AND (INNER_LOOP3_r_11_4_sva_6_0(4));
  and_dcpl_147 <= INNER_LOOP1_stage_0 AND (INNER_LOOP1_r_11_4_sva_6_0(4));
  and_dcpl_150 <= INNER_LOOP2_stage_0_10 AND (butterFly1_15_conc_2_itm_9_2_1(1));
  and_dcpl_152 <= CONV_SL_1_1(INNER_LOOP3_r_11_4_sva_6_0(6 DOWNTO 5)=STD_LOGIC_VECTOR'("01"));
  and_dcpl_154 <= CONV_SL_1_1(INNER_LOOP1_r_11_4_sva_6_0(6 DOWNTO 5)=STD_LOGIC_VECTOR'("01"));
  and_dcpl_161 <= CONV_SL_1_1(INNER_LOOP3_r_11_4_sva_6_0(6 DOWNTO 5)=STD_LOGIC_VECTOR'("10"));
  and_dcpl_163 <= CONV_SL_1_1(INNER_LOOP1_r_11_4_sva_6_0(6 DOWNTO 5)=STD_LOGIC_VECTOR'("10"));
  and_dcpl_167 <= CONV_SL_1_1(INNER_LOOP3_r_11_4_sva_6_0(6 DOWNTO 5)=STD_LOGIC_VECTOR'("11"));
  and_dcpl_169 <= CONV_SL_1_1(INNER_LOOP1_r_11_4_sva_6_0(6 DOWNTO 5)=STD_LOGIC_VECTOR'("11"));
  or_dcpl_298 <= (fsm_output(7)) OR (fsm_output(9));
  or_dcpl_300 <= modulo_add_1_qelse_or_m1c OR or_dcpl_298;
  and_dcpl_173 <= INNER_LOOP1_stage_0 AND (operator_20_false_acc_cse_sva(0));
  and_dcpl_175 <= INNER_LOOP1_stage_0 AND (operator_20_false_acc_cse_sva(1));
  and_dcpl_176 <= INNER_LOOP1_stage_0 AND (operator_33_true_3_lshift_psp_1_0_sva(1));
  or_dcpl_315 <= CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("00"));
  and_dcpl_239 <= NOT((fsm_output(4)) OR (fsm_output(2)));
  or_dcpl_353 <= (fsm_output(2)) OR (fsm_output(7));
  or_dcpl_361 <= (fsm_output(4)) OR (fsm_output(7));
  or_329_cse <= (butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1(2)) OR (butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1(0));
  or_332_nl <= CONV_SL_1_1(INNER_LOOP4_r_11_4_sva_6_0(6 DOWNTO 4)/=STD_LOGIC_VECTOR'("000"));
  mux_3_nl <= MUX_s_1_2_2(not_tmp_25, or_tmp_35, or_332_nl);
  or_331_nl <= CONV_SL_1_1(INNER_LOOP4_r_11_4_sva_6_0(6 DOWNTO 4)/=STD_LOGIC_VECTOR'("000"))
      OR (NOT INNER_LOOP1_stage_0);
  mux_4_nl <= MUX_s_1_2_2(mux_3_nl, or_331_nl, or_329_cse);
  and_344_cse <= (NOT mux_4_nl) AND (fsm_output(9));
  and_346_cse <= (NOT(((butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1(2)) OR
      (butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1(0)) OR (NOT butterFly2_15_conc_2_itm_7_0)
      OR (butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1(1))) AND (CONV_SL_1_1(INNER_LOOP2_r_11_4_sva_6_0(6
      DOWNTO 4)/=STD_LOGIC_VECTOR'("000")) OR (NOT INNER_LOOP1_stage_0)))) AND (fsm_output(4));
  or_359_nl <= CONV_SL_1_1(INNER_LOOP4_r_11_4_sva_6_0(6 DOWNTO 4)/=STD_LOGIC_VECTOR'("001"))
      OR (NOT INNER_LOOP1_stage_0);
  or_357_nl <= CONV_SL_1_1(INNER_LOOP4_r_11_4_sva_6_0(6 DOWNTO 4)/=STD_LOGIC_VECTOR'("001"));
  mux_14_nl <= MUX_s_1_2_2(not_tmp_25, or_tmp_35, or_357_nl);
  nor_3_nl <= NOT((butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1(2)) OR (NOT
      (butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1(0))));
  mux_15_nl <= MUX_s_1_2_2(or_359_nl, mux_14_nl, nor_3_nl);
  and_715_cse <= (NOT mux_15_nl) AND (fsm_output(9));
  and_717_cse <= (NOT(((butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1(2)) OR
      (NOT (butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1(0))) OR (NOT butterFly2_15_conc_2_itm_7_0)
      OR (butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1(1))) AND (CONV_SL_1_1(INNER_LOOP2_r_11_4_sva_6_0(6
      DOWNTO 4)/=STD_LOGIC_VECTOR'("001")) OR (NOT INNER_LOOP1_stage_0)))) AND (fsm_output(4));
  nor_7_nl <= NOT(CONV_SL_1_1(INNER_LOOP4_r_11_4_sva_6_0(6 DOWNTO 4)/=STD_LOGIC_VECTOR'("010")));
  mux_25_nl <= MUX_s_1_2_2(and_8932_cse, or_tmp_82, nor_7_nl);
  nor_64_nl <= NOT((INNER_LOOP4_r_11_4_sva_6_0(4)) OR (INNER_LOOP4_r_11_4_sva_6_0(6))
      OR (NOT nor_tmp_6));
  mux_26_nl <= MUX_s_1_2_2(mux_25_nl, nor_64_nl, or_329_cse);
  and_1022_cse <= mux_26_nl AND (fsm_output(9));
  nand_24_cse <= NOT(butterFly2_15_conc_2_itm_7_0 AND (butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1(1)));
  and_8944_nl <= nand_24_cse AND or_tmp_90;
  mux_29_nl <= MUX_s_1_2_2(and_8944_nl, or_tmp_90, or_329_cse);
  and_1024_cse <= (NOT mux_29_nl) AND (fsm_output(4));
  nor_20_nl <= NOT(CONV_SL_1_1(INNER_LOOP4_r_11_4_sva_6_0(6 DOWNTO 4)/=STD_LOGIC_VECTOR'("011")));
  mux_35_nl <= MUX_s_1_2_2(and_8932_cse, or_tmp_82, nor_20_nl);
  mux_36_nl <= MUX_s_1_2_2((NOT or_tmp_99), mux_35_nl, butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1(0));
  mux_37_nl <= MUX_s_1_2_2(mux_36_nl, (NOT or_tmp_99), butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1(2));
  and_1329_cse <= mux_37_nl AND (fsm_output(9));
  and_8943_nl <= (NOT((butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1(0)) AND
      butterFly2_15_conc_2_itm_7_0 AND (butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1(1))))
      AND or_tmp_104;
  mux_40_nl <= MUX_s_1_2_2(and_8943_nl, or_tmp_104, butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1(2));
  and_1331_cse <= (NOT mux_40_nl) AND (fsm_output(4));
  or_412_cse <= (NOT (butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1(2))) OR (butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1(0));
  or_415_nl <= CONV_SL_1_1(INNER_LOOP4_r_11_4_sva_6_0(6 DOWNTO 4)/=STD_LOGIC_VECTOR'("100"));
  mux_48_nl <= MUX_s_1_2_2(not_tmp_25, or_tmp_35, or_415_nl);
  or_414_nl <= CONV_SL_1_1(INNER_LOOP4_r_11_4_sva_6_0(6 DOWNTO 4)/=STD_LOGIC_VECTOR'("100"))
      OR (NOT INNER_LOOP1_stage_0);
  mux_49_nl <= MUX_s_1_2_2(mux_48_nl, or_414_nl, or_412_cse);
  and_1636_cse <= (NOT mux_49_nl) AND (fsm_output(9));
  and_1638_cse <= (NOT(((NOT (butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1(2)))
      OR (butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1(0)) OR (NOT butterFly2_15_conc_2_itm_7_0)
      OR (butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1(1))) AND (CONV_SL_1_1(INNER_LOOP2_r_11_4_sva_6_0(6
      DOWNTO 4)/=STD_LOGIC_VECTOR'("100")) OR (NOT INNER_LOOP1_stage_0)))) AND (fsm_output(4));
  and_8941_cse <= (butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1(2)) AND (butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1(0));
  nand_17_nl <= NOT(CONV_SL_1_1(INNER_LOOP4_r_11_4_sva_6_0(6 DOWNTO 4)=STD_LOGIC_VECTOR'("101"))
      AND INNER_LOOP1_stage_0);
  or_434_nl <= CONV_SL_1_1(INNER_LOOP4_r_11_4_sva_6_0(6 DOWNTO 4)/=STD_LOGIC_VECTOR'("101"));
  mux_61_nl <= MUX_s_1_2_2(not_tmp_25, or_tmp_35, or_434_nl);
  mux_62_nl <= MUX_s_1_2_2(nand_17_nl, mux_61_nl, and_8941_cse);
  and_2007_cse <= (NOT mux_62_nl) AND (fsm_output(9));
  and_2009_cse <= (NOT((NOT((butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1(2))
      AND (butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1(0)) AND butterFly2_15_conc_2_itm_7_0
      AND (NOT (butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1(1))))) AND (NOT(CONV_SL_1_1(INNER_LOOP2_r_11_4_sva_6_0(6
      DOWNTO 4)=STD_LOGIC_VECTOR'("101")) AND INNER_LOOP1_stage_0)))) AND (fsm_output(4));
  nor_31_nl <= NOT(CONV_SL_1_1(INNER_LOOP4_r_11_4_sva_6_0(6 DOWNTO 4)/=STD_LOGIC_VECTOR'("110")));
  mux_73_nl <= MUX_s_1_2_2(and_8932_cse, or_tmp_82, nor_31_nl);
  nor_63_nl <= NOT((INNER_LOOP4_r_11_4_sva_6_0(4)) OR (NOT(CONV_SL_1_1(INNER_LOOP4_r_11_4_sva_6_0(6
      DOWNTO 5)=STD_LOGIC_VECTOR'("11")) AND INNER_LOOP1_stage_0)));
  mux_74_nl <= MUX_s_1_2_2(mux_73_nl, nor_63_nl, or_412_cse);
  and_2314_cse <= mux_74_nl AND (fsm_output(9));
  and_8942_nl <= nand_24_cse AND or_tmp_156;
  mux_77_nl <= MUX_s_1_2_2(and_8942_nl, or_tmp_156, or_412_cse);
  and_2316_cse <= (NOT mux_77_nl) AND (fsm_output(4));
  mux_85_nl <= MUX_s_1_2_2(and_8932_cse, or_tmp_82, butterFly2_16_f1_butterFly2_16_f1_and_6_cse);
  mux_86_nl <= MUX_s_1_2_2(nor_tmp_43, mux_85_nl, and_8941_cse);
  and_2621_cse <= mux_86_nl AND (fsm_output(9));
  and_2623_cse <= (((butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1(2)) AND (butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1(0))
      AND butterFly2_15_conc_2_itm_7_0 AND (butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1(1)))
      OR nor_tmp_45) AND (fsm_output(4));
  and_6834_cse <= INNER_LOOP1_stage_0 AND (operator_33_true_3_lshift_psp_1_0_sva(0))
      AND (fsm_output(9));
  and_6843_cse <= and_dcpl_176 AND (fsm_output(9));
  and_6852_cse <= and_dcpl_176 AND (operator_33_true_3_lshift_psp_1_0_sva(0)) AND
      (fsm_output(9));
  or_tmp_3231 <= modulo_add_1_qelse_or_m1c OR (fsm_output(9));
  and_7090_cse <= (NOT (operator_33_true_3_lshift_psp_1_0_sva(0))) AND (fsm_output(9));
  or_tmp_3239 <= and_7090_cse OR modulo_add_1_qelse_or_m1c;
  or_tmp_3242 <= (operator_33_true_3_lshift_psp_1_0_sva(0)) AND (fsm_output(9));
  and_7109_cse <= (NOT (operator_33_true_3_lshift_psp_1_0_sva(1))) AND (fsm_output(9));
  or_tmp_3250 <= (operator_20_false_acc_cse_sva(2)) AND (fsm_output(7));
  and_7115_cse <= (NOT (operator_20_false_acc_cse_sva(2))) AND (fsm_output(7));
  or_tmp_3252 <= (operator_33_true_3_lshift_psp_1_0_sva(1)) AND (fsm_output(9));
  or_tmp_3269 <= (operator_20_false_acc_cse_sva(1)) AND (fsm_output(7));
  and_7153_cse <= (NOT (operator_20_false_acc_cse_sva(1))) AND (fsm_output(7));
  or_tmp_3279 <= (operator_20_false_acc_cse_sva(0)) AND (fsm_output(7));
  and_7173_cse <= (NOT (operator_20_false_acc_cse_sva(0))) AND (fsm_output(7));
  or_tmp_3345 <= and_7153_cse OR modulo_add_1_qelse_or_m1c;
  or_tmp_3354 <= and_7173_cse OR modulo_add_1_qelse_or_m1c;
  or_tmp_3597 <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("00"));
  or_tmp_3600 <= CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00"));
  or_tmp_3650 <= and_dcpl_239 AND (NOT (fsm_output(7))) AND (NOT (fsm_output(9)));
  or_tmp_3666 <= (fsm_output(2)) OR (fsm_output(9));
  or_tmp_3717 <= NOT((fsm_output(2)) OR (fsm_output(7)));
  or_tmp_3723 <= NOT((fsm_output(6)) OR (fsm_output(2)) OR (fsm_output(7)));
  or_tmp_3732 <= CONV_SL_1_1(fsm_output(9 DOWNTO 8)/=STD_LOGIC_VECTOR'("00"));
  or_tmp_3755 <= (fsm_output(4)) OR (fsm_output(9));
  or_tmp_3842 <= or_dcpl_361 OR (fsm_output(9));
  INNER_LOOP1_tw_and_nl <= INNER_LOOP2_r_11_4_sva_6_0 AND INNER_LOOP1_r_11_4_sva_6_0;
  INNER_LOOP2_tw_and_nl <= operator_33_true_1_lshift_psp_9_4_sva AND (INNER_LOOP2_r_11_4_sva_6_0(5
      DOWNTO 0));
  INNER_LOOP1_tw_h_mux1h_4_rmff <= MUX1HOT_v_7_4_2(INNER_LOOP1_tw_and_nl, ((INNER_LOOP2_r_11_4_sva_6_0(6))
      & INNER_LOOP2_tw_and_nl), INNER_LOOP3_r_11_4_sva_6_0, INNER_LOOP4_r_11_4_sva_6_0,
      STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  butterFly1_and_ssc <= NOT((z_out_111(31)) OR (fsm_output(7)));
  butterFly1_and_ssc_2 <= (NOT (z_out_125(31))) AND (fsm_output(7));
  butterFly1_1_and_ssc <= NOT((z_out_112(31)) OR (fsm_output(7)));
  butterFly1_1_and_ssc_2 <= (NOT (z_out_126(31))) AND (fsm_output(7));
  butterFly1_1_and_ssc_3 <= (z_out_126(31)) AND (fsm_output(7));
  butterFly1_2_and_ssc <= NOT((z_out_113(31)) OR (fsm_output(7)));
  butterFly1_2_and_ssc_2 <= (NOT (z_out_111(31))) AND (fsm_output(7));
  butterFly1_2_and_ssc_3 <= (z_out_111(31)) AND (fsm_output(7));
  butterFly1_3_and_ssc <= NOT((z_out_114(31)) OR (fsm_output(7)));
  butterFly1_3_and_ssc_2 <= (NOT (z_out_112(31))) AND (fsm_output(7));
  butterFly1_3_and_ssc_3 <= (z_out_112(31)) AND (fsm_output(7));
  butterFly1_4_and_ssc <= NOT((z_out_115(31)) OR (fsm_output(7)));
  butterFly1_4_and_ssc_2 <= (NOT (z_out_113(31))) AND (fsm_output(7));
  butterFly1_4_and_ssc_3 <= (z_out_113(31)) AND (fsm_output(7));
  butterFly1_5_and_ssc <= NOT((z_out_116(31)) OR (fsm_output(7)));
  butterFly1_5_and_ssc_2 <= (NOT (z_out_114(31))) AND (fsm_output(7));
  butterFly1_5_and_ssc_3 <= (z_out_114(31)) AND (fsm_output(7));
  butterFly1_6_and_ssc <= NOT((z_out_117(31)) OR (fsm_output(7)));
  butterFly1_6_and_ssc_2 <= (NOT (z_out_115(31))) AND (fsm_output(7));
  butterFly1_6_and_ssc_3 <= (z_out_115(31)) AND (fsm_output(7));
  butterFly1_7_and_ssc <= NOT((z_out_118(31)) OR (fsm_output(7)));
  butterFly1_7_and_ssc_2 <= (NOT (z_out_116(31))) AND (fsm_output(7));
  butterFly1_7_and_ssc_3 <= (z_out_116(31)) AND (fsm_output(7));
  butterFly1_8_and_ssc <= NOT((z_out_119(31)) OR (fsm_output(7)));
  butterFly1_8_and_ssc_2 <= (NOT (z_out_117(31))) AND (fsm_output(7));
  butterFly1_8_and_ssc_3 <= (z_out_117(31)) AND (fsm_output(7));
  butterFly1_9_and_ssc <= NOT((z_out_120(31)) OR (fsm_output(7)));
  butterFly1_9_and_ssc_2 <= (NOT (z_out_118(31))) AND (fsm_output(7));
  butterFly1_9_and_ssc_3 <= (z_out_118(31)) AND (fsm_output(7));
  butterFly1_10_and_ssc <= NOT((z_out_121(31)) OR (fsm_output(7)));
  butterFly1_10_and_ssc_2 <= (NOT (z_out_119(31))) AND (fsm_output(7));
  butterFly1_10_and_ssc_3 <= (z_out_119(31)) AND (fsm_output(7));
  butterFly1_11_and_ssc <= NOT((z_out_122(31)) OR (fsm_output(7)));
  butterFly1_11_and_ssc_2 <= (NOT (z_out_120(31))) AND (fsm_output(7));
  butterFly1_11_and_ssc_3 <= (z_out_120(31)) AND (fsm_output(7));
  butterFly1_12_and_ssc <= NOT((z_out_123(31)) OR (fsm_output(7)));
  butterFly1_12_and_ssc_2 <= (NOT (z_out_121(31))) AND (fsm_output(7));
  butterFly1_12_and_ssc_3 <= (z_out_121(31)) AND (fsm_output(7));
  butterFly1_13_and_ssc <= NOT((z_out_124(31)) OR (fsm_output(7)));
  butterFly1_13_and_ssc_2 <= (NOT (z_out_122(31))) AND (fsm_output(7));
  butterFly1_13_and_ssc_3 <= (z_out_122(31)) AND (fsm_output(7));
  butterFly1_14_and_ssc <= NOT((z_out_125(31)) OR (fsm_output(7)));
  butterFly1_14_and_ssc_2 <= (NOT (z_out_123(31))) AND (fsm_output(7));
  butterFly1_14_and_ssc_3 <= (z_out_123(31)) AND (fsm_output(7));
  butterFly1_15_and_ssc <= NOT((z_out_126(31)) OR (fsm_output(7)));
  butterFly1_15_and_ssc_2 <= (NOT (z_out_124(31))) AND (fsm_output(7));
  yt_rsc_0_0_i_d_d_pff <= MUX_v_32_2_2(modulo_add_31_qr_lpi_3_dfm_1, modulo_add_10_qr_lpi_3_dfm_1,
      fsm_output(7));
  yt_rsc_0_0_i_radr_d_pff <= MUX_v_4_2_2((INNER_LOOP2_r_11_4_sva_6_0(3 DOWNTO 0)),
      (INNER_LOOP4_r_11_4_sva_6_0(3 DOWNTO 0)), fsm_output(9));
  yt_rsc_0_0_i_wadr_d_pff <= MUX_v_4_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_8450_itm_9,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_8833_itm_8, fsm_output(7));
  yt_rsc_0_0_i_we_d_pff <= (and_dcpl_68 AND (fsm_output(7))) OR (and_dcpl_70 AND
      and_dcpl_69 AND (fsm_output(2)));
  yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_pff <= (and_dcpl_73 AND butterFly2_16_f1_nor_1_cse
      AND (fsm_output(9))) OR (and_dcpl_76 AND (NOT (INNER_LOOP2_r_11_4_sva_6_0(6)))
      AND (NOT (INNER_LOOP2_r_11_4_sva_6_0(4))) AND (fsm_output(4)));
  yt_rsc_0_1_i_d_d_pff <= MUX_v_32_2_2(modulo_add_1_qr_lpi_3_dfm_1, modulo_add_11_qr_lpi_3_dfm_1,
      fsm_output(7));
  yt_rsc_0_1_i_wadr_d_pff <= MUX_v_4_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_8961_itm_9,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_9344_itm_8, fsm_output(7));
  yt_rsc_0_2_i_d_d_pff <= MUX_v_32_2_2(modulo_add_23_qr_lpi_3_dfm_1, modulo_add_12_qr_lpi_3_dfm_1,
      fsm_output(7));
  yt_rsc_0_2_i_wadr_d_pff <= MUX_v_4_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_9472_itm_9,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_9855_itm_8, fsm_output(7));
  yt_rsc_0_3_i_d_d_pff <= MUX_v_32_2_2(modulo_add_24_qr_lpi_3_dfm_1, modulo_add_13_qr_lpi_3_dfm_1,
      fsm_output(7));
  yt_rsc_0_3_i_wadr_d_pff <= MUX_v_4_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_10015_itm_9,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_10366_itm_8, fsm_output(7));
  yt_rsc_0_4_i_d_d_pff <= MUX_v_32_2_2(modulo_add_25_qr_lpi_3_dfm_1, modulo_add_14_qr_lpi_3_dfm_1,
      fsm_output(7));
  yt_rsc_0_4_i_wadr_d_pff <= MUX_v_4_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_10494_itm_9,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_10877_itm_8, fsm_output(7));
  yt_rsc_0_5_i_d_d_pff <= MUX_v_32_2_2(modulo_add_26_qr_lpi_3_dfm_1, modulo_add_15_qr_lpi_3_dfm_1,
      fsm_output(7));
  yt_rsc_0_5_i_wadr_d_pff <= MUX_v_4_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_11005_itm_9,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_11388_itm_8, fsm_output(7));
  yt_rsc_0_6_i_d_d_pff <= MUX_v_32_2_2(modulo_add_27_qr_lpi_3_dfm_1, modulo_add_1_qr_lpi_3_dfm_1,
      fsm_output(7));
  yt_rsc_0_6_i_wadr_d_pff <= MUX_v_4_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_11516_itm_9,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_11899_itm_8, fsm_output(7));
  yt_rsc_0_7_i_d_d_pff <= MUX_v_32_2_2(modulo_add_28_qr_lpi_3_dfm_1, modulo_add_23_qr_lpi_3_dfm_1,
      fsm_output(7));
  yt_rsc_0_8_i_d_d_pff <= MUX_v_32_2_2(modulo_add_29_qr_lpi_3_dfm_1, modulo_add_24_qr_lpi_3_dfm_1,
      fsm_output(7));
  yt_rsc_0_9_i_d_d_pff <= MUX_v_32_2_2(modulo_add_30_qr_lpi_3_dfm_1, modulo_add_25_qr_lpi_3_dfm_1,
      fsm_output(7));
  yt_rsc_0_10_i_d_d_pff <= MUX_v_32_2_2(modulo_add_10_qr_lpi_3_dfm_1, modulo_add_26_qr_lpi_3_dfm_1,
      fsm_output(7));
  yt_rsc_0_10_i_wadr_d_pff <= MUX_v_4_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13560_itm_9,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13943_itm_8, fsm_output(7));
  yt_rsc_0_11_i_d_d_pff <= MUX_v_32_2_2(modulo_add_11_qr_lpi_3_dfm_1, modulo_add_27_qr_lpi_3_dfm_1,
      fsm_output(7));
  yt_rsc_0_11_i_wadr_d_pff <= MUX_v_4_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14071_itm_9,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14454_itm_8, fsm_output(7));
  yt_rsc_0_12_i_d_d_pff <= MUX_v_32_2_2(modulo_add_12_qr_lpi_3_dfm_1, modulo_add_28_qr_lpi_3_dfm_1,
      fsm_output(7));
  yt_rsc_0_13_i_d_d_pff <= MUX_v_32_2_2(modulo_add_13_qr_lpi_3_dfm_1, modulo_add_29_qr_lpi_3_dfm_1,
      fsm_output(7));
  yt_rsc_0_14_i_d_d_pff <= MUX_v_32_2_2(modulo_add_14_qr_lpi_3_dfm_1, modulo_add_30_qr_lpi_3_dfm_1,
      fsm_output(7));
  yt_rsc_0_15_i_d_d_pff <= MUX_v_32_2_2(modulo_add_15_qr_lpi_3_dfm_1, modulo_add_31_qr_lpi_3_dfm_1,
      fsm_output(7));
  yt_rsc_0_16_i_we_d_pff <= (and_dcpl_78 AND (fsm_output(7))) OR (and_dcpl_70 AND
      and_dcpl_79 AND (fsm_output(2)));
  yt_rsc_1_0_i_we_d_pff <= (and_dcpl_82 AND (fsm_output(7))) OR (and_dcpl_70 AND
      and_dcpl_83 AND (fsm_output(2)));
  yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_pff <= (and_dcpl_73 AND (NOT (INNER_LOOP4_r_11_4_sva_6_0(6)))
      AND (INNER_LOOP4_r_11_4_sva_6_0(4)) AND (fsm_output(9))) OR (and_dcpl_76 AND
      (NOT (INNER_LOOP2_r_11_4_sva_6_0(6))) AND (INNER_LOOP2_r_11_4_sva_6_0(4)) AND
      (fsm_output(4)));
  yt_rsc_1_16_i_we_d_pff <= (and_dcpl_89 AND (fsm_output(7))) OR (and_dcpl_70 AND
      and_8912_cse AND (fsm_output(2)));
  yt_rsc_2_0_i_we_d_pff <= (and_dcpl_93 AND (fsm_output(7))) OR (nor_tmp_10 AND and_dcpl_69
      AND (fsm_output(2)));
  yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_pff <= (nor_tmp_6 AND butterFly2_16_f1_nor_1_cse
      AND (fsm_output(9))) OR ((NOT or_tmp_90) AND (fsm_output(4)));
  yt_rsc_2_16_i_we_d_pff <= (and_dcpl_96 AND (fsm_output(7))) OR (nor_tmp_10 AND
      and_dcpl_79 AND (fsm_output(2)));
  yt_rsc_3_0_i_we_d_pff <= (and_dcpl_99 AND (fsm_output(7))) OR (nor_tmp_10 AND and_dcpl_83
      AND (fsm_output(2)));
  yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_pff <= ((NOT or_tmp_99) AND (fsm_output(9)))
      OR ((NOT or_tmp_104) AND (fsm_output(4)));
  yt_rsc_3_16_i_we_d_pff <= (nor_tmp_22 AND (fsm_output(7))) OR (and_8913_cse AND
      (fsm_output(2)));
  butterFly1_and_4_nl <= (z_out_108(31)) AND (NOT(butterFly1_and_ssc OR butterFly1_and_ssc_2));
  butterFly1_or_nl <= ((z_out_111(31)) AND (NOT (fsm_output(7)))) OR ((z_out_125(31))
      AND (fsm_output(7)));
  butterFly1_mux1h_nl <= MUX1HOT_v_31_3_2((z_out_111(30 DOWNTO 0)), (z_out_108(30
      DOWNTO 0)), (z_out_125(30 DOWNTO 0)), STD_LOGIC_VECTOR'( butterFly1_and_ssc
      & butterFly1_or_nl & butterFly1_and_ssc_2));
  yt_rsc_4_0_i_d_d_pff <= butterFly1_and_4_nl & butterFly1_mux1h_nl;
  yt_rsc_4_0_i_wadr_d_pff <= MUX_v_4_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_8833_itm_8,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12538_itm_8, fsm_output(7));
  yt_rsc_4_0_i_we_d_pff <= (and_dcpl_102 AND and_dcpl_101 AND (fsm_output(7))) OR
      (and_dcpl_105 AND and_dcpl_104 AND (fsm_output(2)));
  yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_pff <= (and_dcpl_73 AND and_dcpl_107
      AND (fsm_output(9))) OR (and_dcpl_76 AND (INNER_LOOP2_r_11_4_sva_6_0(6)) AND
      (NOT (INNER_LOOP2_r_11_4_sva_6_0(4))) AND (fsm_output(4)));
  butterFly1_1_mux_nl <= MUX_s_1_2_2((z_out_102(31)), (z_out_105(31)), butterFly1_1_and_ssc_3);
  butterFly1_1_and_4_nl <= butterFly1_1_mux_nl AND (NOT(butterFly1_1_and_ssc OR butterFly1_1_and_ssc_2));
  butterFly1_1_and_1_nl <= (z_out_112(31)) AND (NOT (fsm_output(7)));
  butterFly1_1_mux1h_nl <= MUX1HOT_v_31_4_2((z_out_112(30 DOWNTO 0)), (z_out_102(30
      DOWNTO 0)), (z_out_126(30 DOWNTO 0)), (z_out_105(30 DOWNTO 0)), STD_LOGIC_VECTOR'(
      butterFly1_1_and_ssc & butterFly1_1_and_1_nl & butterFly1_1_and_ssc_2 & butterFly1_1_and_ssc_3));
  yt_rsc_4_1_i_d_d_pff <= butterFly1_1_and_4_nl & butterFly1_1_mux1h_nl;
  yt_rsc_4_1_i_wadr_d_pff <= MUX_v_4_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_9344_itm_8,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13049_itm_8, fsm_output(7));
  butterFly1_2_mux_nl <= MUX_s_1_2_2((z_out_97(31)), (z_out_100(31)), butterFly1_2_and_ssc_3);
  butterFly1_2_and_4_nl <= butterFly1_2_mux_nl AND (NOT(butterFly1_2_and_ssc OR butterFly1_2_and_ssc_2));
  butterFly1_2_and_1_nl <= (z_out_113(31)) AND (NOT (fsm_output(7)));
  butterFly1_2_mux1h_nl <= MUX1HOT_v_31_4_2((z_out_113(30 DOWNTO 0)), (z_out_97(30
      DOWNTO 0)), (z_out_111(30 DOWNTO 0)), (z_out_100(30 DOWNTO 0)), STD_LOGIC_VECTOR'(
      butterFly1_2_and_ssc & butterFly1_2_and_1_nl & butterFly1_2_and_ssc_2 & butterFly1_2_and_ssc_3));
  yt_rsc_4_2_i_d_d_pff <= butterFly1_2_and_4_nl & butterFly1_2_mux1h_nl;
  yt_rsc_4_2_i_wadr_d_pff <= MUX_v_4_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_9855_itm_8,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14582_itm_8, fsm_output(7));
  butterFly1_3_mux_nl <= MUX_s_1_2_2((z_out_92(31)), (z_out_94(31)), butterFly1_3_and_ssc_3);
  butterFly1_3_and_4_nl <= butterFly1_3_mux_nl AND (NOT(butterFly1_3_and_ssc OR butterFly1_3_and_ssc_2));
  butterFly1_3_and_1_nl <= (z_out_114(31)) AND (NOT (fsm_output(7)));
  butterFly1_3_mux1h_nl <= MUX1HOT_v_31_4_2((z_out_114(30 DOWNTO 0)), (z_out_92(30
      DOWNTO 0)), (z_out_112(30 DOWNTO 0)), (z_out_94(30 DOWNTO 0)), STD_LOGIC_VECTOR'(
      butterFly1_3_and_ssc & butterFly1_3_and_1_nl & butterFly1_3_and_ssc_2 & butterFly1_3_and_ssc_3));
  yt_rsc_4_3_i_d_d_pff <= butterFly1_3_and_4_nl & butterFly1_3_mux1h_nl;
  yt_rsc_4_3_i_wadr_d_pff <= MUX_v_4_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_10366_itm_8,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15093_itm_8, fsm_output(7));
  butterFly1_4_mux_nl <= MUX_s_1_2_2((z_out_86(31)), (z_out_89(31)), butterFly1_4_and_ssc_3);
  butterFly1_4_and_4_nl <= butterFly1_4_mux_nl AND (NOT(butterFly1_4_and_ssc OR butterFly1_4_and_ssc_2));
  butterFly1_4_and_1_nl <= (z_out_115(31)) AND (NOT (fsm_output(7)));
  butterFly1_4_mux1h_nl <= MUX1HOT_v_31_4_2((z_out_115(30 DOWNTO 0)), (z_out_86(30
      DOWNTO 0)), (z_out_113(30 DOWNTO 0)), (z_out_89(30 DOWNTO 0)), STD_LOGIC_VECTOR'(
      butterFly1_4_and_ssc & butterFly1_4_and_1_nl & butterFly1_4_and_ssc_2 & butterFly1_4_and_ssc_3));
  yt_rsc_4_4_i_d_d_pff <= butterFly1_4_and_4_nl & butterFly1_4_mux1h_nl;
  yt_rsc_4_4_i_wadr_d_pff <= MUX_v_4_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_10877_itm_8,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15604_itm_8, fsm_output(7));
  butterFly1_5_mux_nl <= MUX_s_1_2_2((z_out_81(31)), (z_out_84(31)), butterFly1_5_and_ssc_3);
  butterFly1_5_and_4_nl <= butterFly1_5_mux_nl AND (NOT(butterFly1_5_and_ssc OR butterFly1_5_and_ssc_2));
  butterFly1_5_and_1_nl <= (z_out_116(31)) AND (NOT (fsm_output(7)));
  butterFly1_5_mux1h_nl <= MUX1HOT_v_31_4_2((z_out_116(30 DOWNTO 0)), (z_out_81(30
      DOWNTO 0)), (z_out_114(30 DOWNTO 0)), (z_out_84(30 DOWNTO 0)), STD_LOGIC_VECTOR'(
      butterFly1_5_and_ssc & butterFly1_5_and_1_nl & butterFly1_5_and_ssc_2 & butterFly1_5_and_ssc_3));
  yt_rsc_4_5_i_d_d_pff <= butterFly1_5_and_4_nl & butterFly1_5_mux1h_nl;
  yt_rsc_4_5_i_wadr_d_pff <= MUX_v_4_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_11388_itm_8,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16115_itm_8, fsm_output(7));
  butterFly1_6_mux_nl <= MUX_s_1_2_2((z_out_76(31)), (z_out_78(31)), butterFly1_6_and_ssc_3);
  butterFly1_6_and_4_nl <= butterFly1_6_mux_nl AND (NOT(butterFly1_6_and_ssc OR butterFly1_6_and_ssc_2));
  butterFly1_6_and_1_nl <= (z_out_117(31)) AND (NOT (fsm_output(7)));
  butterFly1_6_mux1h_nl <= MUX1HOT_v_31_4_2((z_out_117(30 DOWNTO 0)), (z_out_76(30
      DOWNTO 0)), (z_out_115(30 DOWNTO 0)), (z_out_78(30 DOWNTO 0)), STD_LOGIC_VECTOR'(
      butterFly1_6_and_ssc & butterFly1_6_and_1_nl & butterFly1_6_and_ssc_2 & butterFly1_6_and_ssc_3));
  yt_rsc_4_6_i_d_d_pff <= butterFly1_6_and_4_nl & butterFly1_6_mux1h_nl;
  yt_rsc_4_6_i_wadr_d_pff <= MUX_v_4_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_11899_itm_8,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12027_itm_8, fsm_output(7));
  butterFly1_7_mux_nl <= MUX_s_1_2_2((z_out_70(31)), (z_out_73(31)), butterFly1_7_and_ssc_3);
  butterFly1_7_and_4_nl <= butterFly1_7_mux_nl AND (NOT(butterFly1_7_and_ssc OR butterFly1_7_and_ssc_2));
  butterFly1_7_and_1_nl <= (z_out_118(31)) AND (NOT (fsm_output(7)));
  butterFly1_7_mux1h_nl <= MUX1HOT_v_31_4_2((z_out_118(30 DOWNTO 0)), (z_out_70(30
      DOWNTO 0)), (z_out_116(30 DOWNTO 0)), (z_out_73(30 DOWNTO 0)), STD_LOGIC_VECTOR'(
      butterFly1_7_and_ssc & butterFly1_7_and_1_nl & butterFly1_7_and_ssc_2 & butterFly1_7_and_ssc_3));
  yt_rsc_4_7_i_d_d_pff <= butterFly1_7_and_4_nl & butterFly1_7_mux1h_nl;
  butterFly1_8_mux_nl <= MUX_s_1_2_2((z_out_105(31)), (z_out_102(31)), butterFly1_8_and_ssc_3);
  butterFly1_8_and_4_nl <= butterFly1_8_mux_nl AND (NOT(butterFly1_8_and_ssc OR butterFly1_8_and_ssc_2));
  butterFly1_8_and_1_nl <= (z_out_119(31)) AND (NOT (fsm_output(7)));
  butterFly1_8_mux1h_nl <= MUX1HOT_v_31_4_2((z_out_119(30 DOWNTO 0)), (z_out_105(30
      DOWNTO 0)), (z_out_117(30 DOWNTO 0)), (z_out_102(30 DOWNTO 0)), STD_LOGIC_VECTOR'(
      butterFly1_8_and_ssc & butterFly1_8_and_1_nl & butterFly1_8_and_ssc_2 & butterFly1_8_and_ssc_3));
  yt_rsc_4_8_i_d_d_pff <= butterFly1_8_and_4_nl & butterFly1_8_mux1h_nl;
  butterFly1_9_mux_nl <= MUX_s_1_2_2((z_out_100(31)), (z_out_97(31)), butterFly1_9_and_ssc_3);
  butterFly1_9_and_4_nl <= butterFly1_9_mux_nl AND (NOT(butterFly1_9_and_ssc OR butterFly1_9_and_ssc_2));
  butterFly1_9_and_1_nl <= (z_out_120(31)) AND (NOT (fsm_output(7)));
  butterFly1_9_mux1h_272_nl <= MUX1HOT_v_31_4_2((z_out_120(30 DOWNTO 0)), (z_out_100(30
      DOWNTO 0)), (z_out_118(30 DOWNTO 0)), (z_out_97(30 DOWNTO 0)), STD_LOGIC_VECTOR'(
      butterFly1_9_and_ssc & butterFly1_9_and_1_nl & butterFly1_9_and_ssc_2 & butterFly1_9_and_ssc_3));
  yt_rsc_4_9_i_d_d_pff <= butterFly1_9_and_4_nl & butterFly1_9_mux1h_272_nl;
  yt_rsc_4_9_i_wadr_d_pff <= MUX_v_4_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_9855_itm_8,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13560_itm_8, fsm_output(7));
  butterFly1_10_mux_nl <= MUX_s_1_2_2((z_out_94(31)), (z_out_92(31)), butterFly1_10_and_ssc_3);
  butterFly1_10_and_4_nl <= butterFly1_10_mux_nl AND (NOT(butterFly1_10_and_ssc OR
      butterFly1_10_and_ssc_2));
  butterFly1_10_and_1_nl <= (z_out_121(31)) AND (NOT (fsm_output(7)));
  butterFly1_10_mux1h_nl <= MUX1HOT_v_31_4_2((z_out_121(30 DOWNTO 0)), (z_out_94(30
      DOWNTO 0)), (z_out_119(30 DOWNTO 0)), (z_out_92(30 DOWNTO 0)), STD_LOGIC_VECTOR'(
      butterFly1_10_and_ssc & butterFly1_10_and_1_nl & butterFly1_10_and_ssc_2 &
      butterFly1_10_and_ssc_3));
  yt_rsc_4_10_i_d_d_pff <= butterFly1_10_and_4_nl & butterFly1_10_mux1h_nl;
  yt_rsc_4_10_i_wadr_d_pff <= MUX_v_4_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13943_itm_8,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14071_itm_8, fsm_output(7));
  butterFly1_11_mux_nl <= MUX_s_1_2_2((z_out_89(31)), (z_out_86(31)), butterFly1_11_and_ssc_3);
  butterFly1_11_and_4_nl <= butterFly1_11_mux_nl AND (NOT(butterFly1_11_and_ssc OR
      butterFly1_11_and_ssc_2));
  butterFly1_11_and_1_nl <= (z_out_122(31)) AND (NOT (fsm_output(7)));
  butterFly1_11_mux1h_nl <= MUX1HOT_v_31_4_2((z_out_122(30 DOWNTO 0)), (z_out_89(30
      DOWNTO 0)), (z_out_120(30 DOWNTO 0)), (z_out_86(30 DOWNTO 0)), STD_LOGIC_VECTOR'(
      butterFly1_11_and_ssc & butterFly1_11_and_1_nl & butterFly1_11_and_ssc_2 &
      butterFly1_11_and_ssc_3));
  yt_rsc_4_11_i_d_d_pff <= butterFly1_11_and_4_nl & butterFly1_11_mux1h_nl;
  yt_rsc_4_11_i_wadr_d_pff <= MUX_v_4_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14454_itm_8,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14582_itm_8, fsm_output(7));
  butterFly1_12_mux_nl <= MUX_s_1_2_2((z_out_84(31)), (z_out_81(31)), butterFly1_12_and_ssc_3);
  butterFly1_12_and_4_nl <= butterFly1_12_mux_nl AND (NOT(butterFly1_12_and_ssc OR
      butterFly1_12_and_ssc_2));
  butterFly1_12_and_1_nl <= (z_out_123(31)) AND (NOT (fsm_output(7)));
  butterFly1_12_mux1h_nl <= MUX1HOT_v_31_4_2((z_out_123(30 DOWNTO 0)), (z_out_84(30
      DOWNTO 0)), (z_out_121(30 DOWNTO 0)), (z_out_81(30 DOWNTO 0)), STD_LOGIC_VECTOR'(
      butterFly1_12_and_ssc & butterFly1_12_and_1_nl & butterFly1_12_and_ssc_2 &
      butterFly1_12_and_ssc_3));
  yt_rsc_4_12_i_d_d_pff <= butterFly1_12_and_4_nl & butterFly1_12_mux1h_nl;
  butterFly1_13_mux_nl <= MUX_s_1_2_2((z_out_78(31)), (z_out_76(31)), butterFly1_13_and_ssc_3);
  butterFly1_13_and_4_nl <= butterFly1_13_mux_nl AND (NOT(butterFly1_13_and_ssc OR
      butterFly1_13_and_ssc_2));
  butterFly1_13_and_1_nl <= (z_out_124(31)) AND (NOT (fsm_output(7)));
  butterFly1_13_mux1h_nl <= MUX1HOT_v_31_4_2((z_out_124(30 DOWNTO 0)), (z_out_78(30
      DOWNTO 0)), (z_out_122(30 DOWNTO 0)), (z_out_76(30 DOWNTO 0)), STD_LOGIC_VECTOR'(
      butterFly1_13_and_ssc & butterFly1_13_and_1_nl & butterFly1_13_and_ssc_2 &
      butterFly1_13_and_ssc_3));
  yt_rsc_4_13_i_d_d_pff <= butterFly1_13_and_4_nl & butterFly1_13_mux1h_nl;
  butterFly1_14_mux_nl <= MUX_s_1_2_2((z_out_73(31)), (z_out_70(31)), butterFly1_14_and_ssc_3);
  butterFly1_14_and_4_nl <= butterFly1_14_mux_nl AND (NOT(butterFly1_14_and_ssc OR
      butterFly1_14_and_ssc_2));
  butterFly1_14_and_1_nl <= (z_out_125(31)) AND (NOT (fsm_output(7)));
  butterFly1_14_mux1h_nl <= MUX1HOT_v_31_4_2((z_out_125(30 DOWNTO 0)), (z_out_73(30
      DOWNTO 0)), (z_out_123(30 DOWNTO 0)), (z_out_70(30 DOWNTO 0)), STD_LOGIC_VECTOR'(
      butterFly1_14_and_ssc & butterFly1_14_and_1_nl & butterFly1_14_and_ssc_2 &
      butterFly1_14_and_ssc_3));
  yt_rsc_4_14_i_d_d_pff <= butterFly1_14_and_4_nl & butterFly1_14_mux1h_nl;
  butterFly1_15_and_5_nl <= (z_out_68(31)) AND (NOT(butterFly1_15_and_ssc OR butterFly1_15_and_ssc_2));
  butterFly1_15_or_nl <= ((z_out_126(31)) AND (NOT (fsm_output(7)))) OR ((z_out_124(31))
      AND (fsm_output(7)));
  butterFly1_15_mux1h_nl <= MUX1HOT_v_31_3_2((z_out_126(30 DOWNTO 0)), (z_out_68(30
      DOWNTO 0)), (z_out_124(30 DOWNTO 0)), STD_LOGIC_VECTOR'( butterFly1_15_and_ssc
      & butterFly1_15_or_nl & butterFly1_15_and_ssc_2));
  yt_rsc_4_15_i_d_d_pff <= butterFly1_15_and_5_nl & butterFly1_15_mux1h_nl;
  yt_rsc_4_16_i_we_d_pff <= (nor_tmp_25 AND and_dcpl_101 AND (fsm_output(7))) OR
      (and_dcpl_105 AND and_dcpl_112 AND (fsm_output(2)));
  yt_rsc_5_0_i_we_d_pff <= (and_dcpl_102 AND and_dcpl_114 AND (fsm_output(7))) OR
      (and_dcpl_105 AND and_dcpl_116 AND (fsm_output(2)));
  yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_pff <= (and_dcpl_73 AND (INNER_LOOP4_r_11_4_sva_6_0(6))
      AND (INNER_LOOP4_r_11_4_sva_6_0(4)) AND (fsm_output(9))) OR (and_dcpl_76 AND
      (INNER_LOOP2_r_11_4_sva_6_0(6)) AND (INNER_LOOP2_r_11_4_sva_6_0(4)) AND (fsm_output(4)));
  yt_rsc_5_16_i_we_d_pff <= (nor_tmp_25 AND and_dcpl_114 AND (fsm_output(7))) OR
      (and_dcpl_105 AND and_dcpl_123 AND (fsm_output(2)));
  yt_rsc_6_0_i_we_d_pff <= (and_dcpl_102 AND and_dcpl_125 AND (fsm_output(7))) OR
      (nor_tmp_32 AND and_dcpl_104 AND (fsm_output(2)));
  yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_pff <= (nor_tmp_6 AND and_dcpl_107
      AND (fsm_output(9))) OR ((NOT or_tmp_156) AND (fsm_output(4)));
  yt_rsc_6_16_i_we_d_pff <= (nor_tmp_25 AND and_dcpl_125 AND (fsm_output(7))) OR
      (nor_tmp_32 AND and_dcpl_112 AND (fsm_output(2)));
  yt_rsc_7_0_i_we_d_pff <= (and_dcpl_102 AND CONV_SL_1_1(butterFly2_15_conc_2_itm_8_2_1=STD_LOGIC_VECTOR'("11"))
      AND (fsm_output(7))) OR (nor_tmp_32 AND and_dcpl_116 AND (fsm_output(2)));
  yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_pff <= (nor_tmp_43 AND (fsm_output(9)))
      OR (nor_tmp_45 AND (fsm_output(4)));
  yt_rsc_7_16_i_we_d_pff <= (nor_tmp_46 AND (fsm_output(7))) OR (nor_tmp_32 AND and_dcpl_123
      AND (fsm_output(2)));
  xt_rsc_0_0_i_adra_d_pff <= MUX1HOT_v_4_4_2((INNER_LOOP1_r_11_4_sva_6_0(3 DOWNTO
      0)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12538_itm_5, (INNER_LOOP3_r_11_4_sva_6_0(3
      DOWNTO 0)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12921_itm_5, STD_LOGIC_VECTOR'(
      (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  xt_rsc_0_0_i_da_d_pff <= modulo_add_10_qr_lpi_3_dfm_1;
  xt_rsc_0_0_i_wea_d_pff <= (and_dcpl_68 AND (fsm_output(9))) OR (and_dcpl_135 AND
      and_dcpl_69 AND (fsm_output(4)));
  xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff <= (and_dcpl_138 AND butterFly2_f1_nor_cse
      AND (fsm_output(7))) OR (and_dcpl_141 AND butterFly1_f1_nor_cse AND (fsm_output(2)));
  xt_rsc_0_1_i_adra_d_pff <= MUX1HOT_v_4_4_2((INNER_LOOP1_r_11_4_sva_6_0(3 DOWNTO
      0)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13049_itm_6, (INNER_LOOP3_r_11_4_sva_6_0(3
      DOWNTO 0)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13432_itm_6, STD_LOGIC_VECTOR'(
      (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  xt_rsc_0_1_i_da_d_pff <= modulo_add_11_qr_lpi_3_dfm_1;
  xt_rsc_0_2_i_adra_d_pff <= MUX1HOT_v_4_4_2((INNER_LOOP1_r_11_4_sva_6_0(3 DOWNTO
      0)), INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9472_itm_9, (INNER_LOOP3_r_11_4_sva_6_0(3
      DOWNTO 0)), INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9855_itm_9, STD_LOGIC_VECTOR'(
      (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  xt_rsc_0_2_i_da_d_pff <= modulo_add_12_qr_lpi_3_dfm_1;
  xt_rsc_0_3_i_adra_d_pff <= MUX1HOT_v_4_4_2((INNER_LOOP1_r_11_4_sva_6_0(3 DOWNTO
      0)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_10015_itm_9, (INNER_LOOP3_r_11_4_sva_6_0(3
      DOWNTO 0)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15093_itm_1, STD_LOGIC_VECTOR'(
      (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  xt_rsc_0_3_i_da_d_pff <= modulo_add_13_qr_lpi_3_dfm_1;
  xt_rsc_0_4_i_adra_d_pff <= MUX1HOT_v_4_4_2((INNER_LOOP1_r_11_4_sva_6_0(3 DOWNTO
      0)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15476_itm_1, (INNER_LOOP3_r_11_4_sva_6_0(3
      DOWNTO 0)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15604_itm_2, STD_LOGIC_VECTOR'(
      (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  xt_rsc_0_4_i_da_d_pff <= modulo_add_14_qr_lpi_3_dfm_1;
  xt_rsc_0_5_i_adra_d_pff <= MUX1HOT_v_4_4_2((INNER_LOOP1_r_11_4_sva_6_0(3 DOWNTO
      0)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15987_itm_2, (INNER_LOOP3_r_11_4_sva_6_0(3
      DOWNTO 0)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16115_itm_3, STD_LOGIC_VECTOR'(
      (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  xt_rsc_0_5_i_da_d_pff <= modulo_add_15_qr_lpi_3_dfm_1;
  xt_rsc_0_6_i_adra_d_pff <= MUX1HOT_v_4_4_2((INNER_LOOP1_r_11_4_sva_6_0(3 DOWNTO
      0)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16498_itm_3, (INNER_LOOP3_r_11_4_sva_6_0(3
      DOWNTO 0)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12027_itm_4, STD_LOGIC_VECTOR'(
      (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  xt_rsc_0_6_i_da_d_pff <= modulo_add_1_qr_lpi_3_dfm_1;
  xt_rsc_0_7_i_adra_d_pff <= MUX1HOT_v_4_4_2((INNER_LOOP1_r_11_4_sva_6_0(3 DOWNTO
      0)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12410_itm_4, (INNER_LOOP3_r_11_4_sva_6_0(3
      DOWNTO 0)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12538_itm_5, STD_LOGIC_VECTOR'(
      (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  xt_rsc_0_7_i_da_d_pff <= modulo_add_23_qr_lpi_3_dfm_1;
  xt_rsc_0_8_i_adra_d_pff <= MUX1HOT_v_4_4_2((INNER_LOOP1_r_11_4_sva_6_0(3 DOWNTO
      0)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12921_itm_5, (INNER_LOOP3_r_11_4_sva_6_0(3
      DOWNTO 0)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13049_itm_6, STD_LOGIC_VECTOR'(
      (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  xt_rsc_0_8_i_da_d_pff <= modulo_add_24_qr_lpi_3_dfm_1;
  xt_rsc_0_9_i_adra_d_pff <= MUX1HOT_v_4_4_2((INNER_LOOP1_r_11_4_sva_6_0(3 DOWNTO
      0)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13432_itm_6, (INNER_LOOP3_r_11_4_sva_6_0(3
      DOWNTO 0)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13560_itm_7, STD_LOGIC_VECTOR'(
      (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  xt_rsc_0_9_i_da_d_pff <= modulo_add_25_qr_lpi_3_dfm_1;
  xt_rsc_0_10_i_adra_d_pff <= MUX1HOT_v_4_4_2((INNER_LOOP1_r_11_4_sva_6_0(3 DOWNTO
      0)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13943_itm_7, (INNER_LOOP3_r_11_4_sva_6_0(3
      DOWNTO 0)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14071_itm_8, STD_LOGIC_VECTOR'(
      (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  xt_rsc_0_10_i_da_d_pff <= modulo_add_26_qr_lpi_3_dfm_1;
  xt_rsc_0_11_i_adra_d_pff <= MUX1HOT_v_4_4_2((INNER_LOOP1_r_11_4_sva_6_0(3 DOWNTO
      0)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14454_itm_8, (INNER_LOOP3_r_11_4_sva_6_0(3
      DOWNTO 0)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_10015_itm_9, STD_LOGIC_VECTOR'(
      (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  xt_rsc_0_11_i_da_d_pff <= modulo_add_27_qr_lpi_3_dfm_1;
  xt_rsc_0_12_i_adra_d_pff <= MUX1HOT_v_4_4_2((INNER_LOOP1_r_11_4_sva_6_0(3 DOWNTO
      0)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15093_itm_1, (INNER_LOOP3_r_11_4_sva_6_0(3
      DOWNTO 0)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15476_itm_1, STD_LOGIC_VECTOR'(
      (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  xt_rsc_0_12_i_da_d_pff <= modulo_add_28_qr_lpi_3_dfm_1;
  xt_rsc_0_13_i_adra_d_pff <= MUX1HOT_v_4_4_2((INNER_LOOP1_r_11_4_sva_6_0(3 DOWNTO
      0)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15604_itm_2, (INNER_LOOP3_r_11_4_sva_6_0(3
      DOWNTO 0)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15987_itm_2, STD_LOGIC_VECTOR'(
      (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  xt_rsc_0_13_i_da_d_pff <= modulo_add_29_qr_lpi_3_dfm_1;
  xt_rsc_0_14_i_adra_d_pff <= MUX1HOT_v_4_4_2((INNER_LOOP1_r_11_4_sva_6_0(3 DOWNTO
      0)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16115_itm_3, (INNER_LOOP3_r_11_4_sva_6_0(3
      DOWNTO 0)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16498_itm_3, STD_LOGIC_VECTOR'(
      (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  xt_rsc_0_14_i_da_d_pff <= modulo_add_30_qr_lpi_3_dfm_1;
  xt_rsc_0_15_i_adra_d_pff <= MUX1HOT_v_4_4_2((INNER_LOOP1_r_11_4_sva_6_0(3 DOWNTO
      0)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12027_itm_4, (INNER_LOOP3_r_11_4_sva_6_0(3
      DOWNTO 0)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12410_itm_4, STD_LOGIC_VECTOR'(
      (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  xt_rsc_0_15_i_da_d_pff <= modulo_add_31_qr_lpi_3_dfm_1;
  xt_rsc_0_16_i_wea_d_pff <= (and_dcpl_78 AND (fsm_output(9))) OR (and_dcpl_135 AND
      and_dcpl_79 AND (fsm_output(4)));
  xt_rsc_1_0_i_wea_d_pff <= (and_dcpl_82 AND (fsm_output(9))) OR (and_dcpl_135 AND
      and_dcpl_83 AND (fsm_output(4)));
  xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff <= (and_dcpl_145 AND butterFly2_f1_nor_cse
      AND (fsm_output(7))) OR (and_dcpl_147 AND butterFly1_f1_nor_cse AND (fsm_output(2)));
  xt_rsc_1_16_i_wea_d_pff <= (and_dcpl_89 AND (fsm_output(9))) OR (and_dcpl_135 AND
      and_8912_cse AND (fsm_output(4)));
  xt_rsc_2_0_i_wea_d_pff <= (and_dcpl_93 AND (fsm_output(9))) OR (and_dcpl_150 AND
      and_dcpl_69 AND (fsm_output(4)));
  xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff <= (and_dcpl_138 AND and_dcpl_152
      AND (fsm_output(7))) OR (and_dcpl_141 AND and_dcpl_154 AND (fsm_output(2)));
  xt_rsc_2_16_i_wea_d_pff <= (and_dcpl_96 AND (fsm_output(9))) OR (and_dcpl_150 AND
      and_dcpl_79 AND (fsm_output(4)));
  xt_rsc_3_0_i_wea_d_pff <= (and_dcpl_99 AND (fsm_output(9))) OR (and_dcpl_150 AND
      and_dcpl_83 AND (fsm_output(4)));
  xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff <= (and_dcpl_145 AND and_dcpl_152
      AND (fsm_output(7))) OR (and_dcpl_147 AND and_dcpl_154 AND (fsm_output(2)));
  xt_rsc_3_16_i_wea_d_pff <= (nor_tmp_22 AND (fsm_output(9))) OR (and_dcpl_150 AND
      and_8912_cse AND (fsm_output(4)));
  xt_rsc_4_0_i_da_d_pff <= reg_modulo_sub_16_qr_lpi_3_dfm_1_ftd & reg_modulo_sub_16_qr_lpi_3_dfm_1_ftd_1;
  xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff <= (and_dcpl_138 AND and_dcpl_161
      AND (fsm_output(7))) OR (and_dcpl_141 AND and_dcpl_163 AND (fsm_output(2)));
  xt_rsc_4_1_i_adra_d_pff <= MUX1HOT_v_4_4_2((INNER_LOOP1_r_11_4_sva_6_0(3 DOWNTO
      0)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13432_itm_6, (INNER_LOOP3_r_11_4_sva_6_0(3
      DOWNTO 0)), INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9472_itm_9, STD_LOGIC_VECTOR'(
      (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  xt_rsc_4_1_i_da_d_pff <= reg_modulo_sub_17_qr_lpi_3_dfm_1_ftd & reg_modulo_sub_17_qr_lpi_3_dfm_1_ftd_1;
  xt_rsc_4_2_i_adra_d_pff <= MUX1HOT_v_4_4_2((INNER_LOOP1_r_11_4_sva_6_0(3 DOWNTO
      0)), INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9855_itm_9, (INNER_LOOP3_r_11_4_sva_6_0(3
      DOWNTO 0)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_10015_itm_9, STD_LOGIC_VECTOR'(
      (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  xt_rsc_4_2_i_da_d_pff <= reg_modulo_sub_18_qr_lpi_3_dfm_1_ftd & reg_modulo_sub_18_qr_lpi_3_dfm_1_ftd_1;
  xt_rsc_4_3_i_da_d_pff <= reg_modulo_sub_19_qr_lpi_3_dfm_1_ftd & reg_modulo_sub_19_qr_lpi_3_dfm_1_ftd_1;
  xt_rsc_4_4_i_da_d_pff <= reg_modulo_sub_20_qr_lpi_3_dfm_1_ftd & reg_modulo_sub_20_qr_lpi_3_dfm_1_ftd_1;
  xt_rsc_4_5_i_da_d_pff <= reg_modulo_sub_21_qr_lpi_3_dfm_1_ftd & reg_modulo_sub_21_qr_lpi_3_dfm_1_ftd_1;
  xt_rsc_4_6_i_da_d_pff <= reg_modulo_sub_22_qr_lpi_3_dfm_1_ftd & reg_modulo_sub_22_qr_lpi_3_dfm_1_ftd_1;
  xt_rsc_4_7_i_da_d_pff <= reg_modulo_sub_23_qr_lpi_3_dfm_1_ftd & reg_modulo_sub_23_qr_lpi_3_dfm_1_ftd_1;
  xt_rsc_4_8_i_da_d_pff <= reg_modulo_sub_24_qr_lpi_3_dfm_1_ftd & reg_modulo_sub_24_qr_lpi_3_dfm_1_ftd_1;
  xt_rsc_4_9_i_adra_d_pff <= MUX1HOT_v_4_4_2((INNER_LOOP1_r_11_4_sva_6_0(3 DOWNTO
      0)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13560_itm_7, (INNER_LOOP3_r_11_4_sva_6_0(3
      DOWNTO 0)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13943_itm_7, STD_LOGIC_VECTOR'(
      (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  xt_rsc_4_9_i_da_d_pff <= reg_modulo_sub_25_qr_lpi_3_dfm_1_ftd & reg_modulo_sub_25_qr_lpi_3_dfm_1_ftd_1;
  xt_rsc_4_10_i_adra_d_pff <= MUX1HOT_v_4_4_2((INNER_LOOP1_r_11_4_sva_6_0(3 DOWNTO
      0)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14071_itm_8, (INNER_LOOP3_r_11_4_sva_6_0(3
      DOWNTO 0)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14454_itm_8, STD_LOGIC_VECTOR'(
      (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  xt_rsc_4_10_i_da_d_pff <= reg_modulo_sub_26_qr_lpi_3_dfm_1_ftd & reg_modulo_sub_26_qr_lpi_3_dfm_1_ftd_1;
  xt_rsc_4_11_i_da_d_pff <= reg_modulo_sub_27_qr_lpi_3_dfm_1_ftd & reg_modulo_sub_27_qr_lpi_3_dfm_1_ftd_1;
  xt_rsc_4_12_i_da_d_pff <= reg_modulo_sub_28_qr_lpi_3_dfm_1_ftd & reg_modulo_sub_28_qr_lpi_3_dfm_1_ftd_1;
  xt_rsc_4_13_i_da_d_pff <= reg_modulo_sub_29_qr_lpi_3_dfm_1_ftd & reg_modulo_sub_29_qr_lpi_3_dfm_1_ftd_1;
  xt_rsc_4_14_i_da_d_pff <= reg_modulo_sub_30_qr_lpi_3_dfm_1_ftd & reg_modulo_sub_30_qr_lpi_3_dfm_1_ftd_1;
  xt_rsc_4_15_i_da_d_pff <= reg_modulo_sub_31_qr_lpi_3_dfm_1_ftd & reg_modulo_sub_31_qr_lpi_3_dfm_1_ftd_1;
  xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff <= (and_dcpl_145 AND and_dcpl_161
      AND (fsm_output(7))) OR (and_dcpl_147 AND and_dcpl_163 AND (fsm_output(2)));
  xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff <= (and_dcpl_138 AND and_dcpl_167
      AND (fsm_output(7))) OR (and_dcpl_141 AND and_dcpl_169 AND (fsm_output(2)));
  xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff <= (and_dcpl_145 AND and_dcpl_167
      AND (fsm_output(7))) OR (and_dcpl_147 AND and_dcpl_169 AND (fsm_output(2)));
  twiddle_rsc_0_0_i_adra_d <= '0' & INNER_LOOP1_tw_h_mux1h_4_rmff;
  twiddle_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' &
      and_6824_rmff);
  twiddle_rsc_0_1_i_adra_d <= '0' & butterFly2_1_tw_butterFly2_1_tw_mux_rmff;
  twiddle_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' &
      or_3498_rmff);
  twiddle_rsc_0_2_i_adra_d <= '0' & butterFly2_1_tw_butterFly2_1_tw_mux_rmff;
  twiddle_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' &
      or_3502_rmff);
  twiddle_rsc_0_3_i_adra_d <= '0' & butterFly2_1_tw_butterFly2_1_tw_mux_rmff;
  twiddle_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' &
      or_3506_rmff);
  twiddle_rsc_0_4_i_adra_d <= '0' & butterFly2_1_tw_butterFly2_1_tw_mux_rmff;
  twiddle_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' &
      or_3510_rmff);
  twiddle_rsc_0_5_i_adra_d <= '0' & butterFly2_1_tw_butterFly2_1_tw_mux_rmff;
  twiddle_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' &
      or_3514_rmff);
  twiddle_rsc_0_6_i_adra_d <= '0' & butterFly2_1_tw_butterFly2_1_tw_mux_rmff;
  twiddle_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' &
      or_3518_rmff);
  twiddle_rsc_0_7_i_adra_d <= '0' & butterFly2_1_tw_butterFly2_1_tw_mux_rmff;
  twiddle_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' &
      or_3522_rmff);
  twiddle_rsc_0_8_i_adra_d <= '0' & butterFly2_1_tw_butterFly2_1_tw_mux_rmff;
  twiddle_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' &
      and_6895_rmff);
  twiddle_rsc_0_9_i_adra_d <= '0' & butterFly2_1_tw_butterFly2_1_tw_mux_rmff;
  twiddle_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' &
      or_3498_rmff);
  twiddle_rsc_0_10_i_adra_d <= '0' & butterFly2_1_tw_butterFly2_1_tw_mux_rmff;
  twiddle_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' &
      or_3502_rmff);
  twiddle_rsc_0_11_i_adra_d <= '0' & butterFly2_1_tw_butterFly2_1_tw_mux_rmff;
  twiddle_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' &
      or_3506_rmff);
  twiddle_rsc_0_12_i_adra_d <= '0' & butterFly2_1_tw_butterFly2_1_tw_mux_rmff;
  twiddle_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' &
      or_3510_rmff);
  twiddle_rsc_0_13_i_adra_d <= '0' & butterFly2_1_tw_butterFly2_1_tw_mux_rmff;
  twiddle_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' &
      or_3514_rmff);
  twiddle_rsc_0_14_i_adra_d <= '0' & butterFly2_1_tw_butterFly2_1_tw_mux_rmff;
  twiddle_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' &
      or_3518_rmff);
  twiddle_rsc_0_15_i_adra_d <= '0' & butterFly2_1_tw_butterFly2_1_tw_mux_rmff;
  twiddle_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' &
      or_3522_rmff);
  twiddle_h_rsc_0_0_i_adra_d <= '0' & INNER_LOOP1_tw_h_mux1h_4_rmff;
  twiddle_h_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0'
      & and_6824_rmff);
  twiddle_h_rsc_0_1_i_adra_d <= '0' & butterFly2_1_tw_butterFly2_1_tw_mux_rmff;
  twiddle_h_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0'
      & or_3498_rmff);
  twiddle_h_rsc_0_2_i_adra_d <= '0' & butterFly2_1_tw_butterFly2_1_tw_mux_rmff;
  twiddle_h_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0'
      & or_3502_rmff);
  twiddle_h_rsc_0_3_i_adra_d <= '0' & butterFly2_1_tw_butterFly2_1_tw_mux_rmff;
  twiddle_h_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0'
      & or_3506_rmff);
  twiddle_h_rsc_0_4_i_adra_d <= '0' & butterFly2_1_tw_butterFly2_1_tw_mux_rmff;
  twiddle_h_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0'
      & or_3510_rmff);
  twiddle_h_rsc_0_5_i_adra_d <= '0' & butterFly2_1_tw_butterFly2_1_tw_mux_rmff;
  twiddle_h_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0'
      & or_3514_rmff);
  twiddle_h_rsc_0_6_i_adra_d <= '0' & butterFly2_1_tw_butterFly2_1_tw_mux_rmff;
  twiddle_h_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0'
      & or_3518_rmff);
  twiddle_h_rsc_0_7_i_adra_d <= '0' & butterFly2_1_tw_butterFly2_1_tw_mux_rmff;
  twiddle_h_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0'
      & or_3522_rmff);
  twiddle_h_rsc_0_8_i_adra_d <= '0' & butterFly2_1_tw_butterFly2_1_tw_mux_rmff;
  twiddle_h_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0'
      & and_6895_rmff);
  twiddle_h_rsc_0_9_i_adra_d <= '0' & butterFly2_1_tw_butterFly2_1_tw_mux_rmff;
  twiddle_h_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0'
      & or_3498_rmff);
  twiddle_h_rsc_0_10_i_adra_d <= '0' & butterFly2_1_tw_butterFly2_1_tw_mux_rmff;
  twiddle_h_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0'
      & or_3502_rmff);
  twiddle_h_rsc_0_11_i_adra_d <= '0' & butterFly2_1_tw_butterFly2_1_tw_mux_rmff;
  twiddle_h_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0'
      & or_3506_rmff);
  twiddle_h_rsc_0_12_i_adra_d <= '0' & butterFly2_1_tw_butterFly2_1_tw_mux_rmff;
  twiddle_h_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0'
      & or_3510_rmff);
  twiddle_h_rsc_0_13_i_adra_d <= '0' & butterFly2_1_tw_butterFly2_1_tw_mux_rmff;
  twiddle_h_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0'
      & or_3514_rmff);
  twiddle_h_rsc_0_14_i_adra_d <= '0' & butterFly2_1_tw_butterFly2_1_tw_mux_rmff;
  twiddle_h_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0'
      & or_3518_rmff);
  twiddle_h_rsc_0_15_i_adra_d <= '0' & butterFly2_1_tw_butterFly2_1_tw_mux_rmff;
  twiddle_h_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0'
      & or_3522_rmff);
  butterFly1_15_f1_mux_cse <= MUX_s_1_2_2(butterFly1_15_f1_equal_tmp_1, butterFly2_15_f1_equal_tmp_1,
      fsm_output(7));
  butterFly1_15_f1_mux_1_cse <= MUX_s_1_2_2(butterFly1_15_f1_equal_tmp_1_1, butterFly1_15_f1_equal_tmp_3_1,
      fsm_output(7));
  butterFly1_15_f1_mux_2_cse <= MUX_s_1_2_2(butterFly1_15_f1_equal_tmp_2_1, butterFly1_15_f1_equal_tmp_4_1,
      fsm_output(7));
  butterFly1_15_f1_mux_3_cse <= MUX_s_1_2_2(butterFly1_15_f1_equal_tmp_3_1, butterFly1_15_f1_equal_tmp_5_1,
      fsm_output(7));
  butterFly1_15_f1_mux_4_cse <= MUX_s_1_2_2(butterFly1_15_f1_equal_tmp_4_1, butterFly1_15_f1_equal_tmp_6_1,
      fsm_output(7));
  butterFly1_15_f1_mux_5_cse <= MUX_s_1_2_2(butterFly1_15_f1_equal_tmp_5_1, butterFly1_15_f1_equal_tmp_7_1,
      fsm_output(7));
  butterFly1_15_f1_mux_6_cse <= MUX_s_1_2_2(butterFly1_15_f1_equal_tmp_6_1, butterFly1_15_f1_equal_tmp_1,
      fsm_output(7));
  butterFly1_15_f1_mux_7_cse <= MUX_s_1_2_2(butterFly1_15_f1_equal_tmp_7_1, butterFly2_15_f1_equal_tmp_7_1,
      fsm_output(7));
  butterFly1_31_f1_mux_cse <= MUX_s_1_2_2(butterFly1_15_f1_equal_tmp_1, butterFly2_15_f1_equal_tmp_1,
      fsm_output(9));
  butterFly1_31_f1_mux_1_cse <= MUX_s_1_2_2(butterFly1_15_f1_equal_tmp_1_1, butterFly1_15_f1_equal_tmp_3_1,
      fsm_output(9));
  butterFly1_31_f1_mux_2_cse <= MUX_s_1_2_2(butterFly1_15_f1_equal_tmp_2_1, butterFly1_15_f1_equal_tmp_4_1,
      fsm_output(9));
  butterFly1_31_f1_mux_3_cse <= MUX_s_1_2_2(butterFly1_15_f1_equal_tmp_3_1, butterFly1_15_f1_equal_tmp_5_1,
      fsm_output(9));
  butterFly1_31_f1_mux_4_cse <= MUX_s_1_2_2(butterFly1_15_f1_equal_tmp_4_1, butterFly1_15_f1_equal_tmp_6_1,
      fsm_output(9));
  butterFly1_31_f1_mux_5_cse <= MUX_s_1_2_2(butterFly1_15_f1_equal_tmp_5_1, butterFly1_15_f1_equal_tmp_7_1,
      fsm_output(9));
  butterFly1_31_f1_mux_6_cse <= MUX_s_1_2_2(butterFly1_15_f1_equal_tmp_6_1, butterFly1_15_f1_equal_tmp_1,
      fsm_output(9));
  butterFly1_31_f1_mux_7_cse <= MUX_s_1_2_2(butterFly1_15_f1_equal_tmp_7_1, butterFly2_15_f1_equal_tmp_7_1,
      fsm_output(9));
  butterFly2_f1_mux_cse <= MUX_s_1_2_2(butterFly2_15_f1_equal_tmp_1, butterFly1_15_f1_equal_tmp_1,
      fsm_output(2));
  butterFly2_f1_mux_1_cse <= MUX_s_1_2_2(butterFly1_15_f1_equal_tmp_3_1, butterFly1_15_f1_equal_tmp_1_1,
      fsm_output(2));
  butterFly2_f1_mux_2_cse <= MUX_s_1_2_2(butterFly1_15_f1_equal_tmp_4_1, butterFly1_15_f1_equal_tmp_2_1,
      fsm_output(2));
  butterFly2_f1_mux_3_cse <= MUX_s_1_2_2(butterFly1_15_f1_equal_tmp_5_1, butterFly1_15_f1_equal_tmp_3_1,
      fsm_output(2));
  butterFly2_f1_mux_4_cse <= MUX_s_1_2_2(butterFly1_15_f1_equal_tmp_6_1, butterFly1_15_f1_equal_tmp_4_1,
      fsm_output(2));
  butterFly2_f1_mux_5_cse <= MUX_s_1_2_2(butterFly1_15_f1_equal_tmp_7_1, butterFly1_15_f1_equal_tmp_5_1,
      fsm_output(2));
  butterFly2_f1_mux_6_cse <= MUX_s_1_2_2(butterFly1_15_f1_equal_tmp_1, butterFly1_15_f1_equal_tmp_6_1,
      fsm_output(2));
  butterFly2_f1_mux_7_cse <= MUX_s_1_2_2(butterFly2_15_f1_equal_tmp_7_1, butterFly1_15_f1_equal_tmp_7_1,
      fsm_output(2));
  butterFly2_21_f1_mux_cse <= MUX_s_1_2_2(butterFly2_15_f1_equal_tmp_1, butterFly1_15_f1_equal_tmp_1,
      fsm_output(4));
  butterFly2_21_f1_mux_1_cse <= MUX_s_1_2_2(butterFly1_15_f1_equal_tmp_3_1, butterFly1_15_f1_equal_tmp_1_1,
      fsm_output(4));
  butterFly2_21_f1_mux_2_cse <= MUX_s_1_2_2(butterFly1_15_f1_equal_tmp_4_1, butterFly1_15_f1_equal_tmp_2_1,
      fsm_output(4));
  butterFly2_21_f1_mux_3_cse <= MUX_s_1_2_2(butterFly1_15_f1_equal_tmp_5_1, butterFly1_15_f1_equal_tmp_3_1,
      fsm_output(4));
  butterFly2_21_f1_mux_4_cse <= MUX_s_1_2_2(butterFly1_15_f1_equal_tmp_6_1, butterFly1_15_f1_equal_tmp_4_1,
      fsm_output(4));
  butterFly2_21_f1_mux_5_cse <= MUX_s_1_2_2(butterFly1_15_f1_equal_tmp_7_1, butterFly1_15_f1_equal_tmp_5_1,
      fsm_output(4));
  butterFly2_21_f1_mux_6_cse <= MUX_s_1_2_2(butterFly1_15_f1_equal_tmp_1, butterFly1_15_f1_equal_tmp_6_1,
      fsm_output(4));
  butterFly2_21_f1_mux_7_cse <= MUX_s_1_2_2(butterFly2_15_f1_equal_tmp_7_1, butterFly1_15_f1_equal_tmp_7_1,
      fsm_output(4));
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( or_4976_cse = '1' ) THEN
        p_sva <= p_rsci_idat;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        c_1_sva <= '0';
      ELSIF ( ((fsm_output(0)) OR (fsm_output(5)) OR (fsm_output(9))) = '1' ) THEN
        c_1_sva <= c_mux_nl AND (NOT (fsm_output(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_yt_rsc_0_0_cgo_cse <= '0';
        reg_yt_rsc_0_16_cgo_cse <= '0';
        reg_yt_rsc_1_0_cgo_cse <= '0';
        reg_yt_rsc_1_16_cgo_cse <= '0';
        reg_yt_rsc_2_0_cgo_cse <= '0';
        reg_yt_rsc_2_16_cgo_cse <= '0';
        reg_yt_rsc_3_0_cgo_cse <= '0';
        reg_yt_rsc_3_16_cgo_cse <= '0';
        reg_yt_rsc_4_0_cgo_cse <= '0';
        reg_yt_rsc_4_16_cgo_cse <= '0';
        reg_yt_rsc_5_0_cgo_cse <= '0';
        reg_yt_rsc_5_16_cgo_cse <= '0';
        reg_yt_rsc_6_0_cgo_cse <= '0';
        reg_yt_rsc_6_16_cgo_cse <= '0';
        reg_yt_rsc_7_0_cgo_cse <= '0';
        reg_yt_rsc_7_16_cgo_cse <= '0';
        reg_xt_rsc_triosy_7_31_obj_ld_cse <= '0';
        reg_ensig_cgo_cse <= '0';
        reg_ensig_cgo_17_cse <= '0';
        butterFly1_15_conc_2_itm_2_1 <= STD_LOGIC_VECTOR'( "00");
        butterFly1_15_conc_2_itm_9_0 <= '0';
        butterFly1_15_conc_2_itm_8_0 <= '0';
        butterFly1_15_f1_equal_tmp_1 <= '0';
        butterFly1_15_f1_equal_tmp_1_1 <= '0';
        butterFly1_15_f1_equal_tmp_2_1 <= '0';
        butterFly1_15_f1_equal_tmp_3_1 <= '0';
        butterFly1_15_f1_equal_tmp_4_1 <= '0';
        butterFly1_15_f1_equal_tmp_5_1 <= '0';
        butterFly1_15_f1_equal_tmp_6_1 <= '0';
        butterFly1_15_f1_equal_tmp_7_1 <= '0';
        INNER_LOOP1_stage_0 <= '0';
        INNER_LOOP1_r_11_4_sva_6_0 <= STD_LOGIC_VECTOR'( "0000000");
        INNER_LOOP1_stage_0_2 <= '0';
        INNER_LOOP1_stage_0_3 <= '0';
        INNER_LOOP1_stage_0_10 <= '0';
        INNER_LOOP1_stage_0_11 <= '0';
        butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm <= STD_LOGIC_VECTOR'( "000");
        butterFly1_15_conc_2_itm_7_0 <= '0';
        butterFly1_15_conc_2_itm_6_0 <= '0';
        butterFly1_15_conc_2_itm_5_0 <= '0';
        butterFly1_15_conc_2_itm_4_2_1 <= STD_LOGIC_VECTOR'( "00");
        butterFly1_15_conc_2_itm_4_0 <= '0';
        butterFly1_15_conc_2_itm_3_0 <= '0';
        butterFly1_15_conc_2_itm_2_2_1 <= STD_LOGIC_VECTOR'( "00");
        butterFly1_15_conc_2_itm_2_0 <= '0';
        butterFly1_15_conc_2_itm_1_0 <= '0';
        butterFly1_15_conc_2_itm_0 <= '0';
        butterFly2_15_conc_2_itm_0 <= '0';
        butterFly2_15_conc_2_itm_1_0 <= '0';
        butterFly2_15_conc_2_itm_2_0 <= '0';
        butterFly2_15_conc_2_itm_3_0 <= '0';
        butterFly2_15_conc_2_itm_4_0 <= '0';
        butterFly2_15_conc_2_itm_5_0 <= '0';
        INNER_LOOP2_stage_0_10 <= '0';
        butterFly2_15_conc_2_itm_7_0 <= '0';
        butterFly2_15_conc_2_itm_8_0 <= '0';
        butterFly2_15_conc_itm_10_2_1 <= STD_LOGIC_VECTOR'( "00");
        butterFly2_15_f1_equal_tmp_1 <= '0';
        butterFly2_15_f1_equal_tmp_7_1 <= '0';
        INNER_LOOP3_r_11_4_sva_6_0 <= STD_LOGIC_VECTOR'( "0000000");
        INNER_LOOP4_r_11_4_sva_6_0 <= STD_LOGIC_VECTOR'( "0000000");
      ELSE
        reg_yt_rsc_0_0_cgo_cse <= or_553_rmff;
        reg_yt_rsc_0_16_cgo_cse <= or_652_rmff;
        reg_yt_rsc_1_0_cgo_cse <= or_718_rmff;
        reg_yt_rsc_1_16_cgo_cse <= or_785_rmff;
        reg_yt_rsc_2_0_cgo_cse <= or_851_rmff;
        reg_yt_rsc_2_16_cgo_cse <= or_918_rmff;
        reg_yt_rsc_3_0_cgo_cse <= or_984_rmff;
        reg_yt_rsc_3_16_cgo_cse <= or_1051_rmff;
        reg_yt_rsc_4_0_cgo_cse <= or_1117_rmff;
        reg_yt_rsc_4_16_cgo_cse <= or_1216_rmff;
        reg_yt_rsc_5_0_cgo_cse <= or_1282_rmff;
        reg_yt_rsc_5_16_cgo_cse <= or_1349_rmff;
        reg_yt_rsc_6_0_cgo_cse <= or_1415_rmff;
        reg_yt_rsc_6_16_cgo_cse <= or_1482_rmff;
        reg_yt_rsc_7_0_cgo_cse <= or_1548_rmff;
        reg_yt_rsc_7_16_cgo_cse <= or_1615_rmff;
        reg_xt_rsc_triosy_7_31_obj_ld_cse <= and_dcpl_62 AND (fsm_output(9));
        reg_ensig_cgo_cse <= or_3599_rmff;
        reg_ensig_cgo_17_cse <= or_3759_rmff;
        butterFly1_15_conc_2_itm_2_1 <= MUX_v_2_2_2(STAGE_LOOP_mux1h_nl, STD_LOGIC_VECTOR'("11"),
            or_4976_cse);
        butterFly1_15_conc_2_itm_9_0 <= butterFly1_15_conc_2_itm_8_0 AND (NOT or_tmp_3650);
        butterFly1_15_conc_2_itm_8_0 <= butterFly1_15_conc_2_itm_7_0 AND (NOT or_tmp_3650);
        butterFly1_15_f1_equal_tmp_1 <= MUX1HOT_s_1_4_2(butterFly1_f1_butterFly1_f1_nor_nl,
            butterFly1_16_f1_butterFly1_16_f1_nor_nl, butterFly2_f1_butterFly2_f1_and_5_nl,
            butterFly2_16_f1_butterFly2_16_f1_and_5_nl, STD_LOGIC_VECTOR'( (fsm_output(2))
            & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
        butterFly1_15_f1_equal_tmp_1_1 <= MUX1HOT_s_1_3_2(butterFly1_f1_butterFly1_f1_and_nl,
            butterFly1_16_f1_butterFly1_16_f1_and_nl, butterFly2_15_conc_2_itm_8_0,
            STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & or_dcpl_298));
        butterFly1_15_f1_equal_tmp_2_1 <= MUX1HOT_s_1_3_2(butterFly1_f1_butterFly1_f1_and_1_nl,
            butterFly1_16_f1_butterFly1_16_f1_and_1_nl, butterFly1_15_f1_equal_tmp_1_1,
            STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7))));
        butterFly1_15_f1_equal_tmp_3_1 <= MUX1HOT_s_1_4_2(butterFly1_f1_butterFly1_f1_and_2_nl,
            butterFly1_16_f1_butterFly1_16_f1_and_2_nl, butterFly2_f1_butterFly2_f1_and_nl,
            butterFly2_16_f1_butterFly2_16_f1_and_nl, STD_LOGIC_VECTOR'( (fsm_output(2))
            & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
        butterFly1_15_f1_equal_tmp_4_1 <= MUX1HOT_s_1_4_2(butterFly1_f1_butterFly1_f1_and_3_nl,
            butterFly1_16_f1_butterFly1_16_f1_and_3_nl, butterFly2_f1_butterFly2_f1_and_1_nl,
            butterFly2_16_f1_butterFly2_16_f1_and_1_nl, STD_LOGIC_VECTOR'( (fsm_output(2))
            & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
        butterFly1_15_f1_equal_tmp_5_1 <= MUX1HOT_s_1_4_2(butterFly1_f1_butterFly1_f1_and_4_nl,
            butterFly1_16_f1_butterFly1_16_f1_and_4_nl, butterFly2_f1_butterFly2_f1_and_2_nl,
            butterFly2_16_f1_butterFly2_16_f1_and_2_nl, STD_LOGIC_VECTOR'( (fsm_output(2))
            & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
        butterFly1_15_f1_equal_tmp_6_1 <= MUX1HOT_s_1_4_2(butterFly1_f1_butterFly1_f1_and_5_nl,
            butterFly1_16_f1_butterFly1_16_f1_and_5_nl, butterFly2_f1_butterFly2_f1_and_3_nl,
            butterFly2_16_f1_butterFly2_16_f1_and_3_nl, STD_LOGIC_VECTOR'( (fsm_output(2))
            & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
        butterFly1_15_f1_equal_tmp_7_1 <= MUX1HOT_s_1_4_2(butterFly1_f1_butterFly1_f1_and_6_nl,
            butterFly1_16_f1_butterFly1_16_f1_and_6_nl, butterFly2_f1_butterFly2_f1_and_4_nl,
            butterFly2_16_f1_butterFly2_16_f1_and_4_nl, STD_LOGIC_VECTOR'( (fsm_output(2))
            & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
        INNER_LOOP1_stage_0 <= (INNER_LOOP1_stage_0 AND (NOT (z_out_62(7)))) OR or_tmp_3650;
        INNER_LOOP1_r_11_4_sva_6_0 <= INNER_LOOP1_r_INNER_LOOP1_r_and_cse;
        INNER_LOOP1_stage_0_2 <= INNER_LOOP1_mux_nl AND (NOT or_tmp_3717);
        INNER_LOOP1_stage_0_3 <= INNER_LOOP1_mux_4_nl AND (NOT or_tmp_3717);
        INNER_LOOP1_stage_0_10 <= INNER_LOOP1_mux_5_nl AND (NOT or_tmp_3723);
        INNER_LOOP1_stage_0_11 <= INNER_LOOP1_mux_6_nl AND (NOT or_tmp_3723);
        butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm <= MUX1HOT_v_3_4_2((INNER_LOOP1_r_INNER_LOOP1_r_and_cse(6
            DOWNTO 4)), (INNER_LOOP2_r_11_4_sva_6_0_mx1(6 DOWNTO 4)), (INNER_LOOP1_r_INNER_LOOP1_r_and_3_cse(6
            DOWNTO 4)), (INNER_LOOP1_r_INNER_LOOP1_r_and_5_cse(6 DOWNTO 4)), STD_LOGIC_VECTOR'(
            or_tmp_3597 & or_dcpl_315 & or_tmp_3600 & or_tmp_3732));
        butterFly1_15_conc_2_itm_7_0 <= butterFly1_15_conc_2_itm_6_0 AND (NOT or_tmp_3650);
        butterFly1_15_conc_2_itm_6_0 <= butterFly1_15_conc_2_itm_5_0 AND (NOT or_tmp_3650);
        butterFly1_15_conc_2_itm_5_0 <= butterFly1_15_conc_2_itm_4_0 AND (NOT or_tmp_3650);
        butterFly1_15_conc_2_itm_4_2_1 <= MUX1HOT_v_2_3_2(butterFly1_15_conc_2_itm_3_2_1,
            (INNER_LOOP1_r_INNER_LOOP1_r_and_3_cse(6 DOWNTO 5)), (INNER_LOOP1_r_INNER_LOOP1_r_and_5_cse(6
            DOWNTO 5)), STD_LOGIC_VECTOR'( modulo_add_1_qelse_or_m1c & or_tmp_3600
            & or_tmp_3732));
        butterFly1_15_conc_2_itm_4_0 <= butterFly1_15_conc_2_itm_3_0 AND (NOT or_tmp_3650);
        butterFly1_15_conc_2_itm_3_0 <= butterFly1_15_conc_2_itm_2_0 AND (NOT or_tmp_3650);
        butterFly1_15_conc_2_itm_2_2_1 <= MUX1HOT_v_2_4_2(butterFly1_15_conc_2_itm_1_2_1,
            (operator_33_true_2_lshift_psp_2_0_sva_mx0(2 DOWNTO 1)), operator_33_true_3_lshift_psp_1_0_sva_mx0w5,
            operator_33_true_3_lshift_psp_1_0_sva, STD_LOGIC_VECTOR'( modulo_add_1_qelse_or_m1c
            & or_tmp_3600 & (fsm_output(8)) & (fsm_output(9))));
        butterFly1_15_conc_2_itm_2_0 <= butterFly1_15_mux_9_nl AND (NOT or_tmp_3650);
        butterFly1_15_conc_2_itm_1_0 <= butterFly1_15_conc_2_itm_0 AND (NOT(and_dcpl_239
            AND (NOT (fsm_output(7)))));
        butterFly1_15_conc_2_itm_0 <= butterFly1_15_mux1h_47_nl AND (NOT(or_4976_cse
            OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(8))));
        butterFly2_15_conc_2_itm_0 <= butterFly2_15_mux1h_3_nl AND (NOT((fsm_output(3))
            OR (fsm_output(10)) OR (fsm_output(0)) OR (fsm_output(1)) OR (fsm_output(5))));
        butterFly2_15_conc_2_itm_1_0 <= butterFly2_15_conc_2_itm_0 AND or_dcpl_300;
        butterFly2_15_conc_2_itm_2_0 <= butterFly2_15_conc_2_itm_1_0 AND or_dcpl_300;
        butterFly2_15_conc_2_itm_3_0 <= butterFly2_15_conc_2_itm_2_0 AND or_dcpl_300;
        butterFly2_15_conc_2_itm_4_0 <= butterFly2_15_conc_2_itm_3_0 AND or_dcpl_300;
        butterFly2_15_conc_2_itm_5_0 <= butterFly2_15_conc_2_itm_4_0 AND or_dcpl_300;
        INNER_LOOP2_stage_0_10 <= butterFly1_15_mux_10_nl AND (NOT or_tmp_3650);
        butterFly2_15_conc_2_itm_7_0 <= INNER_LOOP1_mux_7_nl AND ((fsm_output(4))
            OR (fsm_output(7)) OR (fsm_output(9)));
        butterFly2_15_conc_2_itm_8_0 <= butterFly2_15_conc_2_itm_7_0 AND or_tmp_3842;
        butterFly2_15_conc_itm_10_2_1 <= MUX1HOT_v_2_3_2(butterFly2_15_conc_2_itm_9_2_1,
            operator_33_true_3_lshift_psp_1_0_sva_mx0w5, operator_33_true_3_lshift_psp_1_0_sva,
            STD_LOGIC_VECTOR'( (fsm_output(7)) & (fsm_output(8)) & (fsm_output(9))));
        butterFly2_15_f1_equal_tmp_1 <= MUX_s_1_2_2(butterFly2_f1_butterFly2_f1_nor_nl,
            butterFly2_16_f1_butterFly2_16_f1_nor_nl, fsm_output(9));
        butterFly2_15_f1_equal_tmp_7_1 <= MUX_s_1_2_2(butterFly2_f1_butterFly2_f1_and_6_nl,
            butterFly2_16_f1_butterFly2_16_f1_and_6_cse, fsm_output(9));
        INNER_LOOP3_r_11_4_sva_6_0 <= INNER_LOOP1_r_INNER_LOOP1_r_and_3_cse;
        INNER_LOOP4_r_11_4_sva_6_0 <= INNER_LOOP1_r_INNER_LOOP1_r_and_5_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_8450_itm_9 <= MUX_v_4_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12027_itm_8,
          (INNER_LOOP3_r_11_4_sva_6_0(4 DOWNTO 1)), fsm_output(7));
      modulo_add_1_qr_lpi_3_dfm_1 <= MUX1HOT_v_32_4_2(z_out_141, (acc_2_nl(32 DOWNTO
          1)), z_out_138, z_out_136, STD_LOGIC_VECTOR'( modulo_add_1_qelse_and_nl
          & modulo_add_1_qelse_or_1_nl & modulo_add_1_qelse_and_4_nl & modulo_add_1_qelse_and_5_nl));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_8961_itm_9 <= MUX_v_4_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12538_itm_8,
          (INNER_LOOP3_r_11_4_sva_6_0(4 DOWNTO 1)), fsm_output(7));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_9472_itm_9 <= MUX_v_4_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13049_itm_8,
          (INNER_LOOP3_r_11_4_sva_6_0(4 DOWNTO 1)), fsm_output(7));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_10015_itm_9 <= MUX_v_4_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14582_itm_8,
          (INNER_LOOP3_r_11_4_sva_6_0(4 DOWNTO 1)), fsm_output(7));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_10494_itm_9 <= MUX_v_4_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15093_itm_8,
          (INNER_LOOP3_r_11_4_sva_6_0(4 DOWNTO 1)), fsm_output(7));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_11005_itm_9 <= MUX_v_4_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15604_itm_8,
          (INNER_LOOP3_r_11_4_sva_6_0(4 DOWNTO 1)), fsm_output(7));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_11516_itm_9 <= MUX_v_4_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16115_itm_8,
          (INNER_LOOP3_r_11_4_sva_6_0(4 DOWNTO 1)), fsm_output(7));
      modulo_add_10_qr_lpi_3_dfm_1 <= MUX1HOT_v_32_5_2(z_out_132, (acc_3_nl(32 DOWNTO
          1)), z_out_127, z_out_128, z_out_142, STD_LOGIC_VECTOR'( modulo_add_10_qelse_and_nl
          & modulo_add_10_qelse_or_nl & modulo_add_10_qelse_and_5_nl & modulo_add_10_qelse_and_6_nl
          & modulo_add_10_qelse_and_7_nl));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13560_itm_9 <= MUX_v_4_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13560_itm_8,
          (INNER_LOOP3_r_11_4_sva_6_0(4 DOWNTO 1)), fsm_output(7));
      modulo_add_11_qr_lpi_3_dfm_1 <= MUX1HOT_v_32_5_2(z_out_131, (acc_4_nl(32 DOWNTO
          1)), z_out_137, z_out_127, z_out_141, STD_LOGIC_VECTOR'( modulo_add_11_qelse_and_nl
          & modulo_add_11_qelse_or_nl & modulo_add_11_qelse_and_5_nl & modulo_add_11_qelse_and_6_nl
          & modulo_add_11_qelse_and_7_nl));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14071_itm_9 <= MUX1HOT_v_4_4_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14071_itm_8,
          (INNER_LOOP2_r_11_4_sva_6_0(4 DOWNTO 1)), (INNER_LOOP3_r_11_4_sva_6_0(4
          DOWNTO 1)), (INNER_LOOP4_r_11_4_sva_6_0(4 DOWNTO 1)), STD_LOGIC_VECTOR'(
          (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
      modulo_add_12_qr_lpi_3_dfm_1 <= MUX1HOT_v_32_4_2(z_out_130, (acc_5_nl(32 DOWNTO
          1)), z_out_142, z_out_140, STD_LOGIC_VECTOR'( modulo_add_12_qelse_and_nl
          & modulo_add_12_qelse_or_1_nl & modulo_add_12_qelse_and_4_nl & modulo_add_12_qelse_and_5_nl));
      modulo_add_13_qr_lpi_3_dfm_1 <= MUX1HOT_v_32_4_2(z_out_129, (acc_6_nl(32 DOWNTO
          1)), z_out_141, z_out_139, STD_LOGIC_VECTOR'( modulo_add_13_qelse_and_nl
          & modulo_add_13_qelse_or_1_nl & modulo_add_13_qelse_and_4_nl & modulo_add_13_qelse_and_5_nl));
      modulo_add_14_qr_lpi_3_dfm_1 <= MUX1HOT_v_32_4_2(z_out_128, (acc_10_nl(32 DOWNTO
          1)), z_out_140, z_out_138, STD_LOGIC_VECTOR'( modulo_add_14_qelse_and_nl
          & modulo_add_14_qelse_or_1_nl & modulo_add_14_qelse_and_4_nl & modulo_add_14_qelse_and_5_nl));
      modulo_add_15_qr_lpi_3_dfm_1 <= MUX1HOT_v_32_5_2(z_out_127, (acc_14_nl(32 DOWNTO
          1)), z_out_142, z_out_139, z_out_137, STD_LOGIC_VECTOR'( modulo_add_15_qelse_and_nl
          & modulo_add_15_qelse_or_nl & modulo_add_15_qelse_and_5_nl & modulo_add_15_qelse_and_6_nl
          & modulo_add_15_qelse_and_7_nl));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13943_itm_8 <= MUX1HOT_v_4_3_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13943_itm_7,
          (INNER_LOOP2_r_11_4_sva_6_0(4 DOWNTO 1)), (INNER_LOOP4_r_11_4_sva_6_0(4
          DOWNTO 1)), STD_LOGIC_VECTOR'( or_dcpl_353 & (fsm_output(4)) & (fsm_output(9))));
      mult_15_z_asn_itm_3 <= MUX1HOT_v_32_4_2(mult_15_z_asn_itm_2, mult_31_z_asn_itm_2,
          mult_14_z_asn_itm_2, mult_27_z_asn_itm_2, STD_LOGIC_VECTOR'( (fsm_output(2))
          & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
      mult_14_z_asn_itm_3 <= MUX1HOT_v_32_4_2(mult_14_z_asn_itm_2, mult_30_z_asn_itm_2,
          mult_26_z_asn_itm_2, mult_15_z_asn_itm_2, STD_LOGIC_VECTOR'( (fsm_output(2))
          & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
      mult_13_z_asn_itm_3 <= MUX1HOT_v_32_3_2(mult_13_z_asn_itm_2, mult_29_z_asn_itm_2,
          mult_28_z_asn_itm_2, STD_LOGIC_VECTOR'( or_dcpl_353 & (fsm_output(4)) &
          (fsm_output(9))));
      mult_12_z_asn_itm_3 <= MUX1HOT_v_32_3_2(mult_12_z_asn_itm_2, mult_28_z_asn_itm_2,
          mult_29_z_asn_itm_2, STD_LOGIC_VECTOR'( or_tmp_3666 & (fsm_output(4)) &
          (fsm_output(7))));
      mult_11_z_asn_itm_3 <= MUX1HOT_v_32_4_2(mult_11_z_asn_itm_2, mult_27_z_asn_itm_2,
          mult_15_z_asn_itm_2, mult_26_z_asn_itm_2, STD_LOGIC_VECTOR'( (fsm_output(2))
          & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
      mult_10_z_asn_itm_3 <= MUX1HOT_v_32_4_2(mult_10_z_asn_itm_2, mult_26_z_asn_itm_2,
          mult_25_z_asn_itm_2, mult_1_z_asn_itm_2, STD_LOGIC_VECTOR'( (fsm_output(2))
          & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13560_itm_8 <= MUX1HOT_v_4_3_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13560_itm_7,
          (INNER_LOOP2_r_11_4_sva_6_0(4 DOWNTO 1)), (INNER_LOOP4_r_11_4_sva_6_0(4
          DOWNTO 1)), STD_LOGIC_VECTOR'( or_dcpl_353 & (fsm_output(4)) & (fsm_output(9))));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13432_itm_7 <= MUX1HOT_v_4_3_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13432_itm_6,
          (INNER_LOOP2_r_11_4_sva_6_0(4 DOWNTO 1)), (INNER_LOOP4_r_11_4_sva_6_0(4
          DOWNTO 1)), STD_LOGIC_VECTOR'( or_dcpl_353 & (fsm_output(4)) & (fsm_output(9))));
      mult_15_z_asn_itm_1 <= MUX1HOT_v_32_3_2(mult_z_mul_cmp_2_z, mult_z_mul_cmp_22_z,
          mult_z_mul_cmp_20_z, STD_LOGIC_VECTOR'( (fsm_output(2)) & or_dcpl_361 &
          (fsm_output(9))));
      mult_14_z_asn_itm_1 <= MUX1HOT_v_32_3_2(mult_z_mul_cmp_4_z, mult_z_mul_cmp_24_z,
          mult_z_mul_cmp_28_z, STD_LOGIC_VECTOR'( or_tmp_3666 & (fsm_output(4)) &
          (fsm_output(7))));
      mult_13_z_asn_itm_1 <= MUX1HOT_v_32_4_2(mult_z_mul_cmp_6_z, mult_z_mul_cmp_26_z,
          mult_z_mul_cmp_24_z, mult_z_mul_cmp_12_z, STD_LOGIC_VECTOR'( (fsm_output(2))
          & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
      mult_12_z_asn_itm_1 <= MUX1HOT_v_32_3_2(mult_z_mul_cmp_8_z, mult_z_mul_cmp_28_z,
          mult_z_mul_cmp_12_z, STD_LOGIC_VECTOR'( (fsm_output(2)) & or_tmp_3755 &
          (fsm_output(7))));
      mult_11_z_asn_itm_1 <= MUX1HOT_v_32_4_2(mult_z_mul_cmp_10_z, mult_z_mul_cmp_30_z,
          mult_z_mul_cmp_8_z, mult_z_mul_cmp_16_z, STD_LOGIC_VECTOR'( (fsm_output(2))
          & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
      mult_10_z_asn_itm_1 <= MUX1HOT_v_32_3_2(mult_z_mul_cmp_12_z, mult_z_mul_cmp_z,
          mult_z_mul_cmp_2_z, STD_LOGIC_VECTOR'( (fsm_output(2)) & or_tmp_3755 &
          (fsm_output(7))));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13049_itm_7 <= MUX1HOT_v_4_3_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13049_itm_6,
          (INNER_LOOP2_r_11_4_sva_6_0(4 DOWNTO 1)), (INNER_LOOP4_r_11_4_sva_6_0(4
          DOWNTO 1)), STD_LOGIC_VECTOR'( or_dcpl_353 & (fsm_output(4)) & (fsm_output(9))));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12921_itm_6 <= MUX1HOT_v_4_3_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12921_itm_5,
          (INNER_LOOP2_r_11_4_sva_6_0(4 DOWNTO 1)), (INNER_LOOP4_r_11_4_sva_6_0(4
          DOWNTO 1)), STD_LOGIC_VECTOR'( or_dcpl_353 & (fsm_output(4)) & (fsm_output(9))));
      mult_1_z_asn_itm_1 <= MUX1HOT_v_32_4_2(mult_z_mul_cmp_30_z, mult_z_mul_cmp_20_z,
          mult_z_mul_cmp_16_z, mult_z_mul_cmp_26_z, STD_LOGIC_VECTOR'( (fsm_output(2))
          & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12538_itm_6 <= MUX1HOT_v_4_3_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12538_itm_5,
          (INNER_LOOP2_r_11_4_sva_6_0(4 DOWNTO 1)), (INNER_LOOP4_r_11_4_sva_6_0(4
          DOWNTO 1)), STD_LOGIC_VECTOR'( or_dcpl_353 & (fsm_output(4)) & (fsm_output(9))));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12410_itm_5 <= MUX1HOT_v_4_3_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12410_itm_4,
          (INNER_LOOP2_r_11_4_sva_6_0(4 DOWNTO 1)), (INNER_LOOP4_r_11_4_sva_6_0(4
          DOWNTO 1)), STD_LOGIC_VECTOR'( or_dcpl_353 & (fsm_output(4)) & (fsm_output(9))));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16498_itm_4 <= MUX1HOT_v_4_3_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16498_itm_3,
          (INNER_LOOP2_r_11_4_sva_6_0(4 DOWNTO 1)), (INNER_LOOP4_r_11_4_sva_6_0(4
          DOWNTO 1)), STD_LOGIC_VECTOR'( or_dcpl_353 & (fsm_output(4)) & (fsm_output(9))));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12027_itm_5 <= MUX1HOT_v_4_3_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12027_itm_4,
          (INNER_LOOP2_r_11_4_sva_6_0(4 DOWNTO 1)), (INNER_LOOP4_r_11_4_sva_6_0(4
          DOWNTO 1)), STD_LOGIC_VECTOR'( or_dcpl_353 & (fsm_output(4)) & (fsm_output(9))));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16115_itm_4 <= MUX1HOT_v_4_3_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16115_itm_3,
          (INNER_LOOP2_r_11_4_sva_6_0(4 DOWNTO 1)), (INNER_LOOP4_r_11_4_sva_6_0(4
          DOWNTO 1)), STD_LOGIC_VECTOR'( or_dcpl_353 & (fsm_output(4)) & (fsm_output(9))));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15987_itm_3 <= MUX1HOT_v_4_3_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15987_itm_2,
          (INNER_LOOP2_r_11_4_sva_6_0(4 DOWNTO 1)), (INNER_LOOP4_r_11_4_sva_6_0(4
          DOWNTO 1)), STD_LOGIC_VECTOR'( or_dcpl_353 & (fsm_output(4)) & (fsm_output(9))));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15604_itm_3 <= MUX1HOT_v_4_3_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15604_itm_2,
          (INNER_LOOP2_r_11_4_sva_6_0(4 DOWNTO 1)), (INNER_LOOP4_r_11_4_sva_6_0(4
          DOWNTO 1)), STD_LOGIC_VECTOR'( or_dcpl_353 & (fsm_output(4)) & (fsm_output(9))));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15476_itm_2 <= MUX1HOT_v_4_3_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15476_itm_1,
          (INNER_LOOP2_r_11_4_sva_6_0(4 DOWNTO 1)), (INNER_LOOP4_r_11_4_sva_6_0(4
          DOWNTO 1)), STD_LOGIC_VECTOR'( or_dcpl_353 & (fsm_output(4)) & (fsm_output(9))));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16498_itm_1 <= MUX_v_4_2_2((INNER_LOOP1_r_11_4_sva_6_0(4
          DOWNTO 1)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_11516_itm_9, or_tmp_3842);
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15987_itm_1 <= MUX_v_4_2_2((INNER_LOOP1_r_11_4_sva_6_0(4
          DOWNTO 1)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_11005_itm_9, or_tmp_3842);
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15476_itm_1 <= MUX_v_4_2_2((INNER_LOOP1_r_11_4_sva_6_0(4
          DOWNTO 1)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_10494_itm_9, or_tmp_3842);
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15093_itm_2 <= MUX1HOT_v_4_3_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15093_itm_1,
          (INNER_LOOP2_r_11_4_sva_6_0(4 DOWNTO 1)), (INNER_LOOP4_r_11_4_sva_6_0(4
          DOWNTO 1)), STD_LOGIC_VECTOR'( or_dcpl_353 & (fsm_output(4)) & (fsm_output(9))));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14965_itm_1 <= MUX1HOT_v_4_4_2((INNER_LOOP1_r_11_4_sva_6_0(4
          DOWNTO 1)), (INNER_LOOP2_r_11_4_sva_6_0(4 DOWNTO 1)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_10015_itm_9,
          (INNER_LOOP4_r_11_4_sva_6_0(4 DOWNTO 1)), STD_LOGIC_VECTOR'( (fsm_output(2))
          & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14454_itm_1 <= MUX_v_4_2_2((INNER_LOOP1_r_11_4_sva_6_0(4
          DOWNTO 1)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14071_itm_9, or_tmp_3842);
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13943_itm_1 <= MUX_v_4_2_2((INNER_LOOP1_r_11_4_sva_6_0(4
          DOWNTO 1)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13560_itm_9, or_tmp_3842);
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13432_itm_1 <= MUX_v_4_2_2((INNER_LOOP1_r_11_4_sva_6_0(4
          DOWNTO 1)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_9472_itm_9, or_tmp_3842);
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12921_itm_1 <= MUX_v_4_2_2((INNER_LOOP1_r_11_4_sva_6_0(4
          DOWNTO 1)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_8961_itm_9, or_tmp_3842);
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12410_itm_1 <= MUX_v_4_2_2((INNER_LOOP1_r_11_4_sva_6_0(4
          DOWNTO 1)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_8450_itm_9, or_tmp_3842);
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16115_itm_1 <= MUX1HOT_v_4_3_2((INNER_LOOP1_r_11_4_sva_6_0(4
          DOWNTO 1)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_11388_itm_8, (INNER_LOOP3_r_11_4_sva_6_0(4
          DOWNTO 1)), STD_LOGIC_VECTOR'( (fsm_output(2)) & or_tmp_3755 & (fsm_output(7))));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15604_itm_1 <= MUX1HOT_v_4_3_2((INNER_LOOP1_r_11_4_sva_6_0(4
          DOWNTO 1)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_10877_itm_8, (INNER_LOOP3_r_11_4_sva_6_0(4
          DOWNTO 1)), STD_LOGIC_VECTOR'( (fsm_output(2)) & or_tmp_3755 & (fsm_output(7))));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15093_itm_1 <= MUX1HOT_v_4_3_2((INNER_LOOP1_r_11_4_sva_6_0(4
          DOWNTO 1)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_10366_itm_8, (INNER_LOOP3_r_11_4_sva_6_0(4
          DOWNTO 1)), STD_LOGIC_VECTOR'( (fsm_output(2)) & or_tmp_3755 & (fsm_output(7))));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14582_itm_1 <= MUX1HOT_v_4_4_2((INNER_LOOP1_r_11_4_sva_6_0(4
          DOWNTO 1)), (INNER_LOOP2_r_11_4_sva_6_0(4 DOWNTO 1)), (INNER_LOOP3_r_11_4_sva_6_0(4
          DOWNTO 1)), (INNER_LOOP4_r_11_4_sva_6_0(4 DOWNTO 1)), STD_LOGIC_VECTOR'(
          (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14071_itm_1 <= MUX1HOT_v_4_3_2((INNER_LOOP1_r_11_4_sva_6_0(4
          DOWNTO 1)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13943_itm_8, (INNER_LOOP3_r_11_4_sva_6_0(4
          DOWNTO 1)), STD_LOGIC_VECTOR'( (fsm_output(2)) & or_tmp_3755 & (fsm_output(7))));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13560_itm_1 <= MUX1HOT_v_4_3_2((INNER_LOOP1_r_11_4_sva_6_0(4
          DOWNTO 1)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_9855_itm_8, (INNER_LOOP3_r_11_4_sva_6_0(4
          DOWNTO 1)), STD_LOGIC_VECTOR'( (fsm_output(2)) & or_tmp_3755 & (fsm_output(7))));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13049_itm_1 <= MUX1HOT_v_4_3_2((INNER_LOOP1_r_11_4_sva_6_0(4
          DOWNTO 1)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_9344_itm_8, (INNER_LOOP3_r_11_4_sva_6_0(4
          DOWNTO 1)), STD_LOGIC_VECTOR'( (fsm_output(2)) & or_tmp_3755 & (fsm_output(7))));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12538_itm_1 <= MUX1HOT_v_4_3_2((INNER_LOOP1_r_11_4_sva_6_0(4
          DOWNTO 1)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_8833_itm_8, (INNER_LOOP3_r_11_4_sva_6_0(4
          DOWNTO 1)), STD_LOGIC_VECTOR'( (fsm_output(2)) & or_tmp_3755 & (fsm_output(7))));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12027_itm_1 <= MUX1HOT_v_4_3_2((INNER_LOOP1_r_11_4_sva_6_0(4
          DOWNTO 1)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_11899_itm_8, (INNER_LOOP3_r_11_4_sva_6_0(4
          DOWNTO 1)), STD_LOGIC_VECTOR'( (fsm_output(2)) & or_tmp_3755 & (fsm_output(7))));
      mult_16_z_asn_itm_3 <= MUX_v_32_2_2(mult_31_z_asn_itm_2, mult_10_z_asn_itm_2,
          or_dcpl_361);
      mult_17_z_asn_itm_3 <= MUX1HOT_v_32_4_2(mult_1_z_asn_itm_2, mult_11_z_asn_itm_2,
          mult_31_z_asn_itm_2, mult_10_z_asn_itm_2, STD_LOGIC_VECTOR'( (fsm_output(2))
          & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
      mult_18_z_asn_itm_3 <= MUX1HOT_v_32_3_2(mult_23_z_asn_itm_2, mult_12_z_asn_itm_2,
          mult_24_z_asn_itm_2, STD_LOGIC_VECTOR'( or_tmp_3666 & (fsm_output(4)) &
          (fsm_output(7))));
      mult_19_z_asn_itm_3 <= MUX1HOT_v_32_3_2(mult_24_z_asn_itm_2, mult_13_z_asn_itm_2,
          mult_23_z_asn_itm_2, STD_LOGIC_VECTOR'( or_tmp_3666 & (fsm_output(4)) &
          (fsm_output(7))));
      mult_20_z_asn_itm_3 <= MUX1HOT_v_32_4_2(mult_25_z_asn_itm_2, mult_14_z_asn_itm_2,
          mult_28_z_asn_itm_2, mult_13_z_asn_itm_2, STD_LOGIC_VECTOR'( (fsm_output(2))
          & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
      mult_21_z_asn_itm_3 <= MUX1HOT_v_32_4_2(mult_26_z_asn_itm_2, mult_15_z_asn_itm_2,
          mult_11_z_asn_itm_2, mult_30_z_asn_itm_2, STD_LOGIC_VECTOR'( (fsm_output(2))
          & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
      mult_22_z_asn_itm_3 <= MUX1HOT_v_32_3_2(mult_27_z_asn_itm_2, mult_1_z_asn_itm_2,
          mult_14_z_asn_itm_2, STD_LOGIC_VECTOR'( or_dcpl_353 & (fsm_output(4)) &
          (fsm_output(9))));
      mult_23_z_asn_itm_3 <= MUX1HOT_v_32_4_2(mult_28_z_asn_itm_2, mult_23_z_asn_itm_2,
          mult_1_z_asn_itm_2, mult_25_z_asn_itm_2, STD_LOGIC_VECTOR'( (fsm_output(2))
          & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
      mult_24_z_asn_itm_3 <= MUX1HOT_v_32_3_2(mult_29_z_asn_itm_2, mult_24_z_asn_itm_2,
          mult_12_z_asn_itm_2, STD_LOGIC_VECTOR'( or_tmp_3666 & (fsm_output(4)) &
          (fsm_output(7))));
      mult_25_z_asn_itm_3 <= MUX1HOT_v_32_3_2(mult_30_z_asn_itm_2, mult_25_z_asn_itm_2,
          mult_11_z_asn_itm_2, STD_LOGIC_VECTOR'( or_dcpl_353 & (fsm_output(4)) &
          (fsm_output(9))));
      modulo_add_23_qr_lpi_3_dfm_1 <= MUX1HOT_v_32_4_2(z_out_140, (acc_18_nl(32 DOWNTO
          1)), z_out_137, z_out_135, STD_LOGIC_VECTOR'( modulo_add_23_qelse_and_nl
          & modulo_add_23_qelse_or_1_nl & modulo_add_23_qelse_and_4_nl & modulo_add_23_qelse_and_5_nl));
      modulo_add_24_qr_lpi_3_dfm_1 <= MUX1HOT_v_32_4_2(z_out_139, (acc_22_nl(32 DOWNTO
          1)), z_out_136, z_out_134, STD_LOGIC_VECTOR'( modulo_add_24_qelse_and_nl
          & modulo_add_24_qelse_or_1_nl & modulo_add_24_qelse_and_4_nl & modulo_add_24_qelse_and_5_nl));
      modulo_add_25_qr_lpi_3_dfm_1 <= MUX1HOT_v_32_4_2(z_out_138, (acc_26_nl(32 DOWNTO
          1)), z_out_135, z_out_133, STD_LOGIC_VECTOR'( modulo_add_25_qelse_and_nl
          & modulo_add_25_qelse_or_1_nl & modulo_add_25_qelse_and_4_nl & modulo_add_25_qelse_and_5_nl));
      modulo_add_26_qr_lpi_3_dfm_1 <= MUX1HOT_v_32_5_2(z_out_137, (acc_30_nl(32 DOWNTO
          1)), z_out_136, z_out_134, z_out_132, STD_LOGIC_VECTOR'( modulo_add_26_qelse_and_nl
          & modulo_add_26_qelse_or_nl & modulo_add_26_qelse_and_5_nl & modulo_add_26_qelse_and_6_nl
          & modulo_add_26_qelse_and_7_nl));
      modulo_add_27_qr_lpi_3_dfm_1 <= MUX1HOT_v_32_5_2(z_out_136, (acc_34_nl(32 DOWNTO
          1)), z_out_135, z_out_133, z_out_131, STD_LOGIC_VECTOR'( modulo_add_27_qelse_and_nl
          & modulo_add_27_qelse_or_nl & modulo_add_27_qelse_and_5_nl & modulo_add_27_qelse_and_6_nl
          & modulo_add_27_qelse_and_7_nl));
      modulo_add_28_qr_lpi_3_dfm_1 <= MUX1HOT_v_32_5_2(z_out_135, (acc_38_nl(32 DOWNTO
          1)), z_out_134, z_out_132, z_out_130, STD_LOGIC_VECTOR'( modulo_add_28_qelse_and_nl
          & modulo_add_28_qelse_or_nl & modulo_add_28_qelse_and_5_nl & modulo_add_28_qelse_and_6_nl
          & modulo_add_28_qelse_and_7_nl));
      modulo_add_29_qr_lpi_3_dfm_1 <= MUX1HOT_v_32_5_2(z_out_134, (acc_42_nl(32 DOWNTO
          1)), z_out_133, z_out_131, z_out_129, STD_LOGIC_VECTOR'( modulo_add_29_qelse_and_nl
          & modulo_add_29_qelse_or_nl & modulo_add_29_qelse_and_5_nl & modulo_add_29_qelse_and_6_nl
          & modulo_add_29_qelse_and_7_nl));
      modulo_add_30_qr_lpi_3_dfm_1 <= MUX1HOT_v_32_5_2(z_out_133, (acc_46_nl(32 DOWNTO
          1)), z_out_132, z_out_130, z_out_128, STD_LOGIC_VECTOR'( modulo_add_30_qelse_and_nl
          & modulo_add_30_qelse_or_nl & modulo_add_30_qelse_and_5_nl & modulo_add_30_qelse_and_6_nl
          & modulo_add_30_qelse_and_7_nl));
      modulo_add_31_qr_lpi_3_dfm_1 <= MUX1HOT_v_32_5_2(z_out_142, (acc_49_nl(32 DOWNTO
          1)), z_out_131, z_out_129, z_out_127, STD_LOGIC_VECTOR'( modulo_add_31_qelse_and_nl
          & modulo_add_31_qelse_or_nl & modulo_add_31_qelse_and_5_nl & modulo_add_31_qelse_and_6_nl
          & modulo_add_31_qelse_and_7_nl));
      mult_23_z_asn_itm_1 <= MUX1HOT_v_32_4_2(mult_z_mul_cmp_28_z, mult_z_mul_cmp_18_z,
          mult_z_mul_cmp_6_z, mult_z_mul_cmp_10_z, STD_LOGIC_VECTOR'( (fsm_output(2))
          & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
      mult_24_z_asn_itm_1 <= MUX1HOT_v_32_4_2(mult_z_mul_cmp_26_z, mult_z_mul_cmp_16_z,
          mult_z_mul_cmp_10_z, mult_z_mul_cmp_2_z, STD_LOGIC_VECTOR'( (fsm_output(2))
          & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
      mult_25_z_asn_itm_1 <= MUX1HOT_v_32_4_2(mult_z_mul_cmp_24_z, mult_z_mul_cmp_14_z,
          mult_z_mul_cmp_18_z, mult_z_mul_cmp_8_z, STD_LOGIC_VECTOR'( (fsm_output(2))
          & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
      mult_26_z_asn_itm_1 <= MUX1HOT_v_32_4_2(mult_z_mul_cmp_22_z, mult_z_mul_cmp_12_z,
          mult_z_mul_cmp_26_z, mult_z_mul_cmp_18_z, STD_LOGIC_VECTOR'( (fsm_output(2))
          & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
      mult_27_z_asn_itm_1 <= MUX1HOT_v_32_4_2(mult_z_mul_cmp_20_z, mult_z_mul_cmp_10_z,
          mult_z_mul_cmp_30_z, mult_z_mul_cmp_24_z, STD_LOGIC_VECTOR'( (fsm_output(2))
          & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
      mult_28_z_asn_itm_1 <= MUX1HOT_v_32_4_2(mult_z_mul_cmp_18_z, mult_z_mul_cmp_8_z,
          mult_z_mul_cmp_20_z, mult_z_mul_cmp_30_z, STD_LOGIC_VECTOR'( (fsm_output(2))
          & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
      mult_29_z_asn_itm_1 <= MUX1HOT_v_32_4_2(mult_z_mul_cmp_16_z, mult_z_mul_cmp_6_z,
          mult_z_mul_cmp_14_z, mult_z_mul_cmp_22_z, STD_LOGIC_VECTOR'( (fsm_output(2))
          & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
      mult_30_z_asn_itm_1 <= MUX_v_32_2_2(mult_z_mul_cmp_14_z, mult_z_mul_cmp_4_z,
          or_dcpl_361);
      mult_31_z_asn_itm_1 <= MUX1HOT_v_32_3_2(mult_z_mul_cmp_z, mult_z_mul_cmp_2_z,
          mult_z_mul_cmp_6_z, STD_LOGIC_VECTOR'( or_dcpl_353 & (fsm_output(4)) &
          (fsm_output(9))));
      tmp_10_lpi_3_dfm_2 <= MUX1HOT_v_32_4_2(tmp_64_lpi_3_dfm_1, tmp_10_lpi_3_dfm_1,
          tmp_100_lpi_3_dfm_1, tmp_32_lpi_3_dfm_1, STD_LOGIC_VECTOR'( (fsm_output(2))
          & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
      tmp_102_lpi_3_dfm_2 <= MUX1HOT_v_32_4_2(tmp_66_lpi_3_dfm_1, tmp_12_lpi_3_dfm_1,
          tmp_102_lpi_3_dfm_1, tmp_34_lpi_3_dfm_1, STD_LOGIC_VECTOR'( (fsm_output(2))
          & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
      tmp_104_lpi_3_dfm_2 <= MUX1HOT_v_32_4_2(tmp_68_lpi_3_dfm_1, tmp_14_lpi_3_dfm_1,
          tmp_104_lpi_3_dfm_1, tmp_36_lpi_3_dfm_1, STD_LOGIC_VECTOR'( (fsm_output(2))
          & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
      tmp_106_lpi_3_dfm_2 <= MUX1HOT_v_32_4_2(tmp_70_lpi_3_dfm_1, tmp_16_lpi_3_dfm_1,
          tmp_106_lpi_3_dfm_1, tmp_38_lpi_3_dfm_1, STD_LOGIC_VECTOR'( (fsm_output(2))
          & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
      tmp_108_lpi_3_dfm_2 <= MUX1HOT_v_32_4_2(tmp_72_lpi_3_dfm_1, tmp_18_lpi_3_dfm_1,
          tmp_108_lpi_3_dfm_1, tmp_40_lpi_3_dfm_1, STD_LOGIC_VECTOR'( (fsm_output(2))
          & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
      tmp_110_lpi_3_dfm_2 <= MUX1HOT_v_32_4_2(tmp_74_lpi_3_dfm_1, tmp_2_lpi_3_dfm_1,
          tmp_110_lpi_3_dfm_1, tmp_42_lpi_3_dfm_1, STD_LOGIC_VECTOR'( (fsm_output(2))
          & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
      tmp_112_lpi_3_dfm_2 <= MUX1HOT_v_32_4_2(tmp_76_lpi_3_dfm_1, tmp_20_lpi_3_dfm_1,
          tmp_112_lpi_3_dfm_1, tmp_44_lpi_3_dfm_1, STD_LOGIC_VECTOR'( (fsm_output(2))
          & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
      tmp_114_lpi_3_dfm_2 <= MUX1HOT_v_32_4_2(tmp_78_lpi_3_dfm_1, tmp_22_lpi_3_dfm_1,
          tmp_114_lpi_3_dfm_1, tmp_46_lpi_3_dfm_1, STD_LOGIC_VECTOR'( (fsm_output(2))
          & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
      tmp_116_lpi_3_dfm_2 <= MUX1HOT_v_32_4_2(tmp_80_lpi_3_dfm_1, tmp_24_lpi_3_dfm_1,
          tmp_116_lpi_3_dfm_1, tmp_48_lpi_3_dfm_1, STD_LOGIC_VECTOR'( (fsm_output(2))
          & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
      tmp_118_lpi_3_dfm_2 <= MUX1HOT_v_32_4_2(tmp_82_lpi_3_dfm_1, tmp_26_lpi_3_dfm_1,
          tmp_118_lpi_3_dfm_1, tmp_50_lpi_3_dfm_1, STD_LOGIC_VECTOR'( (fsm_output(2))
          & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
      tmp_120_lpi_3_dfm_2 <= MUX1HOT_v_32_4_2(tmp_84_lpi_3_dfm_1, tmp_28_lpi_3_dfm_1,
          tmp_120_lpi_3_dfm_1, tmp_52_lpi_3_dfm_1, STD_LOGIC_VECTOR'( (fsm_output(2))
          & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
      tmp_122_lpi_3_dfm_2 <= MUX1HOT_v_32_4_2(tmp_86_lpi_3_dfm_1, tmp_30_lpi_3_dfm_1,
          tmp_122_lpi_3_dfm_1, tmp_54_lpi_3_dfm_1, STD_LOGIC_VECTOR'( (fsm_output(2))
          & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
      tmp_124_lpi_3_dfm_2 <= MUX1HOT_v_32_4_2(tmp_88_lpi_3_dfm_1, tmp_4_lpi_3_dfm_1,
          tmp_124_lpi_3_dfm_1, tmp_56_lpi_3_dfm_1, STD_LOGIC_VECTOR'( (fsm_output(2))
          & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
      tmp_126_lpi_3_dfm_2 <= MUX1HOT_v_32_4_2(tmp_90_lpi_3_dfm_1, tmp_6_lpi_3_dfm_1,
          tmp_126_lpi_3_dfm_1, tmp_58_lpi_3_dfm_1, STD_LOGIC_VECTOR'( (fsm_output(2))
          & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
      tmp_60_lpi_3_dfm_2 <= MUX1HOT_v_32_4_2(tmp_92_lpi_3_dfm_1, tmp_8_lpi_3_dfm_1,
          tmp_96_lpi_3_dfm_1, tmp_60_lpi_3_dfm_1, STD_LOGIC_VECTOR'( (fsm_output(2))
          & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
      tmp_62_lpi_3_dfm_2 <= MUX1HOT_v_32_4_2(tmp_94_lpi_3_dfm_1, tmp_lpi_3_dfm_1,
          tmp_98_lpi_3_dfm_1, tmp_62_lpi_3_dfm_1, STD_LOGIC_VECTOR'( (fsm_output(2))
          & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
      reg_modulo_sub_16_qr_lpi_3_dfm_1_ftd <= (z_out_109(31)) AND (NOT(modulo_sub_16_qelse_and_ssc
          OR modulo_sub_16_qelse_and_ssc_1));
      reg_modulo_sub_16_qr_lpi_3_dfm_1_ftd_1 <= MUX1HOT_v_31_3_2((z_out_126(30 DOWNTO
          0)), (z_out_109(30 DOWNTO 0)), (z_out_111(30 DOWNTO 0)), STD_LOGIC_VECTOR'(
          modulo_sub_16_qelse_and_ssc & modulo_sub_16_qelse_or_nl & modulo_sub_16_qelse_and_ssc_1));
      reg_modulo_sub_17_qr_lpi_3_dfm_1_ftd <= (z_out_106(31)) AND (NOT(modulo_sub_17_qelse_and_ssc
          OR modulo_sub_17_qelse_and_ssc_1));
      reg_modulo_sub_17_qr_lpi_3_dfm_1_ftd_1 <= MUX1HOT_v_31_3_2((z_out_116(30 DOWNTO
          0)), (z_out_106(30 DOWNTO 0)), (z_out_112(30 DOWNTO 0)), STD_LOGIC_VECTOR'(
          modulo_sub_17_qelse_and_ssc & modulo_sub_17_qelse_or_nl & modulo_sub_17_qelse_and_ssc_1));
      reg_modulo_sub_18_qr_lpi_3_dfm_1_ftd <= (z_out_104(31)) AND (NOT(modulo_sub_18_qelse_and_ssc
          OR modulo_sub_18_qelse_and_ssc_1));
      reg_modulo_sub_18_qr_lpi_3_dfm_1_ftd_1 <= MUX1HOT_v_31_3_2((z_out_123(30 DOWNTO
          0)), (z_out_104(30 DOWNTO 0)), (z_out_113(30 DOWNTO 0)), STD_LOGIC_VECTOR'(
          modulo_sub_18_qelse_and_ssc & modulo_sub_18_qelse_or_nl & modulo_sub_18_qelse_and_ssc_1));
      reg_modulo_sub_19_qr_lpi_3_dfm_1_ftd <= (z_out_101(31)) AND (NOT(modulo_sub_19_qelse_and_ssc
          OR modulo_sub_19_qelse_and_ssc_1));
      reg_modulo_sub_19_qr_lpi_3_dfm_1_ftd_1 <= MUX1HOT_v_31_3_2((z_out_124(30 DOWNTO
          0)), (z_out_101(30 DOWNTO 0)), (z_out_114(30 DOWNTO 0)), STD_LOGIC_VECTOR'(
          modulo_sub_19_qelse_and_ssc & modulo_sub_19_qelse_or_nl & modulo_sub_19_qelse_and_ssc_1));
      reg_modulo_sub_20_qr_lpi_3_dfm_1_ftd <= (z_out_98(31)) AND (NOT(modulo_sub_20_qelse_and_ssc
          OR modulo_sub_20_qelse_and_ssc_1));
      reg_modulo_sub_20_qr_lpi_3_dfm_1_ftd_1 <= MUX1HOT_v_31_3_2((z_out_125(30 DOWNTO
          0)), (z_out_98(30 DOWNTO 0)), (z_out_115(30 DOWNTO 0)), STD_LOGIC_VECTOR'(
          modulo_sub_20_qelse_and_ssc & modulo_sub_20_qelse_or_nl & modulo_sub_20_qelse_and_ssc_1));
      reg_modulo_sub_21_qr_lpi_3_dfm_1_ftd <= (z_out_96(31)) AND (NOT(modulo_sub_21_qelse_and_ssc
          OR modulo_sub_21_qelse_and_ssc_1));
      reg_modulo_sub_21_qr_lpi_3_dfm_1_ftd_1 <= MUX1HOT_v_31_3_2((z_out_111(30 DOWNTO
          0)), (z_out_96(30 DOWNTO 0)), (z_out_116(30 DOWNTO 0)), STD_LOGIC_VECTOR'(
          modulo_sub_21_qelse_and_ssc & modulo_sub_21_qelse_or_nl & modulo_sub_21_qelse_and_ssc_1));
      reg_modulo_sub_22_qr_lpi_3_dfm_1_ftd <= (z_out_93(31)) AND (NOT(modulo_sub_22_qelse_and_ssc
          OR modulo_sub_22_qelse_and_ssc_1));
      reg_modulo_sub_22_qr_lpi_3_dfm_1_ftd_1 <= MUX1HOT_v_31_3_2((z_out_112(30 DOWNTO
          0)), (z_out_93(30 DOWNTO 0)), (z_out_117(30 DOWNTO 0)), STD_LOGIC_VECTOR'(
          modulo_sub_22_qelse_and_ssc & modulo_sub_22_qelse_or_nl & modulo_sub_22_qelse_and_ssc_1));
      reg_modulo_sub_23_qr_lpi_3_dfm_1_ftd <= (z_out_90(31)) AND (NOT(modulo_sub_23_qelse_and_ssc
          OR modulo_sub_23_qelse_and_ssc_1));
      reg_modulo_sub_23_qr_lpi_3_dfm_1_ftd_1 <= MUX1HOT_v_31_3_2((z_out_113(30 DOWNTO
          0)), (z_out_90(30 DOWNTO 0)), (z_out_118(30 DOWNTO 0)), STD_LOGIC_VECTOR'(
          modulo_sub_23_qelse_and_ssc & modulo_sub_23_qelse_or_nl & modulo_sub_23_qelse_and_ssc_1));
      reg_modulo_sub_24_qr_lpi_3_dfm_1_ftd <= (z_out_88(31)) AND (NOT(modulo_sub_24_qelse_and_ssc
          OR modulo_sub_24_qelse_and_ssc_1));
      reg_modulo_sub_24_qr_lpi_3_dfm_1_ftd_1 <= MUX1HOT_v_31_3_2((z_out_114(30 DOWNTO
          0)), (z_out_88(30 DOWNTO 0)), (z_out_119(30 DOWNTO 0)), STD_LOGIC_VECTOR'(
          modulo_sub_24_qelse_and_ssc & modulo_sub_24_qelse_or_nl & modulo_sub_24_qelse_and_ssc_1));
      reg_modulo_sub_25_qr_lpi_3_dfm_1_ftd <= (z_out_85(31)) AND (NOT(modulo_sub_25_qelse_and_ssc
          OR modulo_sub_25_qelse_and_ssc_1));
      reg_modulo_sub_25_qr_lpi_3_dfm_1_ftd_1 <= MUX1HOT_v_31_3_2((z_out_115(30 DOWNTO
          0)), (z_out_85(30 DOWNTO 0)), (z_out_120(30 DOWNTO 0)), STD_LOGIC_VECTOR'(
          modulo_sub_25_qelse_and_ssc & modulo_sub_25_qelse_or_nl & modulo_sub_25_qelse_and_ssc_1));
      reg_modulo_sub_26_qr_lpi_3_dfm_1_ftd <= (z_out_82(31)) AND (NOT(modulo_sub_26_qelse_and_ssc
          OR modulo_sub_26_qelse_and_ssc_1));
      reg_modulo_sub_26_qr_lpi_3_dfm_1_ftd_1 <= MUX1HOT_v_31_3_2((z_out_117(30 DOWNTO
          0)), (z_out_82(30 DOWNTO 0)), (z_out_121(30 DOWNTO 0)), STD_LOGIC_VECTOR'(
          modulo_sub_26_qelse_and_ssc & modulo_sub_26_qelse_or_nl & modulo_sub_26_qelse_and_ssc_1));
      reg_modulo_sub_27_qr_lpi_3_dfm_1_ftd <= (z_out_80(31)) AND (NOT(modulo_sub_27_qelse_and_ssc
          OR modulo_sub_27_qelse_and_ssc_1));
      reg_modulo_sub_27_qr_lpi_3_dfm_1_ftd_1 <= MUX1HOT_v_31_3_2((z_out_118(30 DOWNTO
          0)), (z_out_80(30 DOWNTO 0)), (z_out_122(30 DOWNTO 0)), STD_LOGIC_VECTOR'(
          modulo_sub_27_qelse_and_ssc & modulo_sub_27_qelse_or_nl & modulo_sub_27_qelse_and_ssc_1));
      reg_modulo_sub_28_qr_lpi_3_dfm_1_ftd <= (z_out_77(31)) AND (NOT(modulo_sub_28_qelse_and_ssc
          OR modulo_sub_28_qelse_and_ssc_1));
      reg_modulo_sub_28_qr_lpi_3_dfm_1_ftd_1 <= MUX1HOT_v_31_3_2((z_out_119(30 DOWNTO
          0)), (z_out_77(30 DOWNTO 0)), (z_out_123(30 DOWNTO 0)), STD_LOGIC_VECTOR'(
          modulo_sub_28_qelse_and_ssc & modulo_sub_28_qelse_or_nl & modulo_sub_28_qelse_and_ssc_1));
      reg_modulo_sub_29_qr_lpi_3_dfm_1_ftd <= (z_out_74(31)) AND (NOT(modulo_sub_29_qelse_and_ssc
          OR modulo_sub_29_qelse_and_ssc_1));
      reg_modulo_sub_29_qr_lpi_3_dfm_1_ftd_1 <= MUX1HOT_v_31_3_2((z_out_120(30 DOWNTO
          0)), (z_out_74(30 DOWNTO 0)), (z_out_124(30 DOWNTO 0)), STD_LOGIC_VECTOR'(
          modulo_sub_29_qelse_and_ssc & modulo_sub_29_qelse_or_nl & modulo_sub_29_qelse_and_ssc_1));
      reg_modulo_sub_30_qr_lpi_3_dfm_1_ftd <= (z_out_72(31)) AND (NOT(modulo_sub_30_qelse_and_ssc
          OR modulo_sub_30_qelse_and_ssc_1));
      reg_modulo_sub_30_qr_lpi_3_dfm_1_ftd_1 <= MUX1HOT_v_31_3_2((z_out_121(30 DOWNTO
          0)), (z_out_72(30 DOWNTO 0)), (z_out_125(30 DOWNTO 0)), STD_LOGIC_VECTOR'(
          modulo_sub_30_qelse_and_ssc & modulo_sub_30_qelse_or_nl & modulo_sub_30_qelse_and_ssc_1));
      reg_modulo_sub_31_qr_lpi_3_dfm_1_ftd <= (z_out_69(31)) AND (NOT(modulo_sub_31_qelse_and_ssc
          OR modulo_sub_31_qelse_and_ssc_1));
      reg_modulo_sub_31_qr_lpi_3_dfm_1_ftd_1 <= MUX1HOT_v_31_3_2((z_out_122(30 DOWNTO
          0)), (z_out_69(30 DOWNTO 0)), (z_out_126(30 DOWNTO 0)), STD_LOGIC_VECTOR'(
          modulo_sub_31_qelse_and_ssc & modulo_sub_31_qelse_or_nl & modulo_sub_31_qelse_and_ssc_1));
      INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9472_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_9855_itm_8;
      INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9855_itm_1 <= MUX_v_4_2_2((INNER_LOOP2_r_11_4_sva_6_0(4
          DOWNTO 1)), (INNER_LOOP4_r_11_4_sva_6_0(4 DOWNTO 1)), fsm_output(9));
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        butterFly1_15_conc_2_itm_9_2_1 <= STD_LOGIC_VECTOR'( "00");
      ELSIF ( (butterFly1_15_conc_2_itm_5_0 OR butterFly2_15_conc_2_itm_5_0) = '1'
          ) THEN
        butterFly1_15_conc_2_itm_9_2_1 <= butterFly1_15_conc_2_itm_8_2_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (butterFly1_15_conc_2_itm_4_0 OR butterFly1_15_conc_2_itm_9_0 OR or_dcpl_19)
          = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_8833_itm_8 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12410_itm_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (butterFly1_15_conc_2_itm_3_0 OR butterFly1_15_conc_2_itm_9_0 OR or_dcpl_22)
          = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_9344_itm_8 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12921_itm_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (butterFly1_15_conc_2_itm_2_0 OR butterFly1_15_conc_2_itm_9_0 OR or_dcpl_25)
          = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_9855_itm_8 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13432_itm_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (butterFly1_15_conc_2_itm_8_0 OR butterFly1_15_conc_2_itm_9_0 OR butterFly2_15_conc_2_itm_4_0)
          = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_10366_itm_8 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14965_itm_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (butterFly1_15_conc_2_itm_7_0 OR butterFly1_15_conc_2_itm_9_0 OR or_dcpl_30)
          = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_10877_itm_8 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15476_itm_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (butterFly1_15_conc_2_itm_6_0 OR butterFly1_15_conc_2_itm_9_0 OR or_dcpl_33)
          = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_11388_itm_8 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15987_itm_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (butterFly1_15_conc_2_itm_5_0 OR butterFly1_15_conc_2_itm_9_0 OR or_dcpl_36)
          = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_11899_itm_8 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16498_itm_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (butterFly1_15_conc_2_itm_9_0 OR butterFly2_15_conc_2_itm_4_0 OR butterFly2_15_conc_2_itm_5_0)
          = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14454_itm_8 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14454_itm_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        butterFly1_15_conc_2_itm_8_2_1 <= STD_LOGIC_VECTOR'( "00");
      ELSIF ( (butterFly1_15_conc_2_itm_4_0 OR butterFly2_15_conc_2_itm_4_0) = '1'
          ) THEN
        butterFly1_15_conc_2_itm_8_2_1 <= butterFly1_15_conc_2_itm_7_2_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( butterFly2_15_conc_2_itm_4_0 = '1' ) THEN
        reg_mult_15_res_lpi_3_dfm_1_cse <= mult_15_res_lpi_3_dfm_1_mx0;
        reg_mult_14_res_lpi_3_dfm_1_cse <= mult_14_res_lpi_3_dfm_1_mx0;
        reg_mult_13_res_lpi_3_dfm_1_cse <= mult_13_res_lpi_3_dfm_1_mx0;
        reg_mult_12_res_lpi_3_dfm_1_cse <= mult_12_res_lpi_3_dfm_1_mx0;
        reg_mult_11_res_lpi_3_dfm_1_cse <= mult_11_res_lpi_3_dfm_1_mx0;
        reg_mult_10_res_lpi_3_dfm_1_cse <= mult_10_res_lpi_3_dfm_1_mx0;
        reg_mult_9_res_lpi_3_dfm_1_cse <= mult_9_res_lpi_3_dfm_1_mx0;
        reg_mult_8_res_lpi_3_dfm_1_cse <= mult_8_res_lpi_3_dfm_1_mx0;
        reg_mult_7_res_lpi_3_dfm_1_cse <= mult_7_res_lpi_3_dfm_1_mx0;
        reg_mult_6_res_lpi_3_dfm_1_cse <= mult_6_res_lpi_3_dfm_1_mx0;
        reg_mult_5_res_lpi_3_dfm_1_cse <= mult_5_res_lpi_3_dfm_1_mx0;
        reg_mult_4_res_lpi_3_dfm_1_cse <= mult_4_res_lpi_3_dfm_1_mx0;
        reg_mult_3_res_lpi_3_dfm_1_cse <= mult_3_res_lpi_3_dfm_1_mx0;
        reg_mult_2_res_lpi_3_dfm_1_cse <= mult_2_res_lpi_3_dfm_1_mx0;
        reg_mult_1_res_lpi_3_dfm_1_cse <= mult_1_res_lpi_3_dfm_1_mx0;
        reg_mult_res_lpi_3_dfm_1_cse <= mult_res_lpi_3_dfm_1_mx0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1 <= STD_LOGIC_VECTOR'( "000");
        butterFly1_15_conc_2_itm_1_2_1 <= STD_LOGIC_VECTOR'( "00");
        butterFly2_15_tw_equal_tmp_1 <= '0';
        butterFly2_15_tw_equal_tmp_3_1 <= '0';
        butterFly2_15_tw_equal_tmp_5_1 <= '0';
        butterFly2_15_tw_equal_tmp_6_1 <= '0';
        butterFly2_15_tw_equal_tmp_7_1 <= '0';
      ELSIF ( INNER_LOOP1_stage_0 = '1' ) THEN
        butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1 <= butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm;
        butterFly1_15_conc_2_itm_1_2_1 <= butterFly1_15_conc_2_itm_2_1;
        butterFly2_15_tw_equal_tmp_1 <= NOT(CONV_SL_1_1(operator_20_false_acc_cse_sva/=STD_LOGIC_VECTOR'("000")));
        butterFly2_15_tw_equal_tmp_3_1 <= CONV_SL_1_1(operator_20_false_acc_cse_sva=STD_LOGIC_VECTOR'("011"));
        butterFly2_15_tw_equal_tmp_5_1 <= CONV_SL_1_1(operator_20_false_acc_cse_sva=STD_LOGIC_VECTOR'("101"));
        butterFly2_15_tw_equal_tmp_6_1 <= CONV_SL_1_1(operator_20_false_acc_cse_sva=STD_LOGIC_VECTOR'("110"));
        butterFly2_15_tw_equal_tmp_7_1 <= CONV_SL_1_1(operator_20_false_acc_cse_sva=STD_LOGIC_VECTOR'("111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        operator_20_false_acc_cse_sva <= STD_LOGIC_VECTOR'( "000");
      ELSIF ( (NOT(or_dcpl_315 OR or_dcpl_353)) = '1' ) THEN
        operator_20_false_acc_cse_sva <= MUX_v_3_2_2(z_out_61, (z_out_60(2 DOWNTO
            0)), fsm_output(6));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        butterFly1_15_conc_2_itm_7_2_1 <= STD_LOGIC_VECTOR'( "00");
      ELSIF ( (butterFly1_15_conc_2_itm_3_0 OR butterFly2_15_conc_2_itm_3_0) = '1'
          ) THEN
        butterFly1_15_conc_2_itm_7_2_1 <= butterFly1_15_conc_2_itm_6_2_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (butterFly1_15_conc_2_itm_4_0 OR butterFly2_15_conc_2_itm_3_0 OR butterFly1_15_conc_2_itm_8_0
          OR butterFly2_15_conc_2_itm_0) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16498_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16498_itm_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (butterFly1_15_conc_2_itm_5_0 OR butterFly1_15_conc_2_itm_8_0 OR or_dcpl_36)
          = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16115_itm_8 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16115_itm_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( or_dcpl_12 = '1' ) THEN
        mult_15_z_asn_itm_2 <= mult_15_z_asn_itm_1;
        mult_14_z_asn_itm_2 <= mult_14_z_asn_itm_1;
        mult_13_z_asn_itm_2 <= mult_13_z_asn_itm_1;
        mult_12_z_asn_itm_2 <= mult_12_z_asn_itm_1;
        mult_11_z_asn_itm_2 <= mult_11_z_asn_itm_1;
        mult_10_z_asn_itm_2 <= mult_10_z_asn_itm_1;
        mult_1_z_asn_itm_2 <= mult_1_z_asn_itm_1;
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14582_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14582_itm_5;
        mult_23_z_asn_itm_2 <= mult_23_z_asn_itm_1;
        mult_24_z_asn_itm_2 <= mult_24_z_asn_itm_1;
        mult_25_z_asn_itm_2 <= mult_25_z_asn_itm_1;
        mult_26_z_asn_itm_2 <= mult_26_z_asn_itm_1;
        mult_27_z_asn_itm_2 <= mult_27_z_asn_itm_1;
        mult_28_z_asn_itm_2 <= mult_28_z_asn_itm_1;
        mult_29_z_asn_itm_2 <= mult_29_z_asn_itm_1;
        mult_30_z_asn_itm_2 <= mult_30_z_asn_itm_1;
        mult_31_z_asn_itm_2 <= mult_31_z_asn_itm_1;
        tmp_10_lpi_3_dfm_5 <= tmp_10_lpi_3_dfm_4;
        tmp_102_lpi_3_dfm_5 <= tmp_102_lpi_3_dfm_4;
        tmp_104_lpi_3_dfm_5 <= tmp_104_lpi_3_dfm_4;
        tmp_106_lpi_3_dfm_5 <= tmp_106_lpi_3_dfm_4;
        tmp_108_lpi_3_dfm_5 <= tmp_108_lpi_3_dfm_4;
        tmp_110_lpi_3_dfm_5 <= tmp_110_lpi_3_dfm_4;
        tmp_112_lpi_3_dfm_5 <= tmp_112_lpi_3_dfm_4;
        tmp_114_lpi_3_dfm_5 <= tmp_114_lpi_3_dfm_4;
        tmp_116_lpi_3_dfm_5 <= tmp_116_lpi_3_dfm_4;
        tmp_118_lpi_3_dfm_5 <= tmp_118_lpi_3_dfm_4;
        tmp_120_lpi_3_dfm_5 <= tmp_120_lpi_3_dfm_4;
        tmp_122_lpi_3_dfm_5 <= tmp_122_lpi_3_dfm_4;
        tmp_124_lpi_3_dfm_5 <= tmp_124_lpi_3_dfm_4;
        tmp_126_lpi_3_dfm_5 <= tmp_126_lpi_3_dfm_4;
        tmp_60_lpi_3_dfm_5 <= tmp_60_lpi_3_dfm_4;
        tmp_62_lpi_3_dfm_5 <= tmp_62_lpi_3_dfm_4;
        INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9855_itm_6 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9855_itm_5;
        INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9472_itm_6 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9472_itm_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (butterFly1_15_conc_2_itm_5_0 OR butterFly2_15_conc_2_itm_3_0 OR butterFly1_15_conc_2_itm_8_0
          OR butterFly2_15_conc_2_itm_1_0) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15987_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15987_itm_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (butterFly1_15_conc_2_itm_6_0 OR butterFly1_15_conc_2_itm_8_0 OR or_dcpl_33)
          = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15604_itm_8 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15604_itm_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (butterFly1_15_conc_2_itm_6_0 OR butterFly2_15_conc_2_itm_3_0 OR butterFly1_15_conc_2_itm_8_0
          OR butterFly2_15_conc_2_itm_2_0) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15476_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15476_itm_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_63 OR or_dcpl_30) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15093_itm_8 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15093_itm_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_63 OR butterFly2_15_conc_2_itm_3_0) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14965_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14965_itm_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( or_dcpl_8 = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14582_itm_8 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14582_itm_7;
        tmp_10_lpi_3_dfm_7 <= tmp_10_lpi_3_dfm_6;
        tmp_102_lpi_3_dfm_7 <= tmp_102_lpi_3_dfm_6;
        tmp_104_lpi_3_dfm_7 <= tmp_104_lpi_3_dfm_6;
        tmp_106_lpi_3_dfm_7 <= tmp_106_lpi_3_dfm_6;
        tmp_108_lpi_3_dfm_7 <= tmp_108_lpi_3_dfm_6;
        tmp_110_lpi_3_dfm_7 <= tmp_110_lpi_3_dfm_6;
        tmp_112_lpi_3_dfm_7 <= tmp_112_lpi_3_dfm_6;
        tmp_114_lpi_3_dfm_7 <= tmp_114_lpi_3_dfm_6;
        tmp_116_lpi_3_dfm_7 <= tmp_116_lpi_3_dfm_6;
        tmp_118_lpi_3_dfm_7 <= tmp_118_lpi_3_dfm_6;
        tmp_120_lpi_3_dfm_7 <= tmp_120_lpi_3_dfm_6;
        tmp_122_lpi_3_dfm_7 <= tmp_122_lpi_3_dfm_6;
        tmp_124_lpi_3_dfm_7 <= tmp_124_lpi_3_dfm_6;
        tmp_126_lpi_3_dfm_7 <= tmp_126_lpi_3_dfm_6;
        tmp_60_lpi_3_dfm_7 <= tmp_60_lpi_3_dfm_6;
        tmp_62_lpi_3_dfm_7 <= tmp_62_lpi_3_dfm_6;
        INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9855_itm_8 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9855_itm_7;
        INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9472_itm_8 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9472_itm_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (butterFly1_15_conc_2_itm_8_0 OR butterFly2_15_conc_2_itm_3_0 OR butterFly2_15_conc_2_itm_4_0)
          = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14454_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14454_itm_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_70 OR butterFly2_15_conc_2_itm_4_0 OR butterFly2_15_conc_2_itm_5_0)
          = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14071_itm_8 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14071_itm_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_70 OR or_dcpl_72) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13943_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13943_itm_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_76 OR or_dcpl_25) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13049_itm_8 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13049_itm_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_76 OR or_dcpl_78) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12921_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12921_itm_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_80 OR or_dcpl_22) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12538_itm_8 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12538_itm_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_80 OR or_dcpl_82) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12410_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12410_itm_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (butterFly1_15_conc_2_itm_4_0 OR butterFly1_15_conc_2_itm_8_0 OR or_dcpl_19)
          = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12027_itm_8 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12027_itm_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        butterFly1_15_conc_2_itm_6_2_1 <= STD_LOGIC_VECTOR'( "00");
      ELSIF ( (butterFly1_15_conc_2_itm_2_0 OR butterFly2_15_conc_2_itm_2_0) = '1'
          ) THEN
        butterFly1_15_conc_2_itm_6_2_1 <= butterFly1_15_conc_2_itm_5_2_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_89 OR or_dcpl_88) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16498_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16498_itm_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_10 OR or_dcpl_2) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16115_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16115_itm_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_94 OR or_dcpl_2) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15987_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15987_itm_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_10 OR or_dcpl) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15604_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15604_itm_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_94 OR or_dcpl) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15476_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15476_itm_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_10 OR or_dcpl_12) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15093_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15093_itm_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (butterFly1_15_conc_2_itm_7_0 OR butterFly1_15_conc_2_itm_6_0 OR butterFly2_15_conc_2_itm_2_0)
          = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14965_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14965_itm_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( or_dcpl_10 = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14582_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14582_itm_6;
        tmp_10_lpi_3_dfm_6 <= tmp_10_lpi_3_dfm_5;
        tmp_102_lpi_3_dfm_6 <= tmp_102_lpi_3_dfm_5;
        tmp_104_lpi_3_dfm_6 <= tmp_104_lpi_3_dfm_5;
        tmp_106_lpi_3_dfm_6 <= tmp_106_lpi_3_dfm_5;
        tmp_108_lpi_3_dfm_6 <= tmp_108_lpi_3_dfm_5;
        tmp_110_lpi_3_dfm_6 <= tmp_110_lpi_3_dfm_5;
        tmp_112_lpi_3_dfm_6 <= tmp_112_lpi_3_dfm_5;
        tmp_114_lpi_3_dfm_6 <= tmp_114_lpi_3_dfm_5;
        tmp_116_lpi_3_dfm_6 <= tmp_116_lpi_3_dfm_5;
        tmp_118_lpi_3_dfm_6 <= tmp_118_lpi_3_dfm_5;
        tmp_120_lpi_3_dfm_6 <= tmp_120_lpi_3_dfm_5;
        tmp_122_lpi_3_dfm_6 <= tmp_122_lpi_3_dfm_5;
        tmp_124_lpi_3_dfm_6 <= tmp_124_lpi_3_dfm_5;
        tmp_126_lpi_3_dfm_6 <= tmp_126_lpi_3_dfm_5;
        tmp_60_lpi_3_dfm_6 <= tmp_60_lpi_3_dfm_5;
        tmp_62_lpi_3_dfm_6 <= tmp_62_lpi_3_dfm_5;
        INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9855_itm_7 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9855_itm_6;
        INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9472_itm_7 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9472_itm_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (butterFly1_15_conc_2_itm_7_0 OR butterFly2_15_conc_2_itm_2_0 OR butterFly2_15_conc_2_itm_3_0)
          = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14454_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14454_itm_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_10 OR or_dcpl_8) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14071_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14071_itm_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_94 OR or_dcpl_8) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13943_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13943_itm_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_105 OR or_dcpl_72) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13560_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13560_itm_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_105 OR or_dcpl_107) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13432_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13432_itm_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_109 OR or_dcpl_78) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12538_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12538_itm_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_109 OR or_dcpl_111) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12410_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12410_itm_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_89 OR or_dcpl_82) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12027_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12027_itm_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        butterFly1_15_conc_2_itm_5_2_1 <= STD_LOGIC_VECTOR'( "00");
      ELSIF ( (INNER_LOOP1_stage_0 OR butterFly2_15_conc_2_itm_1_0) = '1' ) THEN
        butterFly1_15_conc_2_itm_5_2_1 <= butterFly1_15_conc_2_itm_4_2_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_117 OR or_dcpl_116) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16498_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16498_itm_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_119 OR or_dcpl_88) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16115_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16115_itm_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_119 OR or_dcpl_121) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15987_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15987_itm_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_12 OR or_dcpl_2) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15604_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15604_itm_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_125 OR or_dcpl_2) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15476_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15476_itm_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_12 OR or_dcpl) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15093_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15093_itm_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (butterFly1_15_conc_2_itm_6_0 OR butterFly1_15_conc_2_itm_5_0 OR butterFly2_15_conc_2_itm_1_0)
          = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14965_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14965_itm_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (butterFly1_15_conc_2_itm_6_0 OR butterFly2_15_conc_2_itm_1_0 OR butterFly2_15_conc_2_itm_2_0)
          = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14454_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14454_itm_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_133 OR butterFly2_15_conc_2_itm_2_0 OR butterFly2_15_conc_2_itm_3_0)
          = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14071_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14071_itm_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_133 OR or_dcpl_135) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13943_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13943_itm_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_12 OR or_dcpl_8) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13560_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13560_itm_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_125 OR or_dcpl_8) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13432_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13432_itm_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_139 OR or_dcpl_107) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13049_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13049_itm_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_139 OR or_dcpl_141) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12921_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12921_itm_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_117 OR or_dcpl_111) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12027_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12027_itm_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_146 OR or_dcpl_116) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16115_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16115_itm_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_146 OR or_dcpl_148) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15987_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15987_itm_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_150 OR or_dcpl_121) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15604_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15604_itm_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_150 OR or_dcpl_152) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15476_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15476_itm_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl OR or_dcpl_2) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15093_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15093_itm_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (butterFly1_15_conc_2_itm_5_0 OR butterFly1_15_conc_2_itm_4_0 OR butterFly2_15_conc_2_itm_0)
          = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14965_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14965_itm_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( or_dcpl = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14582_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14582_itm_4;
        tmp_10_lpi_3_dfm_4 <= tmp_10_lpi_3_dfm_3;
        tmp_102_lpi_3_dfm_4 <= tmp_102_lpi_3_dfm_3;
        tmp_104_lpi_3_dfm_4 <= tmp_104_lpi_3_dfm_3;
        tmp_106_lpi_3_dfm_4 <= tmp_106_lpi_3_dfm_3;
        tmp_108_lpi_3_dfm_4 <= tmp_108_lpi_3_dfm_3;
        tmp_110_lpi_3_dfm_4 <= tmp_110_lpi_3_dfm_3;
        tmp_112_lpi_3_dfm_4 <= tmp_112_lpi_3_dfm_3;
        tmp_114_lpi_3_dfm_4 <= tmp_114_lpi_3_dfm_3;
        tmp_116_lpi_3_dfm_4 <= tmp_116_lpi_3_dfm_3;
        tmp_118_lpi_3_dfm_4 <= tmp_118_lpi_3_dfm_3;
        tmp_120_lpi_3_dfm_4 <= tmp_120_lpi_3_dfm_3;
        tmp_122_lpi_3_dfm_4 <= tmp_122_lpi_3_dfm_3;
        tmp_124_lpi_3_dfm_4 <= tmp_124_lpi_3_dfm_3;
        tmp_126_lpi_3_dfm_4 <= tmp_126_lpi_3_dfm_3;
        tmp_60_lpi_3_dfm_4 <= tmp_60_lpi_3_dfm_3;
        tmp_62_lpi_3_dfm_4 <= tmp_62_lpi_3_dfm_3;
        INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9855_itm_5 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9855_itm_4;
        INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9472_itm_5 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9472_itm_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (butterFly1_15_conc_2_itm_5_0 OR butterFly2_15_conc_2_itm_0 OR butterFly2_15_conc_2_itm_1_0)
          = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14454_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14454_itm_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_161 OR butterFly2_15_conc_2_itm_1_0 OR butterFly2_15_conc_2_itm_2_0)
          = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14071_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14071_itm_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_161 OR or_dcpl_163) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13943_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13943_itm_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_165 OR or_dcpl_135) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13560_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13560_itm_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_165 OR or_dcpl_167) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13432_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13432_itm_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl OR or_dcpl_8) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13049_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13049_itm_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (butterFly1_15_conc_2_itm_5_0 OR butterFly2_15_conc_2_itm_0 OR or_dcpl_8)
          = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12921_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12921_itm_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_171 OR or_dcpl_141) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12538_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12538_itm_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_171 OR or_dcpl_173) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12410_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12410_itm_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        butterFly1_15_conc_2_itm_3_2_1 <= STD_LOGIC_VECTOR'( "00");
      ELSIF ( (INNER_LOOP1_stage_0 OR INNER_LOOP1_stage_0_3 OR butterFly2_15_conc_2_itm_8_0)
          = '1' ) THEN
        butterFly1_15_conc_2_itm_3_2_1 <= butterFly1_15_conc_2_itm_2_2_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_181 OR or_dcpl_180) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16498_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16498_itm_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_185 OR or_dcpl_148) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15604_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15604_itm_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_185 OR or_dcpl_187) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15476_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15476_itm_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_189 OR or_dcpl_152) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15093_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15093_itm_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_189 OR INNER_LOOP1_stage_0_3 OR butterFly2_15_conc_2_itm_8_0)
          = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14965_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14965_itm_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( or_dcpl_2 = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14582_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14582_itm_3;
        tmp_10_lpi_3_dfm_3 <= tmp_10_lpi_3_dfm_2;
        tmp_102_lpi_3_dfm_3 <= tmp_102_lpi_3_dfm_2;
        tmp_104_lpi_3_dfm_3 <= tmp_104_lpi_3_dfm_2;
        tmp_106_lpi_3_dfm_3 <= tmp_106_lpi_3_dfm_2;
        tmp_108_lpi_3_dfm_3 <= tmp_108_lpi_3_dfm_2;
        tmp_110_lpi_3_dfm_3 <= tmp_110_lpi_3_dfm_2;
        tmp_112_lpi_3_dfm_3 <= tmp_112_lpi_3_dfm_2;
        tmp_114_lpi_3_dfm_3 <= tmp_114_lpi_3_dfm_2;
        tmp_116_lpi_3_dfm_3 <= tmp_116_lpi_3_dfm_2;
        tmp_118_lpi_3_dfm_3 <= tmp_118_lpi_3_dfm_2;
        tmp_120_lpi_3_dfm_3 <= tmp_120_lpi_3_dfm_2;
        tmp_122_lpi_3_dfm_3 <= tmp_122_lpi_3_dfm_2;
        tmp_124_lpi_3_dfm_3 <= tmp_124_lpi_3_dfm_2;
        tmp_126_lpi_3_dfm_3 <= tmp_126_lpi_3_dfm_2;
        tmp_60_lpi_3_dfm_3 <= tmp_60_lpi_3_dfm_2;
        tmp_62_lpi_3_dfm_3 <= tmp_62_lpi_3_dfm_2;
        INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9855_itm_4 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9855_itm_3;
        INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9472_itm_4 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9472_itm_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (butterFly1_15_conc_2_itm_4_0 OR INNER_LOOP1_stage_0_3 OR butterFly2_15_conc_2_itm_0)
          = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14454_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14454_itm_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_197 OR butterFly2_15_conc_2_itm_0 OR butterFly2_15_conc_2_itm_1_0)
          = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14071_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14071_itm_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_197 OR or_dcpl_199) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13943_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13943_itm_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_201 OR or_dcpl_163) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13560_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13560_itm_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_201 OR or_dcpl_203) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13432_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13432_itm_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_205 OR or_dcpl_167) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13049_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13049_itm_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_205 OR or_dcpl_207) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12921_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12921_itm_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (butterFly1_15_conc_2_itm_4_0 OR butterFly2_15_conc_2_itm_0 OR or_dcpl_8)
          = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12538_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12538_itm_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (butterFly1_15_conc_2_itm_4_0 OR butterFly1_15_conc_2_itm_8_0 OR or_dcpl_210)
          = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12410_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12410_itm_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_181 OR or_dcpl_173) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12027_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12027_itm_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_80 OR or_dcpl_215) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16498_itm_2 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16498_itm_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_218 OR or_dcpl_180) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16115_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16115_itm_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_218 OR or_dcpl_220) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15987_itm_2 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15987_itm_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_224 OR or_dcpl_187) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15093_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15093_itm_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_224 OR INNER_LOOP1_stage_0_2 OR butterFly2_15_conc_2_itm_7_0)
          = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14965_itm_2 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14965_itm_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (butterFly1_15_conc_2_itm_3_0 OR INNER_LOOP1_stage_0_3 OR butterFly2_15_conc_2_itm_8_0)
          = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14582_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14582_itm_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (butterFly1_15_conc_2_itm_3_0 OR INNER_LOOP1_stage_0_2 OR butterFly2_15_conc_2_itm_8_0)
          = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14454_itm_2 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14454_itm_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_189 OR INNER_LOOP1_stage_0_3 OR butterFly2_15_conc_2_itm_0) =
          '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14071_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14071_itm_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_189 OR or_dcpl_234) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13943_itm_2 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13943_itm_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_150 OR or_dcpl_199) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13560_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13560_itm_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_150 OR or_dcpl_238) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13432_itm_2 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13432_itm_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_119 OR or_dcpl_203) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13049_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13049_itm_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_119 OR or_dcpl_242) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12921_itm_2 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12921_itm_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_89 OR or_dcpl_207) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12538_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12538_itm_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_89 OR or_dcpl_246) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12410_itm_2 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12410_itm_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_80 OR or_dcpl_210) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12027_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12027_itm_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( INNER_LOOP1_stage_0_2 = '1' ) THEN
        tmp_94_lpi_3_dfm_1 <= z_out;
        tmp_92_lpi_3_dfm_1 <= z_out_1;
        tmp_90_lpi_3_dfm_1 <= z_out_2;
        tmp_88_lpi_3_dfm_1 <= z_out_3;
        tmp_86_lpi_3_dfm_1 <= z_out_4;
        tmp_84_lpi_3_dfm_1 <= z_out_5;
        tmp_82_lpi_3_dfm_1 <= z_out_6;
        tmp_80_lpi_3_dfm_1 <= z_out_7;
        tmp_78_lpi_3_dfm_1 <= z_out_8;
        tmp_76_lpi_3_dfm_1 <= z_out_9;
        tmp_74_lpi_3_dfm_1 <= z_out_10;
        tmp_72_lpi_3_dfm_1 <= z_out_11;
        tmp_70_lpi_3_dfm_1 <= z_out_12;
        tmp_68_lpi_3_dfm_1 <= z_out_13;
        tmp_66_lpi_3_dfm_1 <= z_out_14;
        tmp_64_lpi_3_dfm_1 <= z_out_15;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (butterFly1_15_conc_2_itm_2_0 OR butterFly1_15_conc_2_itm_8_0 OR or_dcpl_215)
          = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16115_itm_2 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16115_itm_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (butterFly1_15_conc_2_itm_2_0 OR butterFly1_15_conc_2_itm_9_0 OR or_dcpl_220)
          = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15604_itm_2 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15604_itm_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (butterFly1_15_conc_2_itm_2_0 OR INNER_LOOP1_stage_0_2 OR butterFly2_15_conc_2_itm_7_0)
          = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14582_itm_2 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14582_itm_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (butterFly1_15_conc_2_itm_2_0 OR butterFly1_15_conc_2_itm_3_0 OR INNER_LOOP1_stage_0_2
          OR butterFly2_15_conc_2_itm_8_0) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14071_itm_2 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14071_itm_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (butterFly1_15_conc_2_itm_2_0 OR butterFly1_15_conc_2_itm_4_0 OR or_dcpl_234)
          = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13560_itm_2 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13560_itm_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (butterFly1_15_conc_2_itm_2_0 OR butterFly1_15_conc_2_itm_5_0 OR or_dcpl_238)
          = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13049_itm_2 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13049_itm_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (butterFly1_15_conc_2_itm_2_0 OR butterFly1_15_conc_2_itm_6_0 OR or_dcpl_242)
          = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12538_itm_2 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12538_itm_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (butterFly1_15_conc_2_itm_2_0 OR butterFly1_15_conc_2_itm_7_0 OR or_dcpl_246)
          = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12027_itm_2 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12027_itm_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        INNER_LOOP2_r_11_4_sva_6_0 <= STD_LOGIC_VECTOR'( "0000000");
      ELSIF ( (fsm_output(2)) = '0' ) THEN
        INNER_LOOP2_r_11_4_sva_6_0 <= MUX_v_7_2_2(STD_LOGIC_VECTOR'("0000000"), STAGE_LOOP_base_STAGE_LOOP_base_mux_nl,
            INNER_LOOP2_r_or_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        butterFly2_15_conc_2_itm_6_2_1 <= STD_LOGIC_VECTOR'( "00");
      ELSIF ( (butterFly1_15_conc_2_itm_6_0 OR INNER_LOOP1_stage_0_10) = '1' ) THEN
        butterFly2_15_conc_2_itm_6_2_1 <= butterFly1_15_conc_2_itm_9_2_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( or_dcpl_274 = '1' ) THEN
        INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9472_itm_9 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9472_itm_8;
        INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9855_itm_9 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9855_itm_8;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(4)) = '0' ) THEN
        operator_33_true_1_lshift_psp_9_4_sva <= z_out_60(9 DOWNTO 4);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (butterFly1_15_conc_2_itm_3_0 OR butterFly2_15_conc_2_itm_8_0) = '1' )
          THEN
        INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9855_itm_3 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9855_itm_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( butterFly2_15_conc_2_itm_7_0 = '1' ) THEN
        tmp_30_lpi_3_dfm_1 <= z_out_16;
        tmp_28_lpi_3_dfm_1 <= z_out_17;
        tmp_26_lpi_3_dfm_1 <= z_out_18;
        tmp_24_lpi_3_dfm_1 <= z_out_19;
        tmp_22_lpi_3_dfm_1 <= z_out_20;
        tmp_20_lpi_3_dfm_1 <= z_out_21;
        tmp_18_lpi_3_dfm_1 <= z_out_22;
        tmp_16_lpi_3_dfm_1 <= z_out_23;
        tmp_14_lpi_3_dfm_1 <= z_out_24;
        tmp_12_lpi_3_dfm_1 <= z_out_25;
        tmp_10_lpi_3_dfm_1 <= z_out_26;
        tmp_8_lpi_3_dfm_1 <= z_out_27;
        tmp_6_lpi_3_dfm_1 <= z_out_28;
        tmp_4_lpi_3_dfm_1 <= z_out_29;
        tmp_2_lpi_3_dfm_1 <= z_out_30;
        tmp_lpi_3_dfm_1 <= z_out_31;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (butterFly1_15_conc_2_itm_2_0 OR butterFly2_15_conc_2_itm_7_0) = '1' )
          THEN
        INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9855_itm_2 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9855_itm_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        butterFly2_15_conc_2_itm_9_2_1 <= STD_LOGIC_VECTOR'( "00");
      ELSIF ( butterFly1_15_conc_2_itm_9_0 = '1' ) THEN
        butterFly2_15_conc_2_itm_9_2_1 <= butterFly2_15_conc_2_itm_8_2_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( butterFly1_15_conc_2_itm_8_0 = '1' ) THEN
        reg_mult_47_res_lpi_3_dfm_1_cse <= mult_1_res_lpi_3_dfm_1_mx0;
        reg_mult_46_res_lpi_3_dfm_1_cse <= mult_9_res_lpi_3_dfm_1_mx0;
        reg_mult_45_res_lpi_3_dfm_1_cse <= mult_12_res_lpi_3_dfm_1_mx0;
        reg_mult_44_res_lpi_3_dfm_1_cse <= mult_4_res_lpi_3_dfm_1_mx0;
        reg_mult_43_res_lpi_3_dfm_1_cse <= mult_6_res_lpi_3_dfm_1_mx0;
        reg_mult_42_res_lpi_3_dfm_1_cse <= mult_14_res_lpi_3_dfm_1_mx0;
        reg_mult_41_res_lpi_3_dfm_1_cse <= mult_10_res_lpi_3_dfm_1_mx0;
        reg_mult_40_res_lpi_3_dfm_1_cse <= mult_2_res_lpi_3_dfm_1_mx0;
        reg_mult_39_res_lpi_3_dfm_1_cse <= mult_3_res_lpi_3_dfm_1_mx0;
        reg_mult_38_res_lpi_3_dfm_1_cse <= mult_7_res_lpi_3_dfm_1_mx0;
        reg_mult_37_res_lpi_3_dfm_1_cse <= mult_11_res_lpi_3_dfm_1_mx0;
        reg_mult_36_res_lpi_3_dfm_1_cse <= mult_15_res_lpi_3_dfm_1_mx0;
        reg_mult_35_res_lpi_3_dfm_1_cse <= mult_13_res_lpi_3_dfm_1_mx0;
        reg_mult_34_res_lpi_3_dfm_1_cse <= mult_8_res_lpi_3_dfm_1_mx0;
        reg_mult_33_res_lpi_3_dfm_1_cse <= mult_5_res_lpi_3_dfm_1_mx0;
        reg_mult_32_res_lpi_3_dfm_1_cse <= mult_res_lpi_3_dfm_1_mx0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        butterFly2_15_conc_2_itm_8_2_1 <= STD_LOGIC_VECTOR'( "00");
      ELSIF ( butterFly1_15_conc_2_itm_8_0 = '1' ) THEN
        butterFly2_15_conc_2_itm_8_2_1 <= butterFly2_15_conc_2_itm_7_2_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        butterFly2_15_conc_2_itm_7_2_1 <= STD_LOGIC_VECTOR'( "00");
      ELSIF ( butterFly1_15_conc_2_itm_7_0 = '1' ) THEN
        butterFly2_15_conc_2_itm_7_2_1 <= butterFly2_15_conc_2_itm_6_2_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( butterFly1_15_conc_2_itm_2_0 = '1' ) THEN
        tmp_126_lpi_3_dfm_1 <= z_out;
        tmp_124_lpi_3_dfm_1 <= z_out_1;
        tmp_122_lpi_3_dfm_1 <= z_out_2;
        tmp_120_lpi_3_dfm_1 <= z_out_3;
        tmp_118_lpi_3_dfm_1 <= z_out_4;
        tmp_116_lpi_3_dfm_1 <= z_out_5;
        tmp_114_lpi_3_dfm_1 <= z_out_6;
        tmp_112_lpi_3_dfm_1 <= z_out_7;
        tmp_110_lpi_3_dfm_1 <= z_out_8;
        tmp_108_lpi_3_dfm_1 <= z_out_9;
        tmp_106_lpi_3_dfm_1 <= z_out_10;
        tmp_104_lpi_3_dfm_1 <= z_out_11;
        tmp_102_lpi_3_dfm_1 <= z_out_12;
        tmp_100_lpi_3_dfm_1 <= z_out_13;
        tmp_98_lpi_3_dfm_1 <= z_out_14;
        tmp_96_lpi_3_dfm_1 <= z_out_15;
        tmp_62_lpi_3_dfm_1 <= z_out_16;
        tmp_60_lpi_3_dfm_1 <= z_out_17;
        tmp_58_lpi_3_dfm_1 <= z_out_18;
        tmp_56_lpi_3_dfm_1 <= z_out_19;
        tmp_54_lpi_3_dfm_1 <= z_out_20;
        tmp_52_lpi_3_dfm_1 <= z_out_21;
        tmp_50_lpi_3_dfm_1 <= z_out_22;
        tmp_48_lpi_3_dfm_1 <= z_out_23;
        tmp_46_lpi_3_dfm_1 <= z_out_24;
        tmp_44_lpi_3_dfm_1 <= z_out_25;
        tmp_42_lpi_3_dfm_1 <= z_out_26;
        tmp_40_lpi_3_dfm_1 <= z_out_27;
        tmp_38_lpi_3_dfm_1 <= z_out_28;
        tmp_36_lpi_3_dfm_1 <= z_out_29;
        tmp_34_lpi_3_dfm_1 <= z_out_30;
        tmp_32_lpi_3_dfm_1 <= z_out_31;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        operator_33_true_3_lshift_psp_1_0_sva <= STD_LOGIC_VECTOR'( "00");
      ELSIF ( (fsm_output(9)) = '0' ) THEN
        operator_33_true_3_lshift_psp_1_0_sva <= operator_33_true_3_lshift_psp_1_0_sva_mx0w5;
      END IF;
    END IF;
  END PROCESS;
  butterFly2_21_tw_butterFly2_21_tw_or_nl <= c_1_sva OR INNER_LOOP4_nor_tmp;
  c_mux_nl <= MUX_s_1_2_2((operator_20_false_acc_cse_sva(0)), butterFly2_21_tw_butterFly2_21_tw_or_nl,
      fsm_output(9));
  STAGE_LOOP_mux1h_nl <= MUX1HOT_v_2_6_2((INNER_LOOP1_r_INNER_LOOP1_r_and_cse(6 DOWNTO
      5)), (INNER_LOOP2_r_11_4_sva_6_0_mx1(6 DOWNTO 5)), (operator_20_false_acc_cse_sva(2
      DOWNTO 1)), (operator_33_true_2_lshift_psp_2_0_sva_mx0(1 DOWNTO 0)), operator_33_true_3_lshift_psp_1_0_sva_mx0w5,
      operator_33_true_3_lshift_psp_1_0_sva, STD_LOGIC_VECTOR'( or_tmp_3597 & or_dcpl_315
      & (fsm_output(5)) & or_tmp_3600 & (fsm_output(8)) & (fsm_output(9))));
  modulo_add_1_qif_mux1h_2_nl <= MUX1HOT_v_32_3_2(z_out_141, z_out_138, z_out_136,
      STD_LOGIC_VECTOR'( modulo_add_1_qelse_or_m1c & (fsm_output(7)) & (fsm_output(9))));
  acc_2_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_1_qif_mux1h_2_nl
      & '1') + UNSIGNED((NOT p_sva) & '1'), 33));
  modulo_add_1_qelse_and_nl <= (NOT z_out_143_32) AND modulo_add_1_qelse_or_m1c;
  modulo_add_1_qelse_or_1_nl <= (z_out_143_32 AND modulo_add_1_qelse_or_m1c) OR (z_out_143_32
      AND (fsm_output(7))) OR (z_out_145_32 AND (fsm_output(9)));
  modulo_add_1_qelse_and_4_nl <= (NOT z_out_143_32) AND (fsm_output(7));
  modulo_add_1_qelse_and_5_nl <= (NOT z_out_145_32) AND (fsm_output(9));
  modulo_add_10_qif_mux1h_2_nl <= MUX1HOT_v_32_4_2(z_out_132, z_out_127, z_out_128,
      z_out_142, STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7))
      & (fsm_output(9))));
  acc_3_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_10_qif_mux1h_2_nl
      & '1') + UNSIGNED((NOT p_sva) & '1'), 33));
  modulo_add_10_qelse_and_nl <= (NOT z_out_144_32) AND (fsm_output(2));
  modulo_add_10_qelse_or_nl <= (z_out_144_32 AND (fsm_output(2))) OR (z_out_144_32
      AND (fsm_output(4))) OR (z_out_144_32 AND (fsm_output(7))) OR (z_out_146_32
      AND (fsm_output(9)));
  modulo_add_10_qelse_and_5_nl <= (NOT z_out_144_32) AND (fsm_output(4));
  modulo_add_10_qelse_and_6_nl <= (NOT z_out_144_32) AND (fsm_output(7));
  modulo_add_10_qelse_and_7_nl <= (NOT z_out_146_32) AND (fsm_output(9));
  modulo_add_11_qif_mux1h_2_nl <= MUX1HOT_v_32_4_2(z_out_131, z_out_137, z_out_127,
      z_out_141, STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7))
      & (fsm_output(9))));
  acc_4_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_11_qif_mux1h_2_nl
      & '1') + UNSIGNED((NOT p_sva) & '1'), 33));
  modulo_add_11_qelse_and_nl <= (NOT z_out_146_32) AND (fsm_output(2));
  modulo_add_11_qelse_or_nl <= (z_out_146_32 AND (fsm_output(2))) OR (z_out_146_32
      AND (fsm_output(4))) OR (z_out_147_32 AND (fsm_output(7))) OR (z_out_147_32
      AND (fsm_output(9)));
  modulo_add_11_qelse_and_5_nl <= (NOT z_out_146_32) AND (fsm_output(4));
  modulo_add_11_qelse_and_6_nl <= (NOT z_out_147_32) AND (fsm_output(7));
  modulo_add_11_qelse_and_7_nl <= (NOT z_out_147_32) AND (fsm_output(9));
  modulo_add_12_qif_mux1h_2_nl <= MUX1HOT_v_32_3_2(z_out_130, z_out_142, z_out_140,
      STD_LOGIC_VECTOR'( modulo_add_1_qelse_or_m1c & (fsm_output(7)) & (fsm_output(9))));
  acc_5_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_12_qif_mux1h_2_nl
      & '1') + UNSIGNED((NOT p_sva) & '1'), 33));
  modulo_add_12_qelse_and_nl <= (NOT z_out_147_32) AND modulo_add_1_qelse_or_m1c;
  modulo_add_12_qelse_or_1_nl <= (z_out_147_32 AND modulo_add_1_qelse_or_m1c) OR
      (z_out_148_32 AND (fsm_output(7))) OR (z_out_150_32 AND (fsm_output(9)));
  modulo_add_12_qelse_and_4_nl <= (NOT z_out_148_32) AND (fsm_output(7));
  modulo_add_12_qelse_and_5_nl <= (NOT z_out_150_32) AND (fsm_output(9));
  modulo_add_13_qif_mux1h_2_nl <= MUX1HOT_v_32_3_2(z_out_129, z_out_141, z_out_139,
      STD_LOGIC_VECTOR'( modulo_add_1_qelse_or_m1c & (fsm_output(7)) & (fsm_output(9))));
  acc_6_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_13_qif_mux1h_2_nl
      & '1') + UNSIGNED((NOT p_sva) & '1'), 33));
  modulo_add_13_qelse_and_nl <= (NOT z_out_150_32) AND modulo_add_1_qelse_or_m1c;
  modulo_add_13_qelse_or_1_nl <= (z_out_150_32 AND modulo_add_1_qelse_or_m1c) OR
      (z_out_150_32 AND (fsm_output(7))) OR (z_out_151_32 AND (fsm_output(9)));
  modulo_add_13_qelse_and_4_nl <= (NOT z_out_150_32) AND (fsm_output(7));
  modulo_add_13_qelse_and_5_nl <= (NOT z_out_151_32) AND (fsm_output(9));
  modulo_add_14_qif_mux1h_2_nl <= MUX1HOT_v_32_3_2(z_out_128, z_out_140, z_out_138,
      STD_LOGIC_VECTOR'( modulo_add_1_qelse_or_m1c & (fsm_output(7)) & (fsm_output(9))));
  acc_10_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_14_qif_mux1h_2_nl
      & '1') + UNSIGNED((NOT p_sva) & '1'), 33));
  modulo_add_14_qelse_and_nl <= (NOT z_out_152_32) AND modulo_add_1_qelse_or_m1c;
  modulo_add_14_qelse_or_1_nl <= (z_out_152_32 AND modulo_add_1_qelse_or_m1c) OR
      (z_out_153_32 AND (fsm_output(7))) OR (z_out_154_32 AND (fsm_output(9)));
  modulo_add_14_qelse_and_4_nl <= (NOT z_out_153_32) AND (fsm_output(7));
  modulo_add_14_qelse_and_5_nl <= (NOT z_out_154_32) AND (fsm_output(9));
  modulo_add_15_qif_mux1h_2_nl <= MUX1HOT_v_32_4_2(z_out_127, z_out_142, z_out_139,
      z_out_137, STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7))
      & (fsm_output(9))));
  acc_14_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_15_qif_mux1h_2_nl
      & '1') + UNSIGNED((NOT p_sva) & '1'), 33));
  modulo_add_15_qelse_and_nl <= (NOT z_out_153_32) AND (fsm_output(2));
  modulo_add_15_qelse_or_nl <= (z_out_153_32 AND (fsm_output(2))) OR (z_out_153_32
      AND (fsm_output(4))) OR (z_out_154_32 AND (fsm_output(7))) OR (z_out_157_32
      AND (fsm_output(9)));
  modulo_add_15_qelse_and_5_nl <= (NOT z_out_153_32) AND (fsm_output(4));
  modulo_add_15_qelse_and_6_nl <= (NOT z_out_154_32) AND (fsm_output(7));
  modulo_add_15_qelse_and_7_nl <= (NOT z_out_157_32) AND (fsm_output(9));
  butterFly1_f1_butterFly1_f1_nor_nl <= NOT(CONV_SL_1_1(INNER_LOOP1_r_11_4_sva_6_0(6
      DOWNTO 4)/=STD_LOGIC_VECTOR'("000")));
  butterFly1_16_f1_butterFly1_16_f1_nor_nl <= NOT(CONV_SL_1_1(INNER_LOOP2_r_11_4_sva_6_0(6
      DOWNTO 4)/=STD_LOGIC_VECTOR'("000")));
  butterFly2_f1_butterFly2_f1_and_5_nl <= CONV_SL_1_1(INNER_LOOP3_r_11_4_sva_6_0(6
      DOWNTO 4)=STD_LOGIC_VECTOR'("110"));
  butterFly2_16_f1_butterFly2_16_f1_and_5_nl <= CONV_SL_1_1(INNER_LOOP4_r_11_4_sva_6_0(6
      DOWNTO 4)=STD_LOGIC_VECTOR'("110"));
  butterFly1_f1_butterFly1_f1_and_nl <= (INNER_LOOP1_r_11_4_sva_6_0(4)) AND butterFly1_f1_nor_cse;
  butterFly1_16_f1_butterFly1_16_f1_and_nl <= CONV_SL_1_1(INNER_LOOP2_r_11_4_sva_6_0(6
      DOWNTO 4)=STD_LOGIC_VECTOR'("001"));
  butterFly1_f1_butterFly1_f1_and_1_nl <= CONV_SL_1_1(INNER_LOOP1_r_11_4_sva_6_0(6
      DOWNTO 4)=STD_LOGIC_VECTOR'("010"));
  butterFly1_16_f1_butterFly1_16_f1_and_1_nl <= CONV_SL_1_1(INNER_LOOP2_r_11_4_sva_6_0(6
      DOWNTO 4)=STD_LOGIC_VECTOR'("010"));
  butterFly1_f1_butterFly1_f1_and_2_nl <= CONV_SL_1_1(INNER_LOOP1_r_11_4_sva_6_0(6
      DOWNTO 4)=STD_LOGIC_VECTOR'("011"));
  butterFly1_16_f1_butterFly1_16_f1_and_2_nl <= CONV_SL_1_1(INNER_LOOP2_r_11_4_sva_6_0(6
      DOWNTO 4)=STD_LOGIC_VECTOR'("011"));
  butterFly2_f1_butterFly2_f1_and_nl <= (INNER_LOOP3_r_11_4_sva_6_0(4)) AND butterFly2_f1_nor_cse;
  butterFly2_16_f1_butterFly2_16_f1_and_nl <= CONV_SL_1_1(INNER_LOOP4_r_11_4_sva_6_0(6
      DOWNTO 4)=STD_LOGIC_VECTOR'("001"));
  butterFly1_f1_butterFly1_f1_and_3_nl <= CONV_SL_1_1(INNER_LOOP1_r_11_4_sva_6_0(6
      DOWNTO 4)=STD_LOGIC_VECTOR'("100"));
  butterFly1_16_f1_butterFly1_16_f1_and_3_nl <= CONV_SL_1_1(INNER_LOOP2_r_11_4_sva_6_0(6
      DOWNTO 4)=STD_LOGIC_VECTOR'("100"));
  butterFly2_f1_butterFly2_f1_and_1_nl <= CONV_SL_1_1(INNER_LOOP3_r_11_4_sva_6_0(6
      DOWNTO 4)=STD_LOGIC_VECTOR'("010"));
  butterFly2_16_f1_butterFly2_16_f1_and_1_nl <= (INNER_LOOP4_r_11_4_sva_6_0(5)) AND
      butterFly2_16_f1_nor_1_cse;
  butterFly1_f1_butterFly1_f1_and_4_nl <= CONV_SL_1_1(INNER_LOOP1_r_11_4_sva_6_0(6
      DOWNTO 4)=STD_LOGIC_VECTOR'("101"));
  butterFly1_16_f1_butterFly1_16_f1_and_4_nl <= CONV_SL_1_1(INNER_LOOP2_r_11_4_sva_6_0(6
      DOWNTO 4)=STD_LOGIC_VECTOR'("101"));
  butterFly2_f1_butterFly2_f1_and_2_nl <= CONV_SL_1_1(INNER_LOOP3_r_11_4_sva_6_0(6
      DOWNTO 4)=STD_LOGIC_VECTOR'("011"));
  butterFly2_16_f1_butterFly2_16_f1_and_2_nl <= CONV_SL_1_1(INNER_LOOP4_r_11_4_sva_6_0(6
      DOWNTO 4)=STD_LOGIC_VECTOR'("011"));
  butterFly1_f1_butterFly1_f1_and_5_nl <= CONV_SL_1_1(INNER_LOOP1_r_11_4_sva_6_0(6
      DOWNTO 4)=STD_LOGIC_VECTOR'("110"));
  butterFly1_16_f1_butterFly1_16_f1_and_5_nl <= CONV_SL_1_1(INNER_LOOP2_r_11_4_sva_6_0(6
      DOWNTO 4)=STD_LOGIC_VECTOR'("110"));
  butterFly2_f1_butterFly2_f1_and_3_nl <= CONV_SL_1_1(INNER_LOOP3_r_11_4_sva_6_0(6
      DOWNTO 4)=STD_LOGIC_VECTOR'("100"));
  butterFly2_16_f1_butterFly2_16_f1_and_3_nl <= CONV_SL_1_1(INNER_LOOP4_r_11_4_sva_6_0(6
      DOWNTO 4)=STD_LOGIC_VECTOR'("100"));
  butterFly1_f1_butterFly1_f1_and_6_nl <= CONV_SL_1_1(INNER_LOOP1_r_11_4_sva_6_0(6
      DOWNTO 4)=STD_LOGIC_VECTOR'("111"));
  butterFly1_16_f1_butterFly1_16_f1_and_6_nl <= CONV_SL_1_1(INNER_LOOP2_r_11_4_sva_6_0(6
      DOWNTO 4)=STD_LOGIC_VECTOR'("111"));
  butterFly2_f1_butterFly2_f1_and_4_nl <= CONV_SL_1_1(INNER_LOOP3_r_11_4_sva_6_0(6
      DOWNTO 4)=STD_LOGIC_VECTOR'("101"));
  butterFly2_16_f1_butterFly2_16_f1_and_4_nl <= CONV_SL_1_1(INNER_LOOP4_r_11_4_sva_6_0(6
      DOWNTO 4)=STD_LOGIC_VECTOR'("101"));
  INNER_LOOP1_mux_nl <= MUX_s_1_2_2(INNER_LOOP1_stage_0, INNER_LOOP1_stage_0_10,
      fsm_output(7));
  INNER_LOOP1_mux_4_nl <= MUX_s_1_2_2(INNER_LOOP1_stage_0_2, INNER_LOOP1_stage_0_11,
      fsm_output(7));
  INNER_LOOP1_mux_5_nl <= MUX_s_1_2_2(butterFly2_15_conc_2_itm_5_0, (operator_33_true_2_lshift_psp_2_0_sva_mx0(0)),
      or_tmp_3600);
  INNER_LOOP1_mux_6_nl <= MUX_s_1_2_2(INNER_LOOP1_stage_0_10, (operator_33_true_2_lshift_psp_2_0_sva_mx0(2)),
      or_tmp_3600);
  butterFly1_15_mux_9_nl <= MUX_s_1_2_2(butterFly1_15_conc_2_itm_1_0, INNER_LOOP1_stage_0,
      or_dcpl_298);
  butterFly1_15_mux1h_47_nl <= MUX1HOT_s_1_3_2((INNER_LOOP1_r_INNER_LOOP1_r_and_cse(0)),
      (INNER_LOOP2_r_11_4_sva_6_0_mx1(0)), butterFly1_15_conc_2_itm_9_0, STD_LOGIC_VECTOR'(
      or_tmp_3597 & or_dcpl_315 & or_dcpl_298));
  butterFly2_15_mux1h_3_nl <= MUX1HOT_s_1_4_2(INNER_LOOP1_stage_0_3, butterFly2_15_conc_2_itm_8_0,
      (INNER_LOOP1_r_INNER_LOOP1_r_and_3_cse(0)), (INNER_LOOP1_r_INNER_LOOP1_r_and_5_cse(0)),
      STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & or_tmp_3600 & or_tmp_3732));
  butterFly1_15_mux_10_nl <= MUX_s_1_2_2(butterFly1_15_conc_2_itm_9_0, butterFly2_15_conc_2_itm_5_0,
      or_tmp_3842);
  modulo_add_2_qif_mux1h_2_nl <= MUX1HOT_v_32_3_2(z_out_140, z_out_137, z_out_135,
      STD_LOGIC_VECTOR'( modulo_add_1_qelse_or_m1c & (fsm_output(7)) & (fsm_output(9))));
  acc_18_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_2_qif_mux1h_2_nl
      & '1') + UNSIGNED((NOT p_sva) & '1'), 33));
  modulo_add_23_qelse_and_nl <= (NOT z_out_156_32) AND modulo_add_1_qelse_or_m1c;
  modulo_add_23_qelse_or_1_nl <= (z_out_156_32 AND modulo_add_1_qelse_or_m1c) OR
      (z_out_156_32 AND (fsm_output(7))) OR (z_out_158_32 AND (fsm_output(9)));
  modulo_add_23_qelse_and_4_nl <= (NOT z_out_156_32) AND (fsm_output(7));
  modulo_add_23_qelse_and_5_nl <= (NOT z_out_158_32) AND (fsm_output(9));
  modulo_add_3_qif_mux1h_2_nl <= MUX1HOT_v_32_3_2(z_out_139, z_out_136, z_out_134,
      STD_LOGIC_VECTOR'( modulo_add_1_qelse_or_m1c & (fsm_output(7)) & (fsm_output(9))));
  acc_22_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_3_qif_mux1h_2_nl
      & '1') + UNSIGNED((NOT p_sva) & '1'), 33));
  modulo_add_24_qelse_and_nl <= (NOT z_out_158_32) AND modulo_add_1_qelse_or_m1c;
  modulo_add_24_qelse_or_1_nl <= (z_out_158_32 AND modulo_add_1_qelse_or_m1c) OR
      (z_out_157_32 AND (fsm_output(7))) OR (z_out_156_32 AND (fsm_output(9)));
  modulo_add_24_qelse_and_4_nl <= (NOT z_out_157_32) AND (fsm_output(7));
  modulo_add_24_qelse_and_5_nl <= (NOT z_out_156_32) AND (fsm_output(9));
  modulo_add_4_qif_mux1h_2_nl <= MUX1HOT_v_32_3_2(z_out_138, z_out_135, z_out_133,
      STD_LOGIC_VECTOR'( modulo_add_1_qelse_or_m1c & (fsm_output(7)) & (fsm_output(9))));
  acc_26_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_4_qif_mux1h_2_nl
      & '1') + UNSIGNED((NOT p_sva) & '1'), 33));
  modulo_add_25_qelse_and_nl <= (NOT z_out_157_32) AND modulo_add_1_qelse_or_m1c;
  modulo_add_25_qelse_or_1_nl <= (z_out_157_32 AND modulo_add_1_qelse_or_m1c) OR
      (z_out_155_32 AND (fsm_output(7))) OR (z_out_152_32 AND (fsm_output(9)));
  modulo_add_25_qelse_and_4_nl <= (NOT z_out_155_32) AND (fsm_output(7));
  modulo_add_25_qelse_and_5_nl <= (NOT z_out_152_32) AND (fsm_output(9));
  modulo_add_5_qif_mux1h_2_nl <= MUX1HOT_v_32_4_2(z_out_137, z_out_136, z_out_134,
      z_out_132, STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7))
      & (fsm_output(9))));
  acc_30_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_5_qif_mux1h_2_nl
      & '1') + UNSIGNED((NOT p_sva) & '1'), 33));
  modulo_add_26_qelse_and_nl <= (NOT z_out_151_32) AND (fsm_output(2));
  modulo_add_26_qelse_or_nl <= (z_out_151_32 AND (fsm_output(2))) OR (z_out_151_32
      AND (fsm_output(4))) OR (z_out_151_32 AND (fsm_output(7))) OR (z_out_148_32
      AND (fsm_output(9)));
  modulo_add_26_qelse_and_5_nl <= (NOT z_out_151_32) AND (fsm_output(4));
  modulo_add_26_qelse_and_6_nl <= (NOT z_out_151_32) AND (fsm_output(7));
  modulo_add_26_qelse_and_7_nl <= (NOT z_out_148_32) AND (fsm_output(9));
  modulo_add_6_qif_mux1h_2_nl <= MUX1HOT_v_32_4_2(z_out_136, z_out_135, z_out_133,
      z_out_131, STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7))
      & (fsm_output(9))));
  acc_34_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_6_qif_mux1h_2_nl
      & '1') + UNSIGNED((NOT p_sva) & '1'), 33));
  modulo_add_27_qelse_and_nl <= (NOT z_out_149_32) AND (fsm_output(2));
  modulo_add_27_qelse_or_nl <= (z_out_149_32 AND (fsm_output(2))) OR (z_out_149_32
      AND (fsm_output(4))) OR (z_out_145_32 AND (fsm_output(7))) OR (z_out_144_32
      AND (fsm_output(9)));
  modulo_add_27_qelse_and_5_nl <= (NOT z_out_149_32) AND (fsm_output(4));
  modulo_add_27_qelse_and_6_nl <= (NOT z_out_145_32) AND (fsm_output(7));
  modulo_add_27_qelse_and_7_nl <= (NOT z_out_144_32) AND (fsm_output(9));
  modulo_add_7_qif_mux1h_2_nl <= MUX1HOT_v_32_4_2(z_out_135, z_out_134, z_out_132,
      z_out_130, STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7))
      & (fsm_output(9))));
  acc_38_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_7_qif_mux1h_2_nl
      & '1') + UNSIGNED((NOT p_sva) & '1'), 33));
  modulo_add_28_qelse_and_nl <= (NOT z_out_145_32) AND (fsm_output(2));
  modulo_add_28_qelse_or_nl <= (z_out_145_32 AND (fsm_output(2))) OR (z_out_145_32
      AND (fsm_output(4))) OR (z_out_149_32 AND (fsm_output(7))) OR (z_out_153_32
      AND (fsm_output(9)));
  modulo_add_28_qelse_and_5_nl <= (NOT z_out_145_32) AND (fsm_output(4));
  modulo_add_28_qelse_and_6_nl <= (NOT z_out_149_32) AND (fsm_output(7));
  modulo_add_28_qelse_and_7_nl <= (NOT z_out_153_32) AND (fsm_output(9));
  modulo_add_8_qif_mux1h_2_nl <= MUX1HOT_v_32_4_2(z_out_134, z_out_133, z_out_131,
      z_out_129, STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7))
      & (fsm_output(9))));
  acc_42_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_8_qif_mux1h_2_nl
      & '1') + UNSIGNED((NOT p_sva) & '1'), 33));
  modulo_add_29_qelse_and_nl <= (NOT z_out_155_32) AND (fsm_output(2));
  modulo_add_29_qelse_or_nl <= (z_out_155_32 AND (fsm_output(2))) OR (z_out_155_32
      AND (fsm_output(4))) OR (z_out_158_32 AND (fsm_output(7))) OR (z_out_155_32
      AND (fsm_output(9)));
  modulo_add_29_qelse_and_5_nl <= (NOT z_out_155_32) AND (fsm_output(4));
  modulo_add_29_qelse_and_6_nl <= (NOT z_out_158_32) AND (fsm_output(7));
  modulo_add_29_qelse_and_7_nl <= (NOT z_out_155_32) AND (fsm_output(9));
  modulo_add_9_qif_mux1h_2_nl <= MUX1HOT_v_32_4_2(z_out_133, z_out_132, z_out_130,
      z_out_128, STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7))
      & (fsm_output(9))));
  acc_46_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_9_qif_mux1h_2_nl
      & '1') + UNSIGNED((NOT p_sva) & '1'), 33));
  modulo_add_30_qelse_and_nl <= (NOT z_out_154_32) AND (fsm_output(2));
  modulo_add_30_qelse_or_nl <= (z_out_154_32 AND (fsm_output(2))) OR (z_out_154_32
      AND (fsm_output(4))) OR (z_out_152_32 AND (fsm_output(7))) OR (z_out_149_32
      AND (fsm_output(9)));
  modulo_add_30_qelse_and_5_nl <= (NOT z_out_154_32) AND (fsm_output(4));
  modulo_add_30_qelse_and_6_nl <= (NOT z_out_152_32) AND (fsm_output(7));
  modulo_add_30_qelse_and_7_nl <= (NOT z_out_149_32) AND (fsm_output(9));
  modulo_add_qif_mux1h_2_nl <= MUX1HOT_v_32_4_2(z_out_142, z_out_131, z_out_129,
      z_out_127, STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7))
      & (fsm_output(9))));
  acc_49_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_qif_mux1h_2_nl
      & '1') + UNSIGNED((NOT p_sva) & '1'), 33));
  modulo_add_31_qelse_and_nl <= (NOT z_out_148_32) AND (fsm_output(2));
  modulo_add_31_qelse_or_nl <= (z_out_148_32 AND (fsm_output(2))) OR (z_out_148_32
      AND (fsm_output(4))) OR (z_out_146_32 AND (fsm_output(7))) OR (z_out_143_32
      AND (fsm_output(9)));
  modulo_add_31_qelse_and_5_nl <= (NOT z_out_148_32) AND (fsm_output(4));
  modulo_add_31_qelse_and_6_nl <= (NOT z_out_146_32) AND (fsm_output(7));
  modulo_add_31_qelse_and_7_nl <= (NOT z_out_143_32) AND (fsm_output(9));
  modulo_sub_16_qelse_or_nl <= ((z_out_126(31)) AND (NOT (fsm_output(9)))) OR ((z_out_111(31))
      AND (fsm_output(9)));
  modulo_sub_17_qelse_or_nl <= ((z_out_116(31)) AND (NOT (fsm_output(9)))) OR ((z_out_112(31))
      AND (fsm_output(9)));
  modulo_sub_18_qelse_or_nl <= ((z_out_123(31)) AND (NOT (fsm_output(9)))) OR ((z_out_113(31))
      AND (fsm_output(9)));
  modulo_sub_19_qelse_or_nl <= ((z_out_124(31)) AND (NOT (fsm_output(9)))) OR ((z_out_114(31))
      AND (fsm_output(9)));
  modulo_sub_20_qelse_or_nl <= ((z_out_125(31)) AND (NOT (fsm_output(9)))) OR ((z_out_115(31))
      AND (fsm_output(9)));
  modulo_sub_21_qelse_or_nl <= ((z_out_111(31)) AND (NOT (fsm_output(9)))) OR ((z_out_116(31))
      AND (fsm_output(9)));
  modulo_sub_22_qelse_or_nl <= ((z_out_112(31)) AND (NOT (fsm_output(9)))) OR ((z_out_117(31))
      AND (fsm_output(9)));
  modulo_sub_23_qelse_or_nl <= ((z_out_113(31)) AND (NOT (fsm_output(9)))) OR ((z_out_118(31))
      AND (fsm_output(9)));
  modulo_sub_24_qelse_or_nl <= ((z_out_114(31)) AND (NOT (fsm_output(9)))) OR ((z_out_119(31))
      AND (fsm_output(9)));
  modulo_sub_25_qelse_or_nl <= ((z_out_115(31)) AND (NOT (fsm_output(9)))) OR ((z_out_120(31))
      AND (fsm_output(9)));
  modulo_sub_26_qelse_or_nl <= ((z_out_117(31)) AND (NOT (fsm_output(9)))) OR ((z_out_121(31))
      AND (fsm_output(9)));
  modulo_sub_27_qelse_or_nl <= ((z_out_118(31)) AND (NOT (fsm_output(9)))) OR ((z_out_122(31))
      AND (fsm_output(9)));
  modulo_sub_28_qelse_or_nl <= ((z_out_119(31)) AND (NOT (fsm_output(9)))) OR ((z_out_123(31))
      AND (fsm_output(9)));
  modulo_sub_29_qelse_or_nl <= ((z_out_120(31)) AND (NOT (fsm_output(9)))) OR ((z_out_124(31))
      AND (fsm_output(9)));
  modulo_sub_30_qelse_or_nl <= ((z_out_121(31)) AND (NOT (fsm_output(9)))) OR ((z_out_125(31))
      AND (fsm_output(9)));
  modulo_sub_31_qelse_or_nl <= ((z_out_122(31)) AND (NOT (fsm_output(9)))) OR ((z_out_126(31))
      AND (fsm_output(9)));
  INNER_LOOP1_mux_7_nl <= MUX_s_1_2_2(INNER_LOOP1_stage_0, INNER_LOOP2_stage_0_10,
      or_dcpl_298);
  butterFly2_f1_butterFly2_f1_nor_nl <= NOT(CONV_SL_1_1(INNER_LOOP3_r_11_4_sva_6_0(6
      DOWNTO 4)/=STD_LOGIC_VECTOR'("000")));
  butterFly2_16_f1_butterFly2_16_f1_nor_nl <= NOT(CONV_SL_1_1(INNER_LOOP4_r_11_4_sva_6_0(6
      DOWNTO 4)/=STD_LOGIC_VECTOR'("000")));
  butterFly2_f1_butterFly2_f1_and_6_nl <= CONV_SL_1_1(INNER_LOOP3_r_11_4_sva_6_0(6
      DOWNTO 4)=STD_LOGIC_VECTOR'("111"));
  STAGE_LOOP_base_STAGE_LOOP_base_mux_nl <= MUX_v_7_2_2((z_out_60(10 DOWNTO 4)),
      (z_out_62(6 DOWNTO 0)), fsm_output(4));
  INNER_LOOP2_r_or_nl <= (fsm_output(1)) OR (fsm_output(4)) OR (fsm_output(2));
  operator_20_false_mux_2_nl <= MUX_v_3_2_2((butterFly1_15_conc_2_itm_2_1 & c_1_sva),
      operator_20_false_acc_cse_sva, fsm_output(5));
  z_out_61 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(operator_20_false_mux_2_nl)
      + UNSIGNED'( '1' & (NOT (fsm_output(5))) & '1'), 3));
  operator_20_false_mux1h_2_nl <= MUX1HOT_v_7_4_2(INNER_LOOP1_r_11_4_sva_6_0, INNER_LOOP2_r_11_4_sva_6_0,
      INNER_LOOP3_r_11_4_sva_6_0, INNER_LOOP4_r_11_4_sva_6_0, STD_LOGIC_VECTOR'(
      (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  z_out_62 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(operator_20_false_mux1h_2_nl),
      8) + UNSIGNED'( "00000001"), 8));
  modulo_sub_15_qif_mux_2_nl <= MUX_v_31_2_2((z_out_126(30 DOWNTO 0)), (z_out_124(30
      DOWNTO 0)), fsm_output(7));
  z_out_68 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_15_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_31_qif_mux_2_nl <= MUX_v_31_2_2((z_out_122(30 DOWNTO 0)), (z_out_126(30
      DOWNTO 0)), fsm_output(9));
  z_out_69 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_31_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_7_qif_mux_2_nl <= MUX_v_31_2_2((z_out_118(30 DOWNTO 0)), (z_out_123(30
      DOWNTO 0)), fsm_output(7));
  z_out_70 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_7_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_30_qif_mux_2_nl <= MUX_v_31_2_2((z_out_121(30 DOWNTO 0)), (z_out_125(30
      DOWNTO 0)), fsm_output(9));
  z_out_72 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_30_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_39_qif_mux_2_nl <= MUX_v_31_2_2((z_out_116(30 DOWNTO 0)), (z_out_125(30
      DOWNTO 0)), fsm_output(2));
  z_out_73 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_39_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_29_qif_mux_2_nl <= MUX_v_31_2_2((z_out_120(30 DOWNTO 0)), (z_out_124(30
      DOWNTO 0)), fsm_output(9));
  z_out_74 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_29_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_6_qif_mux_2_nl <= MUX_v_31_2_2((z_out_117(30 DOWNTO 0)), (z_out_122(30
      DOWNTO 0)), fsm_output(7));
  z_out_76 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_6_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_28_qif_mux_2_nl <= MUX_v_31_2_2((z_out_119(30 DOWNTO 0)), (z_out_123(30
      DOWNTO 0)), fsm_output(9));
  z_out_77 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_28_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_38_qif_mux_2_nl <= MUX_v_31_2_2((z_out_115(30 DOWNTO 0)), (z_out_124(30
      DOWNTO 0)), fsm_output(2));
  z_out_78 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_38_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_27_qif_mux_2_nl <= MUX_v_31_2_2((z_out_118(30 DOWNTO 0)), (z_out_122(30
      DOWNTO 0)), fsm_output(9));
  z_out_80 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_27_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_5_qif_mux_2_nl <= MUX_v_31_2_2((z_out_116(30 DOWNTO 0)), (z_out_121(30
      DOWNTO 0)), fsm_output(7));
  z_out_81 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_5_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_26_qif_mux_2_nl <= MUX_v_31_2_2((z_out_117(30 DOWNTO 0)), (z_out_121(30
      DOWNTO 0)), fsm_output(9));
  z_out_82 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_26_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_37_qif_mux_2_nl <= MUX_v_31_2_2((z_out_114(30 DOWNTO 0)), (z_out_123(30
      DOWNTO 0)), fsm_output(2));
  z_out_84 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_37_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_25_qif_mux_2_nl <= MUX_v_31_2_2((z_out_115(30 DOWNTO 0)), (z_out_120(30
      DOWNTO 0)), fsm_output(9));
  z_out_85 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_25_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_4_qif_mux_2_nl <= MUX_v_31_2_2((z_out_115(30 DOWNTO 0)), (z_out_120(30
      DOWNTO 0)), fsm_output(7));
  z_out_86 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_4_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_24_qif_mux_2_nl <= MUX_v_31_2_2((z_out_114(30 DOWNTO 0)), (z_out_119(30
      DOWNTO 0)), fsm_output(9));
  z_out_88 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_24_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_36_qif_mux_2_nl <= MUX_v_31_2_2((z_out_113(30 DOWNTO 0)), (z_out_122(30
      DOWNTO 0)), fsm_output(2));
  z_out_89 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_36_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_23_qif_mux_2_nl <= MUX_v_31_2_2((z_out_113(30 DOWNTO 0)), (z_out_118(30
      DOWNTO 0)), fsm_output(9));
  z_out_90 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_23_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_3_qif_mux_2_nl <= MUX_v_31_2_2((z_out_114(30 DOWNTO 0)), (z_out_119(30
      DOWNTO 0)), fsm_output(7));
  z_out_92 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_3_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_22_qif_mux_2_nl <= MUX_v_31_2_2((z_out_112(30 DOWNTO 0)), (z_out_117(30
      DOWNTO 0)), fsm_output(9));
  z_out_93 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_22_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_35_qif_mux_2_nl <= MUX_v_31_2_2((z_out_112(30 DOWNTO 0)), (z_out_121(30
      DOWNTO 0)), fsm_output(2));
  z_out_94 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_35_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_21_qif_mux_2_nl <= MUX_v_31_2_2((z_out_111(30 DOWNTO 0)), (z_out_116(30
      DOWNTO 0)), fsm_output(9));
  z_out_96 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_21_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_2_qif_mux_2_nl <= MUX_v_31_2_2((z_out_113(30 DOWNTO 0)), (z_out_118(30
      DOWNTO 0)), fsm_output(7));
  z_out_97 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_2_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_20_qif_mux_2_nl <= MUX_v_31_2_2((z_out_125(30 DOWNTO 0)), (z_out_115(30
      DOWNTO 0)), fsm_output(9));
  z_out_98 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_20_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_34_qif_mux_2_nl <= MUX_v_31_2_2((z_out_111(30 DOWNTO 0)), (z_out_120(30
      DOWNTO 0)), fsm_output(2));
  z_out_100 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_34_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_19_qif_mux_2_nl <= MUX_v_31_2_2((z_out_124(30 DOWNTO 0)), (z_out_114(30
      DOWNTO 0)), fsm_output(9));
  z_out_101 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_19_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_1_qif_mux_2_nl <= MUX_v_31_2_2((z_out_112(30 DOWNTO 0)), (z_out_117(30
      DOWNTO 0)), fsm_output(7));
  z_out_102 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_1_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_18_qif_mux_2_nl <= MUX_v_31_2_2((z_out_123(30 DOWNTO 0)), (z_out_113(30
      DOWNTO 0)), fsm_output(9));
  z_out_104 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_18_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_33_qif_mux_2_nl <= MUX_v_31_2_2((z_out_126(30 DOWNTO 0)), (z_out_119(30
      DOWNTO 0)), fsm_output(2));
  z_out_105 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_33_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_17_qif_mux_2_nl <= MUX_v_31_2_2((z_out_116(30 DOWNTO 0)), (z_out_112(30
      DOWNTO 0)), fsm_output(9));
  z_out_106 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_17_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_qif_mux_2_nl <= MUX_v_31_2_2((z_out_111(30 DOWNTO 0)), (z_out_125(30
      DOWNTO 0)), fsm_output(7));
  z_out_108 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_16_qif_mux_2_nl <= MUX_v_31_2_2((z_out_126(30 DOWNTO 0)), (z_out_111(30
      DOWNTO 0)), fsm_output(9));
  z_out_109 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_16_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  butterFly1_mux1h_18_nl <= MUX1HOT_v_32_4_2((NOT reg_mult_res_lpi_3_dfm_1_cse),
      (NOT reg_mult_5_res_lpi_3_dfm_1_cse), (NOT reg_mult_34_res_lpi_3_dfm_1_cse),
      (NOT reg_mult_47_res_lpi_3_dfm_1_cse), STD_LOGIC_VECTOR'( (fsm_output(2)) &
      (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  acc_50_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_10_lpi_3_dfm_7 & '1')
      + UNSIGNED(butterFly1_mux1h_18_nl & '1'), 33));
  z_out_111 <= acc_50_nl(32 DOWNTO 1);
  butterFly1_1_mux1h_18_nl <= MUX1HOT_v_32_4_2((NOT reg_mult_1_res_lpi_3_dfm_1_cse),
      (NOT reg_mult_6_res_lpi_3_dfm_1_cse), (NOT reg_mult_35_res_lpi_3_dfm_1_cse),
      (NOT reg_mult_46_res_lpi_3_dfm_1_cse), STD_LOGIC_VECTOR'( (fsm_output(2)) &
      (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  acc_51_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_102_lpi_3_dfm_7 & '1')
      + UNSIGNED(butterFly1_1_mux1h_18_nl & '1'), 33));
  z_out_112 <= acc_51_nl(32 DOWNTO 1);
  butterFly1_2_mux1h_18_nl <= MUX1HOT_v_32_4_2((NOT reg_mult_2_res_lpi_3_dfm_1_cse),
      (NOT reg_mult_7_res_lpi_3_dfm_1_cse), (NOT reg_mult_36_res_lpi_3_dfm_1_cse),
      (NOT reg_mult_45_res_lpi_3_dfm_1_cse), STD_LOGIC_VECTOR'( (fsm_output(2)) &
      (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  acc_52_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_104_lpi_3_dfm_7 & '1')
      + UNSIGNED(butterFly1_2_mux1h_18_nl & '1'), 33));
  z_out_113 <= acc_52_nl(32 DOWNTO 1);
  butterFly1_3_mux1h_18_nl <= MUX1HOT_v_32_4_2((NOT reg_mult_3_res_lpi_3_dfm_1_cse),
      (NOT reg_mult_8_res_lpi_3_dfm_1_cse), (NOT reg_mult_37_res_lpi_3_dfm_1_cse),
      (NOT reg_mult_44_res_lpi_3_dfm_1_cse), STD_LOGIC_VECTOR'( (fsm_output(2)) &
      (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  acc_53_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_106_lpi_3_dfm_7 & '1')
      + UNSIGNED(butterFly1_3_mux1h_18_nl & '1'), 33));
  z_out_114 <= acc_53_nl(32 DOWNTO 1);
  butterFly1_4_mux1h_18_nl <= MUX1HOT_v_32_4_2((NOT reg_mult_4_res_lpi_3_dfm_1_cse),
      (NOT reg_mult_9_res_lpi_3_dfm_1_cse), (NOT reg_mult_38_res_lpi_3_dfm_1_cse),
      (NOT reg_mult_43_res_lpi_3_dfm_1_cse), STD_LOGIC_VECTOR'( (fsm_output(2)) &
      (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  acc_54_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_108_lpi_3_dfm_7 & '1')
      + UNSIGNED(butterFly1_4_mux1h_18_nl & '1'), 33));
  z_out_115 <= acc_54_nl(32 DOWNTO 1);
  butterFly1_5_mux1h_18_nl <= MUX1HOT_v_32_4_2((NOT reg_mult_5_res_lpi_3_dfm_1_cse),
      (NOT reg_mult_1_res_lpi_3_dfm_1_cse), (NOT reg_mult_39_res_lpi_3_dfm_1_cse),
      (NOT reg_mult_42_res_lpi_3_dfm_1_cse), STD_LOGIC_VECTOR'( (fsm_output(2)) &
      (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  acc_55_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_110_lpi_3_dfm_7 & '1')
      + UNSIGNED(butterFly1_5_mux1h_18_nl & '1'), 33));
  z_out_116 <= acc_55_nl(32 DOWNTO 1);
  butterFly1_6_mux1h_18_nl <= MUX1HOT_v_32_4_2((NOT reg_mult_6_res_lpi_3_dfm_1_cse),
      (NOT reg_mult_10_res_lpi_3_dfm_1_cse), (NOT reg_mult_40_res_lpi_3_dfm_1_cse),
      (NOT reg_mult_41_res_lpi_3_dfm_1_cse), STD_LOGIC_VECTOR'( (fsm_output(2)) &
      (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  acc_56_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_112_lpi_3_dfm_7 & '1')
      + UNSIGNED(butterFly1_6_mux1h_18_nl & '1'), 33));
  z_out_117 <= acc_56_nl(32 DOWNTO 1);
  butterFly1_7_mux1h_18_nl <= MUX1HOT_v_32_4_2((NOT reg_mult_7_res_lpi_3_dfm_1_cse),
      (NOT reg_mult_11_res_lpi_3_dfm_1_cse), (NOT reg_mult_41_res_lpi_3_dfm_1_cse),
      (NOT reg_mult_40_res_lpi_3_dfm_1_cse), STD_LOGIC_VECTOR'( (fsm_output(2)) &
      (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  acc_57_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_114_lpi_3_dfm_7 & '1')
      + UNSIGNED(butterFly1_7_mux1h_18_nl & '1'), 33));
  z_out_118 <= acc_57_nl(32 DOWNTO 1);
  butterFly1_8_mux1h_18_nl <= MUX1HOT_v_32_4_2((NOT reg_mult_8_res_lpi_3_dfm_1_cse),
      (NOT reg_mult_12_res_lpi_3_dfm_1_cse), (NOT reg_mult_42_res_lpi_3_dfm_1_cse),
      (NOT reg_mult_39_res_lpi_3_dfm_1_cse), STD_LOGIC_VECTOR'( (fsm_output(2)) &
      (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  acc_58_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_116_lpi_3_dfm_7 & '1')
      + UNSIGNED(butterFly1_8_mux1h_18_nl & '1'), 33));
  z_out_119 <= acc_58_nl(32 DOWNTO 1);
  butterFly1_9_mux1h_274_nl <= MUX1HOT_v_32_4_2((NOT reg_mult_9_res_lpi_3_dfm_1_cse),
      (NOT reg_mult_13_res_lpi_3_dfm_1_cse), (NOT reg_mult_43_res_lpi_3_dfm_1_cse),
      (NOT reg_mult_38_res_lpi_3_dfm_1_cse), STD_LOGIC_VECTOR'( (fsm_output(2)) &
      (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  acc_59_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_118_lpi_3_dfm_7 & '1')
      + UNSIGNED(butterFly1_9_mux1h_274_nl & '1'), 33));
  z_out_120 <= acc_59_nl(32 DOWNTO 1);
  butterFly1_10_mux1h_18_nl <= MUX1HOT_v_32_4_2((NOT reg_mult_10_res_lpi_3_dfm_1_cse),
      (NOT reg_mult_14_res_lpi_3_dfm_1_cse), (NOT reg_mult_44_res_lpi_3_dfm_1_cse),
      (NOT reg_mult_37_res_lpi_3_dfm_1_cse), STD_LOGIC_VECTOR'( (fsm_output(2)) &
      (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  acc_60_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_120_lpi_3_dfm_7 & '1')
      + UNSIGNED(butterFly1_10_mux1h_18_nl & '1'), 33));
  z_out_121 <= acc_60_nl(32 DOWNTO 1);
  butterFly1_11_mux1h_18_nl <= MUX1HOT_v_32_4_2((NOT reg_mult_11_res_lpi_3_dfm_1_cse),
      (NOT reg_mult_15_res_lpi_3_dfm_1_cse), (NOT reg_mult_45_res_lpi_3_dfm_1_cse),
      (NOT reg_mult_36_res_lpi_3_dfm_1_cse), STD_LOGIC_VECTOR'( (fsm_output(2)) &
      (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  acc_61_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_122_lpi_3_dfm_7 & '1')
      + UNSIGNED(butterFly1_11_mux1h_18_nl & '1'), 33));
  z_out_122 <= acc_61_nl(32 DOWNTO 1);
  butterFly1_12_mux1h_18_nl <= MUX1HOT_v_32_4_2((NOT reg_mult_12_res_lpi_3_dfm_1_cse),
      (NOT reg_mult_2_res_lpi_3_dfm_1_cse), (NOT reg_mult_46_res_lpi_3_dfm_1_cse),
      (NOT reg_mult_35_res_lpi_3_dfm_1_cse), STD_LOGIC_VECTOR'( (fsm_output(2)) &
      (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  acc_62_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_124_lpi_3_dfm_7 & '1')
      + UNSIGNED(butterFly1_12_mux1h_18_nl & '1'), 33));
  z_out_123 <= acc_62_nl(32 DOWNTO 1);
  butterFly1_13_mux1h_18_nl <= MUX1HOT_v_32_4_2((NOT reg_mult_13_res_lpi_3_dfm_1_cse),
      (NOT reg_mult_3_res_lpi_3_dfm_1_cse), (NOT reg_mult_47_res_lpi_3_dfm_1_cse),
      (NOT reg_mult_34_res_lpi_3_dfm_1_cse), STD_LOGIC_VECTOR'( (fsm_output(2)) &
      (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  acc_63_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_126_lpi_3_dfm_7 & '1')
      + UNSIGNED(butterFly1_13_mux1h_18_nl & '1'), 33));
  z_out_124 <= acc_63_nl(32 DOWNTO 1);
  butterFly1_14_mux1h_18_nl <= MUX1HOT_v_32_4_2((NOT reg_mult_14_res_lpi_3_dfm_1_cse),
      (NOT reg_mult_4_res_lpi_3_dfm_1_cse), (NOT reg_mult_32_res_lpi_3_dfm_1_cse),
      (NOT reg_mult_33_res_lpi_3_dfm_1_cse), STD_LOGIC_VECTOR'( (fsm_output(2)) &
      (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  acc_64_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_60_lpi_3_dfm_7 & '1')
      + UNSIGNED(butterFly1_14_mux1h_18_nl & '1'), 33));
  z_out_125 <= acc_64_nl(32 DOWNTO 1);
  butterFly1_15_mux1h_79_nl <= MUX1HOT_v_32_4_2((NOT reg_mult_15_res_lpi_3_dfm_1_cse),
      (NOT reg_mult_res_lpi_3_dfm_1_cse), (NOT reg_mult_33_res_lpi_3_dfm_1_cse),
      (NOT reg_mult_32_res_lpi_3_dfm_1_cse), STD_LOGIC_VECTOR'( (fsm_output(2)) &
      (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  acc_65_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_62_lpi_3_dfm_7 & '1')
      + UNSIGNED(butterFly1_15_mux1h_79_nl & '1'), 33));
  z_out_126 <= acc_65_nl(32 DOWNTO 1);
  butterFly1_15_mux1h_80_nl <= MUX1HOT_v_32_4_2(reg_mult_15_res_lpi_3_dfm_1_cse,
      reg_mult_res_lpi_3_dfm_1_cse, reg_mult_33_res_lpi_3_dfm_1_cse, reg_mult_32_res_lpi_3_dfm_1_cse,
      STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  z_out_127 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_62_lpi_3_dfm_7) + UNSIGNED(butterFly1_15_mux1h_80_nl),
      32));
  butterFly1_14_mux1h_19_nl <= MUX1HOT_v_32_4_2(reg_mult_14_res_lpi_3_dfm_1_cse,
      reg_mult_4_res_lpi_3_dfm_1_cse, reg_mult_32_res_lpi_3_dfm_1_cse, reg_mult_33_res_lpi_3_dfm_1_cse,
      STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  z_out_128 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_60_lpi_3_dfm_7) + UNSIGNED(butterFly1_14_mux1h_19_nl),
      32));
  butterFly1_13_mux1h_19_nl <= MUX1HOT_v_32_4_2(reg_mult_13_res_lpi_3_dfm_1_cse,
      reg_mult_3_res_lpi_3_dfm_1_cse, reg_mult_47_res_lpi_3_dfm_1_cse, reg_mult_34_res_lpi_3_dfm_1_cse,
      STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  z_out_129 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_126_lpi_3_dfm_7) + UNSIGNED(butterFly1_13_mux1h_19_nl),
      32));
  butterFly1_12_mux1h_19_nl <= MUX1HOT_v_32_4_2(reg_mult_12_res_lpi_3_dfm_1_cse,
      reg_mult_2_res_lpi_3_dfm_1_cse, reg_mult_46_res_lpi_3_dfm_1_cse, reg_mult_35_res_lpi_3_dfm_1_cse,
      STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  z_out_130 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_124_lpi_3_dfm_7) + UNSIGNED(butterFly1_12_mux1h_19_nl),
      32));
  butterFly1_11_mux1h_19_nl <= MUX1HOT_v_32_4_2(reg_mult_11_res_lpi_3_dfm_1_cse,
      reg_mult_15_res_lpi_3_dfm_1_cse, reg_mult_45_res_lpi_3_dfm_1_cse, reg_mult_36_res_lpi_3_dfm_1_cse,
      STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  z_out_131 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_122_lpi_3_dfm_7) + UNSIGNED(butterFly1_11_mux1h_19_nl),
      32));
  butterFly1_10_mux1h_19_nl <= MUX1HOT_v_32_4_2(reg_mult_10_res_lpi_3_dfm_1_cse,
      reg_mult_14_res_lpi_3_dfm_1_cse, reg_mult_44_res_lpi_3_dfm_1_cse, reg_mult_37_res_lpi_3_dfm_1_cse,
      STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  z_out_132 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_120_lpi_3_dfm_7) + UNSIGNED(butterFly1_10_mux1h_19_nl),
      32));
  butterFly1_9_mux1h_275_nl <= MUX1HOT_v_32_4_2(reg_mult_9_res_lpi_3_dfm_1_cse, reg_mult_13_res_lpi_3_dfm_1_cse,
      reg_mult_43_res_lpi_3_dfm_1_cse, reg_mult_38_res_lpi_3_dfm_1_cse, STD_LOGIC_VECTOR'(
      (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  z_out_133 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_118_lpi_3_dfm_7) + UNSIGNED(butterFly1_9_mux1h_275_nl),
      32));
  butterFly1_8_mux1h_19_nl <= MUX1HOT_v_32_4_2(reg_mult_8_res_lpi_3_dfm_1_cse, reg_mult_12_res_lpi_3_dfm_1_cse,
      reg_mult_42_res_lpi_3_dfm_1_cse, reg_mult_39_res_lpi_3_dfm_1_cse, STD_LOGIC_VECTOR'(
      (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  z_out_134 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_116_lpi_3_dfm_7) + UNSIGNED(butterFly1_8_mux1h_19_nl),
      32));
  butterFly1_7_mux1h_19_nl <= MUX1HOT_v_32_4_2(reg_mult_7_res_lpi_3_dfm_1_cse, reg_mult_11_res_lpi_3_dfm_1_cse,
      reg_mult_41_res_lpi_3_dfm_1_cse, reg_mult_40_res_lpi_3_dfm_1_cse, STD_LOGIC_VECTOR'(
      (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  z_out_135 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_114_lpi_3_dfm_7) + UNSIGNED(butterFly1_7_mux1h_19_nl),
      32));
  butterFly1_6_mux1h_19_nl <= MUX1HOT_v_32_4_2(reg_mult_6_res_lpi_3_dfm_1_cse, reg_mult_10_res_lpi_3_dfm_1_cse,
      reg_mult_40_res_lpi_3_dfm_1_cse, reg_mult_41_res_lpi_3_dfm_1_cse, STD_LOGIC_VECTOR'(
      (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  z_out_136 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_112_lpi_3_dfm_7) + UNSIGNED(butterFly1_6_mux1h_19_nl),
      32));
  butterFly1_5_mux1h_19_nl <= MUX1HOT_v_32_4_2(reg_mult_5_res_lpi_3_dfm_1_cse, reg_mult_1_res_lpi_3_dfm_1_cse,
      reg_mult_39_res_lpi_3_dfm_1_cse, reg_mult_42_res_lpi_3_dfm_1_cse, STD_LOGIC_VECTOR'(
      (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  z_out_137 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_110_lpi_3_dfm_7) + UNSIGNED(butterFly1_5_mux1h_19_nl),
      32));
  butterFly1_4_mux1h_19_nl <= MUX1HOT_v_32_4_2(reg_mult_4_res_lpi_3_dfm_1_cse, reg_mult_9_res_lpi_3_dfm_1_cse,
      reg_mult_38_res_lpi_3_dfm_1_cse, reg_mult_43_res_lpi_3_dfm_1_cse, STD_LOGIC_VECTOR'(
      (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  z_out_138 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_108_lpi_3_dfm_7) + UNSIGNED(butterFly1_4_mux1h_19_nl),
      32));
  butterFly1_3_mux1h_19_nl <= MUX1HOT_v_32_4_2(reg_mult_3_res_lpi_3_dfm_1_cse, reg_mult_8_res_lpi_3_dfm_1_cse,
      reg_mult_37_res_lpi_3_dfm_1_cse, reg_mult_44_res_lpi_3_dfm_1_cse, STD_LOGIC_VECTOR'(
      (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  z_out_139 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_106_lpi_3_dfm_7) + UNSIGNED(butterFly1_3_mux1h_19_nl),
      32));
  butterFly1_2_mux1h_19_nl <= MUX1HOT_v_32_4_2(reg_mult_2_res_lpi_3_dfm_1_cse, reg_mult_7_res_lpi_3_dfm_1_cse,
      reg_mult_36_res_lpi_3_dfm_1_cse, reg_mult_45_res_lpi_3_dfm_1_cse, STD_LOGIC_VECTOR'(
      (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  z_out_140 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_104_lpi_3_dfm_7) + UNSIGNED(butterFly1_2_mux1h_19_nl),
      32));
  butterFly1_1_mux1h_19_nl <= MUX1HOT_v_32_4_2(reg_mult_1_res_lpi_3_dfm_1_cse, reg_mult_6_res_lpi_3_dfm_1_cse,
      reg_mult_35_res_lpi_3_dfm_1_cse, reg_mult_46_res_lpi_3_dfm_1_cse, STD_LOGIC_VECTOR'(
      (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  z_out_141 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_102_lpi_3_dfm_7) + UNSIGNED(butterFly1_1_mux1h_19_nl),
      32));
  butterFly1_mux1h_19_nl <= MUX1HOT_v_32_4_2(reg_mult_res_lpi_3_dfm_1_cse, reg_mult_5_res_lpi_3_dfm_1_cse,
      reg_mult_34_res_lpi_3_dfm_1_cse, reg_mult_47_res_lpi_3_dfm_1_cse, STD_LOGIC_VECTOR'(
      (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  z_out_142 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_10_lpi_3_dfm_7) + UNSIGNED(butterFly1_mux1h_19_nl),
      32));
  modulo_add_1_mux1h_3_nl <= MUX1HOT_v_32_3_2((NOT z_out_141), (NOT z_out_138), (NOT
      z_out_127), STD_LOGIC_VECTOR'( modulo_add_1_qelse_or_m1c & (fsm_output(7))
      & (fsm_output(9))));
  acc_82_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & p_sva & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(modulo_add_1_mux1h_3_nl
      & '1'), 33), 34), 34));
  z_out_143_32 <= acc_82_nl(33);
  modulo_add_10_mux1h_3_nl <= MUX1HOT_v_32_4_2((NOT z_out_132), (NOT z_out_127),
      (NOT z_out_128), (NOT z_out_131), STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4))
      & (fsm_output(7)) & (fsm_output(9))));
  acc_83_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & p_sva & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(modulo_add_10_mux1h_3_nl
      & '1'), 33), 34), 34));
  z_out_144_32 <= acc_83_nl(33);
  modulo_add_54_mux1h_3_nl <= MUX1HOT_v_32_4_2((NOT z_out_136), (NOT z_out_133),
      (NOT z_out_135), (NOT z_out_134), STD_LOGIC_VECTOR'( (fsm_output(9)) & (fsm_output(7))
      & (fsm_output(2)) & (fsm_output(4))));
  acc_84_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & p_sva & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(modulo_add_54_mux1h_3_nl
      & '1'), 33), 34), 34));
  z_out_145_32 <= acc_84_nl(33);
  modulo_add_48_mux1h_3_nl <= MUX1HOT_v_32_4_2((NOT z_out_142), (NOT z_out_131),
      (NOT z_out_137), (NOT z_out_129), STD_LOGIC_VECTOR'( (fsm_output(9)) & (fsm_output(2))
      & (fsm_output(4)) & (fsm_output(7))));
  acc_85_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & p_sva & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(modulo_add_48_mux1h_3_nl
      & '1'), 33), 34), 34));
  z_out_146_32 <= acc_85_nl(33);
  modulo_add_33_mux1h_3_nl <= MUX1HOT_v_32_3_2((NOT z_out_127), (NOT z_out_141),
      (NOT z_out_130), STD_LOGIC_VECTOR'( (fsm_output(7)) & (fsm_output(9)) & modulo_add_1_qelse_or_m1c));
  acc_86_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & p_sva & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(modulo_add_33_mux1h_3_nl
      & '1'), 33), 34), 34));
  z_out_147_32 <= acc_86_nl(33);
  modulo_add_34_mux1h_3_nl <= MUX1HOT_v_32_3_2((NOT z_out_142), (NOT z_out_132),
      (NOT z_out_131), STD_LOGIC_VECTOR'( or_dcpl_353 & (fsm_output(9)) & (fsm_output(4))));
  acc_87_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & p_sva & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(modulo_add_34_mux1h_3_nl
      & '1'), 33), 34), 34));
  z_out_148_32 <= acc_87_nl(33);
  modulo_add_6_mux1h_3_nl <= MUX1HOT_v_32_4_2((NOT z_out_136), (NOT z_out_135), (NOT
      z_out_132), (NOT z_out_128), STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4))
      & (fsm_output(7)) & (fsm_output(9))));
  acc_88_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & p_sva & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(modulo_add_6_mux1h_3_nl
      & '1'), 33), 34), 34));
  z_out_149_32 <= acc_88_nl(33);
  modulo_add_50_mux1h_3_nl <= MUX1HOT_v_32_3_2((NOT z_out_140), (NOT z_out_129),
      (NOT z_out_141), STD_LOGIC_VECTOR'( (fsm_output(9)) & modulo_add_1_qelse_or_m1c
      & (fsm_output(7))));
  acc_89_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & p_sva & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(modulo_add_50_mux1h_3_nl
      & '1'), 33), 34), 34));
  z_out_150_32 <= acc_89_nl(33);
  modulo_add_51_mux1h_3_nl <= MUX1HOT_v_32_4_2((NOT z_out_139), (NOT z_out_137),
      (NOT z_out_136), (NOT z_out_134), STD_LOGIC_VECTOR'( (fsm_output(9)) & (fsm_output(2))
      & (fsm_output(4)) & (fsm_output(7))));
  acc_90_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & p_sva & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(modulo_add_51_mux1h_3_nl
      & '1'), 33), 34), 34));
  z_out_151_32 <= acc_90_nl(33);
  modulo_add_14_mux1h_3_nl <= MUX1HOT_v_32_3_2((NOT z_out_128), (NOT z_out_133),
      (NOT z_out_130), STD_LOGIC_VECTOR'( modulo_add_1_qelse_or_m1c & (fsm_output(9))
      & (fsm_output(7))));
  acc_91_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & p_sva & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(modulo_add_14_mux1h_3_nl
      & '1'), 33), 34), 34));
  z_out_152_32 <= acc_91_nl(33);
  modulo_add_36_mux1h_3_nl <= MUX1HOT_v_32_4_2((NOT z_out_140), (NOT z_out_127),
      (NOT z_out_142), (NOT z_out_130), STD_LOGIC_VECTOR'( (fsm_output(7)) & (fsm_output(2))
      & (fsm_output(4)) & (fsm_output(9))));
  acc_92_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & p_sva & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(modulo_add_36_mux1h_3_nl
      & '1'), 33), 34), 34));
  z_out_153_32 <= acc_92_nl(33);
  modulo_add_52_mux1h_3_nl <= MUX1HOT_v_32_4_2((NOT z_out_138), (NOT z_out_139),
      (NOT z_out_133), (NOT z_out_132), STD_LOGIC_VECTOR'( (fsm_output(9)) & (fsm_output(7))
      & (fsm_output(2)) & (fsm_output(4))));
  acc_93_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & p_sva & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(modulo_add_52_mux1h_3_nl
      & '1'), 33), 34), 34));
  z_out_154_32 <= acc_93_nl(33);
  modulo_add_41_mux1h_3_nl <= MUX1HOT_v_32_4_2((NOT z_out_135), (NOT z_out_134),
      (NOT z_out_133), (NOT z_out_129), STD_LOGIC_VECTOR'( (fsm_output(7)) & (fsm_output(2))
      & (fsm_output(4)) & (fsm_output(9))));
  acc_94_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & p_sva & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(modulo_add_41_mux1h_3_nl
      & '1'), 33), 34), 34));
  z_out_155_32 <= acc_94_nl(33);
  modulo_add_2_mux1h_3_nl <= MUX1HOT_v_32_3_2((NOT z_out_140), (NOT z_out_137), (NOT
      z_out_134), STD_LOGIC_VECTOR'( modulo_add_1_qelse_or_m1c & (fsm_output(7))
      & (fsm_output(9))));
  acc_95_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & p_sva & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(modulo_add_2_mux1h_3_nl
      & '1'), 33), 34), 34));
  z_out_156_32 <= acc_95_nl(33);
  modulo_add_53_mux1h_3_nl <= MUX1HOT_v_32_3_2((NOT z_out_137), (NOT z_out_136),
      (NOT z_out_138), STD_LOGIC_VECTOR'( (fsm_output(9)) & (fsm_output(7)) & modulo_add_1_qelse_or_m1c));
  acc_96_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & p_sva & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(modulo_add_53_mux1h_3_nl
      & '1'), 33), 34), 34));
  z_out_157_32 <= acc_96_nl(33);
  modulo_add_55_mux1h_3_nl <= MUX1HOT_v_32_3_2((NOT z_out_135), (NOT z_out_139),
      (NOT z_out_131), STD_LOGIC_VECTOR'( (fsm_output(9)) & modulo_add_1_qelse_or_m1c
      & (fsm_output(7))));
  acc_97_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & p_sva & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(modulo_add_55_mux1h_3_nl
      & '1'), 33), 34), 34));
  z_out_158_32 <= acc_97_nl(33);
  z_out <= MUX1HOT_v_32_8_2(xt_rsc_0_30_i_qa_d, xt_rsc_1_30_i_qa_d, xt_rsc_2_30_i_qa_d,
      xt_rsc_3_30_i_qa_d, xt_rsc_4_30_i_qa_d, xt_rsc_5_30_i_qa_d, xt_rsc_6_30_i_qa_d,
      xt_rsc_7_30_i_qa_d, STD_LOGIC_VECTOR'( butterFly1_15_f1_mux_cse & butterFly1_15_f1_mux_1_cse
      & butterFly1_15_f1_mux_2_cse & butterFly1_15_f1_mux_3_cse & butterFly1_15_f1_mux_4_cse
      & butterFly1_15_f1_mux_5_cse & butterFly1_15_f1_mux_6_cse & butterFly1_15_f1_mux_7_cse));
  z_out_1 <= MUX1HOT_v_32_8_2(xt_rsc_0_28_i_qa_d, xt_rsc_1_28_i_qa_d, xt_rsc_2_28_i_qa_d,
      xt_rsc_3_28_i_qa_d, xt_rsc_4_28_i_qa_d, xt_rsc_5_28_i_qa_d, xt_rsc_6_28_i_qa_d,
      xt_rsc_7_28_i_qa_d, STD_LOGIC_VECTOR'( butterFly1_15_f1_mux_cse & butterFly1_15_f1_mux_1_cse
      & butterFly1_15_f1_mux_2_cse & butterFly1_15_f1_mux_3_cse & butterFly1_15_f1_mux_4_cse
      & butterFly1_15_f1_mux_5_cse & butterFly1_15_f1_mux_6_cse & butterFly1_15_f1_mux_7_cse));
  z_out_2 <= MUX1HOT_v_32_8_2(xt_rsc_0_26_i_qa_d, xt_rsc_1_26_i_qa_d, xt_rsc_2_26_i_qa_d,
      xt_rsc_3_26_i_qa_d, xt_rsc_4_26_i_qa_d, xt_rsc_5_26_i_qa_d, xt_rsc_6_26_i_qa_d,
      xt_rsc_7_26_i_qa_d, STD_LOGIC_VECTOR'( butterFly1_15_f1_mux_cse & butterFly1_15_f1_mux_1_cse
      & butterFly1_15_f1_mux_2_cse & butterFly1_15_f1_mux_3_cse & butterFly1_15_f1_mux_4_cse
      & butterFly1_15_f1_mux_5_cse & butterFly1_15_f1_mux_6_cse & butterFly1_15_f1_mux_7_cse));
  z_out_3 <= MUX1HOT_v_32_8_2(xt_rsc_0_24_i_qa_d, xt_rsc_1_24_i_qa_d, xt_rsc_2_24_i_qa_d,
      xt_rsc_3_24_i_qa_d, xt_rsc_4_24_i_qa_d, xt_rsc_5_24_i_qa_d, xt_rsc_6_24_i_qa_d,
      xt_rsc_7_24_i_qa_d, STD_LOGIC_VECTOR'( butterFly1_15_f1_mux_cse & butterFly1_15_f1_mux_1_cse
      & butterFly1_15_f1_mux_2_cse & butterFly1_15_f1_mux_3_cse & butterFly1_15_f1_mux_4_cse
      & butterFly1_15_f1_mux_5_cse & butterFly1_15_f1_mux_6_cse & butterFly1_15_f1_mux_7_cse));
  z_out_4 <= MUX1HOT_v_32_8_2(xt_rsc_0_22_i_qa_d, xt_rsc_1_22_i_qa_d, xt_rsc_2_22_i_qa_d,
      xt_rsc_3_22_i_qa_d, xt_rsc_4_22_i_qa_d, xt_rsc_5_22_i_qa_d, xt_rsc_6_22_i_qa_d,
      xt_rsc_7_22_i_qa_d, STD_LOGIC_VECTOR'( butterFly1_15_f1_mux_cse & butterFly1_15_f1_mux_1_cse
      & butterFly1_15_f1_mux_2_cse & butterFly1_15_f1_mux_3_cse & butterFly1_15_f1_mux_4_cse
      & butterFly1_15_f1_mux_5_cse & butterFly1_15_f1_mux_6_cse & butterFly1_15_f1_mux_7_cse));
  z_out_5 <= MUX1HOT_v_32_8_2(xt_rsc_0_20_i_qa_d, xt_rsc_1_20_i_qa_d, xt_rsc_2_20_i_qa_d,
      xt_rsc_3_20_i_qa_d, xt_rsc_4_20_i_qa_d, xt_rsc_5_20_i_qa_d, xt_rsc_6_20_i_qa_d,
      xt_rsc_7_20_i_qa_d, STD_LOGIC_VECTOR'( butterFly1_15_f1_mux_cse & butterFly1_15_f1_mux_1_cse
      & butterFly1_15_f1_mux_2_cse & butterFly1_15_f1_mux_3_cse & butterFly1_15_f1_mux_4_cse
      & butterFly1_15_f1_mux_5_cse & butterFly1_15_f1_mux_6_cse & butterFly1_15_f1_mux_7_cse));
  z_out_6 <= MUX1HOT_v_32_8_2(xt_rsc_0_18_i_qa_d, xt_rsc_1_18_i_qa_d, xt_rsc_2_18_i_qa_d,
      xt_rsc_3_18_i_qa_d, xt_rsc_4_18_i_qa_d, xt_rsc_5_18_i_qa_d, xt_rsc_6_18_i_qa_d,
      xt_rsc_7_18_i_qa_d, STD_LOGIC_VECTOR'( butterFly1_15_f1_mux_cse & butterFly1_15_f1_mux_1_cse
      & butterFly1_15_f1_mux_2_cse & butterFly1_15_f1_mux_3_cse & butterFly1_15_f1_mux_4_cse
      & butterFly1_15_f1_mux_5_cse & butterFly1_15_f1_mux_6_cse & butterFly1_15_f1_mux_7_cse));
  z_out_7 <= MUX1HOT_v_32_8_2(xt_rsc_0_16_i_qa_d, xt_rsc_1_16_i_qa_d, xt_rsc_2_16_i_qa_d,
      xt_rsc_3_16_i_qa_d, xt_rsc_4_16_i_qa_d, xt_rsc_5_16_i_qa_d, xt_rsc_6_16_i_qa_d,
      xt_rsc_7_16_i_qa_d, STD_LOGIC_VECTOR'( butterFly1_15_f1_mux_cse & butterFly1_15_f1_mux_1_cse
      & butterFly1_15_f1_mux_2_cse & butterFly1_15_f1_mux_3_cse & butterFly1_15_f1_mux_4_cse
      & butterFly1_15_f1_mux_5_cse & butterFly1_15_f1_mux_6_cse & butterFly1_15_f1_mux_7_cse));
  z_out_8 <= MUX1HOT_v_32_8_2(xt_rsc_0_14_i_qa_d, xt_rsc_1_14_i_qa_d, xt_rsc_2_14_i_qa_d,
      xt_rsc_3_14_i_qa_d, xt_rsc_4_14_i_qa_d, xt_rsc_5_14_i_qa_d, xt_rsc_6_14_i_qa_d,
      xt_rsc_7_14_i_qa_d, STD_LOGIC_VECTOR'( butterFly1_15_f1_mux_cse & butterFly1_15_f1_mux_1_cse
      & butterFly1_15_f1_mux_2_cse & butterFly1_15_f1_mux_3_cse & butterFly1_15_f1_mux_4_cse
      & butterFly1_15_f1_mux_5_cse & butterFly1_15_f1_mux_6_cse & butterFly1_15_f1_mux_7_cse));
  z_out_9 <= MUX1HOT_v_32_8_2(xt_rsc_0_12_i_qa_d, xt_rsc_1_12_i_qa_d, xt_rsc_2_12_i_qa_d,
      xt_rsc_3_12_i_qa_d, xt_rsc_4_12_i_qa_d, xt_rsc_5_12_i_qa_d, xt_rsc_6_12_i_qa_d,
      xt_rsc_7_12_i_qa_d, STD_LOGIC_VECTOR'( butterFly1_15_f1_mux_cse & butterFly1_15_f1_mux_1_cse
      & butterFly1_15_f1_mux_2_cse & butterFly1_15_f1_mux_3_cse & butterFly1_15_f1_mux_4_cse
      & butterFly1_15_f1_mux_5_cse & butterFly1_15_f1_mux_6_cse & butterFly1_15_f1_mux_7_cse));
  z_out_10 <= MUX1HOT_v_32_8_2(xt_rsc_0_10_i_qa_d, xt_rsc_1_10_i_qa_d, xt_rsc_2_10_i_qa_d,
      xt_rsc_3_10_i_qa_d, xt_rsc_4_10_i_qa_d, xt_rsc_5_10_i_qa_d, xt_rsc_6_10_i_qa_d,
      xt_rsc_7_10_i_qa_d, STD_LOGIC_VECTOR'( butterFly1_15_f1_mux_cse & butterFly1_15_f1_mux_1_cse
      & butterFly1_15_f1_mux_2_cse & butterFly1_15_f1_mux_3_cse & butterFly1_15_f1_mux_4_cse
      & butterFly1_15_f1_mux_5_cse & butterFly1_15_f1_mux_6_cse & butterFly1_15_f1_mux_7_cse));
  z_out_11 <= MUX1HOT_v_32_8_2(xt_rsc_0_8_i_qa_d, xt_rsc_1_8_i_qa_d, xt_rsc_2_8_i_qa_d,
      xt_rsc_3_8_i_qa_d, xt_rsc_4_8_i_qa_d, xt_rsc_5_8_i_qa_d, xt_rsc_6_8_i_qa_d,
      xt_rsc_7_8_i_qa_d, STD_LOGIC_VECTOR'( butterFly1_15_f1_mux_cse & butterFly1_15_f1_mux_1_cse
      & butterFly1_15_f1_mux_2_cse & butterFly1_15_f1_mux_3_cse & butterFly1_15_f1_mux_4_cse
      & butterFly1_15_f1_mux_5_cse & butterFly1_15_f1_mux_6_cse & butterFly1_15_f1_mux_7_cse));
  z_out_12 <= MUX1HOT_v_32_8_2(xt_rsc_0_6_i_qa_d, xt_rsc_1_6_i_qa_d, xt_rsc_2_6_i_qa_d,
      xt_rsc_3_6_i_qa_d, xt_rsc_4_6_i_qa_d, xt_rsc_5_6_i_qa_d, xt_rsc_6_6_i_qa_d,
      xt_rsc_7_6_i_qa_d, STD_LOGIC_VECTOR'( butterFly1_15_f1_mux_cse & butterFly1_15_f1_mux_1_cse
      & butterFly1_15_f1_mux_2_cse & butterFly1_15_f1_mux_3_cse & butterFly1_15_f1_mux_4_cse
      & butterFly1_15_f1_mux_5_cse & butterFly1_15_f1_mux_6_cse & butterFly1_15_f1_mux_7_cse));
  z_out_13 <= MUX1HOT_v_32_8_2(xt_rsc_0_4_i_qa_d, xt_rsc_1_4_i_qa_d, xt_rsc_2_4_i_qa_d,
      xt_rsc_3_4_i_qa_d, xt_rsc_4_4_i_qa_d, xt_rsc_5_4_i_qa_d, xt_rsc_6_4_i_qa_d,
      xt_rsc_7_4_i_qa_d, STD_LOGIC_VECTOR'( butterFly1_15_f1_mux_cse & butterFly1_15_f1_mux_1_cse
      & butterFly1_15_f1_mux_2_cse & butterFly1_15_f1_mux_3_cse & butterFly1_15_f1_mux_4_cse
      & butterFly1_15_f1_mux_5_cse & butterFly1_15_f1_mux_6_cse & butterFly1_15_f1_mux_7_cse));
  z_out_14 <= MUX1HOT_v_32_8_2(xt_rsc_0_2_i_qa_d, xt_rsc_1_2_i_qa_d, xt_rsc_2_2_i_qa_d,
      xt_rsc_3_2_i_qa_d, xt_rsc_4_2_i_qa_d, xt_rsc_5_2_i_qa_d, xt_rsc_6_2_i_qa_d,
      xt_rsc_7_2_i_qa_d, STD_LOGIC_VECTOR'( butterFly1_15_f1_mux_cse & butterFly1_15_f1_mux_1_cse
      & butterFly1_15_f1_mux_2_cse & butterFly1_15_f1_mux_3_cse & butterFly1_15_f1_mux_4_cse
      & butterFly1_15_f1_mux_5_cse & butterFly1_15_f1_mux_6_cse & butterFly1_15_f1_mux_7_cse));
  z_out_15 <= MUX1HOT_v_32_8_2(xt_rsc_0_0_i_qa_d, xt_rsc_1_0_i_qa_d, xt_rsc_2_0_i_qa_d,
      xt_rsc_3_0_i_qa_d, xt_rsc_4_0_i_qa_d, xt_rsc_5_0_i_qa_d, xt_rsc_6_0_i_qa_d,
      xt_rsc_7_0_i_qa_d, STD_LOGIC_VECTOR'( butterFly1_15_f1_mux_cse & butterFly1_15_f1_mux_1_cse
      & butterFly1_15_f1_mux_2_cse & butterFly1_15_f1_mux_3_cse & butterFly1_15_f1_mux_4_cse
      & butterFly1_15_f1_mux_5_cse & butterFly1_15_f1_mux_6_cse & butterFly1_15_f1_mux_7_cse));
  z_out_16 <= MUX1HOT_v_32_8_2(yt_rsc_0_30_i_q_d, yt_rsc_1_30_i_q_d, yt_rsc_2_30_i_q_d,
      yt_rsc_3_30_i_q_d, yt_rsc_4_30_i_q_d, yt_rsc_5_30_i_q_d, yt_rsc_6_30_i_q_d,
      yt_rsc_7_30_i_q_d, STD_LOGIC_VECTOR'( butterFly1_31_f1_mux_cse & butterFly1_31_f1_mux_1_cse
      & butterFly1_31_f1_mux_2_cse & butterFly1_31_f1_mux_3_cse & butterFly1_31_f1_mux_4_cse
      & butterFly1_31_f1_mux_5_cse & butterFly1_31_f1_mux_6_cse & butterFly1_31_f1_mux_7_cse));
  z_out_17 <= MUX1HOT_v_32_8_2(yt_rsc_0_28_i_q_d, yt_rsc_1_28_i_q_d, yt_rsc_2_28_i_q_d,
      yt_rsc_3_28_i_q_d, yt_rsc_4_28_i_q_d, yt_rsc_5_28_i_q_d, yt_rsc_6_28_i_q_d,
      yt_rsc_7_28_i_q_d, STD_LOGIC_VECTOR'( butterFly1_31_f1_mux_cse & butterFly1_31_f1_mux_1_cse
      & butterFly1_31_f1_mux_2_cse & butterFly1_31_f1_mux_3_cse & butterFly1_31_f1_mux_4_cse
      & butterFly1_31_f1_mux_5_cse & butterFly1_31_f1_mux_6_cse & butterFly1_31_f1_mux_7_cse));
  z_out_18 <= MUX1HOT_v_32_8_2(yt_rsc_0_26_i_q_d, yt_rsc_1_26_i_q_d, yt_rsc_2_26_i_q_d,
      yt_rsc_3_26_i_q_d, yt_rsc_4_26_i_q_d, yt_rsc_5_26_i_q_d, yt_rsc_6_26_i_q_d,
      yt_rsc_7_26_i_q_d, STD_LOGIC_VECTOR'( butterFly1_31_f1_mux_cse & butterFly1_31_f1_mux_1_cse
      & butterFly1_31_f1_mux_2_cse & butterFly1_31_f1_mux_3_cse & butterFly1_31_f1_mux_4_cse
      & butterFly1_31_f1_mux_5_cse & butterFly1_31_f1_mux_6_cse & butterFly1_31_f1_mux_7_cse));
  z_out_19 <= MUX1HOT_v_32_8_2(yt_rsc_0_24_i_q_d, yt_rsc_1_24_i_q_d, yt_rsc_2_24_i_q_d,
      yt_rsc_3_24_i_q_d, yt_rsc_4_24_i_q_d, yt_rsc_5_24_i_q_d, yt_rsc_6_24_i_q_d,
      yt_rsc_7_24_i_q_d, STD_LOGIC_VECTOR'( butterFly1_31_f1_mux_cse & butterFly1_31_f1_mux_1_cse
      & butterFly1_31_f1_mux_2_cse & butterFly1_31_f1_mux_3_cse & butterFly1_31_f1_mux_4_cse
      & butterFly1_31_f1_mux_5_cse & butterFly1_31_f1_mux_6_cse & butterFly1_31_f1_mux_7_cse));
  z_out_20 <= MUX1HOT_v_32_8_2(yt_rsc_0_22_i_q_d, yt_rsc_1_22_i_q_d, yt_rsc_2_22_i_q_d,
      yt_rsc_3_22_i_q_d, yt_rsc_4_22_i_q_d, yt_rsc_5_22_i_q_d, yt_rsc_6_22_i_q_d,
      yt_rsc_7_22_i_q_d, STD_LOGIC_VECTOR'( butterFly1_31_f1_mux_cse & butterFly1_31_f1_mux_1_cse
      & butterFly1_31_f1_mux_2_cse & butterFly1_31_f1_mux_3_cse & butterFly1_31_f1_mux_4_cse
      & butterFly1_31_f1_mux_5_cse & butterFly1_31_f1_mux_6_cse & butterFly1_31_f1_mux_7_cse));
  z_out_21 <= MUX1HOT_v_32_8_2(yt_rsc_0_20_i_q_d, yt_rsc_1_20_i_q_d, yt_rsc_2_20_i_q_d,
      yt_rsc_3_20_i_q_d, yt_rsc_4_20_i_q_d, yt_rsc_5_20_i_q_d, yt_rsc_6_20_i_q_d,
      yt_rsc_7_20_i_q_d, STD_LOGIC_VECTOR'( butterFly1_31_f1_mux_cse & butterFly1_31_f1_mux_1_cse
      & butterFly1_31_f1_mux_2_cse & butterFly1_31_f1_mux_3_cse & butterFly1_31_f1_mux_4_cse
      & butterFly1_31_f1_mux_5_cse & butterFly1_31_f1_mux_6_cse & butterFly1_31_f1_mux_7_cse));
  z_out_22 <= MUX1HOT_v_32_8_2(yt_rsc_0_18_i_q_d, yt_rsc_1_18_i_q_d, yt_rsc_2_18_i_q_d,
      yt_rsc_3_18_i_q_d, yt_rsc_4_18_i_q_d, yt_rsc_5_18_i_q_d, yt_rsc_6_18_i_q_d,
      yt_rsc_7_18_i_q_d, STD_LOGIC_VECTOR'( butterFly1_31_f1_mux_cse & butterFly1_31_f1_mux_1_cse
      & butterFly1_31_f1_mux_2_cse & butterFly1_31_f1_mux_3_cse & butterFly1_31_f1_mux_4_cse
      & butterFly1_31_f1_mux_5_cse & butterFly1_31_f1_mux_6_cse & butterFly1_31_f1_mux_7_cse));
  z_out_23 <= MUX1HOT_v_32_8_2(yt_rsc_0_16_i_q_d, yt_rsc_1_16_i_q_d, yt_rsc_2_16_i_q_d,
      yt_rsc_3_16_i_q_d, yt_rsc_4_16_i_q_d, yt_rsc_5_16_i_q_d, yt_rsc_6_16_i_q_d,
      yt_rsc_7_16_i_q_d, STD_LOGIC_VECTOR'( butterFly1_31_f1_mux_cse & butterFly1_31_f1_mux_1_cse
      & butterFly1_31_f1_mux_2_cse & butterFly1_31_f1_mux_3_cse & butterFly1_31_f1_mux_4_cse
      & butterFly1_31_f1_mux_5_cse & butterFly1_31_f1_mux_6_cse & butterFly1_31_f1_mux_7_cse));
  z_out_24 <= MUX1HOT_v_32_8_2(yt_rsc_0_14_i_q_d, yt_rsc_1_14_i_q_d, yt_rsc_2_14_i_q_d,
      yt_rsc_3_14_i_q_d, yt_rsc_4_14_i_q_d, yt_rsc_5_14_i_q_d, yt_rsc_6_14_i_q_d,
      yt_rsc_7_14_i_q_d, STD_LOGIC_VECTOR'( butterFly1_31_f1_mux_cse & butterFly1_31_f1_mux_1_cse
      & butterFly1_31_f1_mux_2_cse & butterFly1_31_f1_mux_3_cse & butterFly1_31_f1_mux_4_cse
      & butterFly1_31_f1_mux_5_cse & butterFly1_31_f1_mux_6_cse & butterFly1_31_f1_mux_7_cse));
  z_out_25 <= MUX1HOT_v_32_8_2(yt_rsc_0_12_i_q_d, yt_rsc_1_12_i_q_d, yt_rsc_2_12_i_q_d,
      yt_rsc_3_12_i_q_d, yt_rsc_4_12_i_q_d, yt_rsc_5_12_i_q_d, yt_rsc_6_12_i_q_d,
      yt_rsc_7_12_i_q_d, STD_LOGIC_VECTOR'( butterFly1_31_f1_mux_cse & butterFly1_31_f1_mux_1_cse
      & butterFly1_31_f1_mux_2_cse & butterFly1_31_f1_mux_3_cse & butterFly1_31_f1_mux_4_cse
      & butterFly1_31_f1_mux_5_cse & butterFly1_31_f1_mux_6_cse & butterFly1_31_f1_mux_7_cse));
  z_out_26 <= MUX1HOT_v_32_8_2(yt_rsc_0_10_i_q_d, yt_rsc_1_10_i_q_d, yt_rsc_2_10_i_q_d,
      yt_rsc_3_10_i_q_d, yt_rsc_4_10_i_q_d, yt_rsc_5_10_i_q_d, yt_rsc_6_10_i_q_d,
      yt_rsc_7_10_i_q_d, STD_LOGIC_VECTOR'( butterFly1_31_f1_mux_cse & butterFly1_31_f1_mux_1_cse
      & butterFly1_31_f1_mux_2_cse & butterFly1_31_f1_mux_3_cse & butterFly1_31_f1_mux_4_cse
      & butterFly1_31_f1_mux_5_cse & butterFly1_31_f1_mux_6_cse & butterFly1_31_f1_mux_7_cse));
  z_out_27 <= MUX1HOT_v_32_8_2(yt_rsc_0_8_i_q_d, yt_rsc_1_8_i_q_d, yt_rsc_2_8_i_q_d,
      yt_rsc_3_8_i_q_d, yt_rsc_4_8_i_q_d, yt_rsc_5_8_i_q_d, yt_rsc_6_8_i_q_d, yt_rsc_7_8_i_q_d,
      STD_LOGIC_VECTOR'( butterFly1_31_f1_mux_cse & butterFly1_31_f1_mux_1_cse &
      butterFly1_31_f1_mux_2_cse & butterFly1_31_f1_mux_3_cse & butterFly1_31_f1_mux_4_cse
      & butterFly1_31_f1_mux_5_cse & butterFly1_31_f1_mux_6_cse & butterFly1_31_f1_mux_7_cse));
  z_out_28 <= MUX1HOT_v_32_8_2(yt_rsc_0_6_i_q_d, yt_rsc_1_6_i_q_d, yt_rsc_2_6_i_q_d,
      yt_rsc_3_6_i_q_d, yt_rsc_4_6_i_q_d, yt_rsc_5_6_i_q_d, yt_rsc_6_6_i_q_d, yt_rsc_7_6_i_q_d,
      STD_LOGIC_VECTOR'( butterFly1_31_f1_mux_cse & butterFly1_31_f1_mux_1_cse &
      butterFly1_31_f1_mux_2_cse & butterFly1_31_f1_mux_3_cse & butterFly1_31_f1_mux_4_cse
      & butterFly1_31_f1_mux_5_cse & butterFly1_31_f1_mux_6_cse & butterFly1_31_f1_mux_7_cse));
  z_out_29 <= MUX1HOT_v_32_8_2(yt_rsc_0_4_i_q_d, yt_rsc_1_4_i_q_d, yt_rsc_2_4_i_q_d,
      yt_rsc_3_4_i_q_d, yt_rsc_4_4_i_q_d, yt_rsc_5_4_i_q_d, yt_rsc_6_4_i_q_d, yt_rsc_7_4_i_q_d,
      STD_LOGIC_VECTOR'( butterFly1_31_f1_mux_cse & butterFly1_31_f1_mux_1_cse &
      butterFly1_31_f1_mux_2_cse & butterFly1_31_f1_mux_3_cse & butterFly1_31_f1_mux_4_cse
      & butterFly1_31_f1_mux_5_cse & butterFly1_31_f1_mux_6_cse & butterFly1_31_f1_mux_7_cse));
  z_out_30 <= MUX1HOT_v_32_8_2(yt_rsc_0_2_i_q_d, yt_rsc_1_2_i_q_d, yt_rsc_2_2_i_q_d,
      yt_rsc_3_2_i_q_d, yt_rsc_4_2_i_q_d, yt_rsc_5_2_i_q_d, yt_rsc_6_2_i_q_d, yt_rsc_7_2_i_q_d,
      STD_LOGIC_VECTOR'( butterFly1_31_f1_mux_cse & butterFly1_31_f1_mux_1_cse &
      butterFly1_31_f1_mux_2_cse & butterFly1_31_f1_mux_3_cse & butterFly1_31_f1_mux_4_cse
      & butterFly1_31_f1_mux_5_cse & butterFly1_31_f1_mux_6_cse & butterFly1_31_f1_mux_7_cse));
  z_out_31 <= MUX1HOT_v_32_8_2(yt_rsc_0_0_i_q_d, yt_rsc_1_0_i_q_d, yt_rsc_2_0_i_q_d,
      yt_rsc_3_0_i_q_d, yt_rsc_4_0_i_q_d, yt_rsc_5_0_i_q_d, yt_rsc_6_0_i_q_d, yt_rsc_7_0_i_q_d,
      STD_LOGIC_VECTOR'( butterFly1_31_f1_mux_cse & butterFly1_31_f1_mux_1_cse &
      butterFly1_31_f1_mux_2_cse & butterFly1_31_f1_mux_3_cse & butterFly1_31_f1_mux_4_cse
      & butterFly1_31_f1_mux_5_cse & butterFly1_31_f1_mux_6_cse & butterFly1_31_f1_mux_7_cse));
  z_out_32 <= MUX1HOT_v_32_8_2(yt_rsc_0_3_i_q_d, yt_rsc_1_3_i_q_d, yt_rsc_2_3_i_q_d,
      yt_rsc_3_3_i_q_d, yt_rsc_4_3_i_q_d, yt_rsc_5_3_i_q_d, yt_rsc_6_3_i_q_d, yt_rsc_7_3_i_q_d,
      STD_LOGIC_VECTOR'( butterFly1_31_f1_mux_cse & butterFly1_31_f1_mux_1_cse &
      butterFly1_31_f1_mux_2_cse & butterFly1_31_f1_mux_3_cse & butterFly1_31_f1_mux_4_cse
      & butterFly1_31_f1_mux_5_cse & butterFly1_31_f1_mux_6_cse & butterFly1_31_f1_mux_7_cse));
  z_out_33 <= MUX1HOT_v_32_8_2(yt_rsc_0_5_i_q_d, yt_rsc_1_5_i_q_d, yt_rsc_2_5_i_q_d,
      yt_rsc_3_5_i_q_d, yt_rsc_4_5_i_q_d, yt_rsc_5_5_i_q_d, yt_rsc_6_5_i_q_d, yt_rsc_7_5_i_q_d,
      STD_LOGIC_VECTOR'( butterFly1_31_f1_mux_cse & butterFly1_31_f1_mux_1_cse &
      butterFly1_31_f1_mux_2_cse & butterFly1_31_f1_mux_3_cse & butterFly1_31_f1_mux_4_cse
      & butterFly1_31_f1_mux_5_cse & butterFly1_31_f1_mux_6_cse & butterFly1_31_f1_mux_7_cse));
  z_out_34 <= MUX1HOT_v_32_8_2(yt_rsc_0_7_i_q_d, yt_rsc_1_7_i_q_d, yt_rsc_2_7_i_q_d,
      yt_rsc_3_7_i_q_d, yt_rsc_4_7_i_q_d, yt_rsc_5_7_i_q_d, yt_rsc_6_7_i_q_d, yt_rsc_7_7_i_q_d,
      STD_LOGIC_VECTOR'( butterFly1_31_f1_mux_cse & butterFly1_31_f1_mux_1_cse &
      butterFly1_31_f1_mux_2_cse & butterFly1_31_f1_mux_3_cse & butterFly1_31_f1_mux_4_cse
      & butterFly1_31_f1_mux_5_cse & butterFly1_31_f1_mux_6_cse & butterFly1_31_f1_mux_7_cse));
  z_out_35 <= MUX1HOT_v_32_8_2(yt_rsc_0_31_i_q_d, yt_rsc_1_31_i_q_d, yt_rsc_2_31_i_q_d,
      yt_rsc_3_31_i_q_d, yt_rsc_4_31_i_q_d, yt_rsc_5_31_i_q_d, yt_rsc_6_31_i_q_d,
      yt_rsc_7_31_i_q_d, STD_LOGIC_VECTOR'( butterFly1_31_f1_mux_cse & butterFly1_31_f1_mux_1_cse
      & butterFly1_31_f1_mux_2_cse & butterFly1_31_f1_mux_3_cse & butterFly1_31_f1_mux_4_cse
      & butterFly1_31_f1_mux_5_cse & butterFly1_31_f1_mux_6_cse & butterFly1_31_f1_mux_7_cse));
  z_out_36 <= MUX1HOT_v_32_8_2(xt_rsc_0_11_i_qa_d, xt_rsc_1_11_i_qa_d, xt_rsc_2_11_i_qa_d,
      xt_rsc_3_11_i_qa_d, xt_rsc_4_11_i_qa_d, xt_rsc_5_11_i_qa_d, xt_rsc_6_11_i_qa_d,
      xt_rsc_7_11_i_qa_d, STD_LOGIC_VECTOR'( butterFly1_15_f1_mux_cse & butterFly1_15_f1_mux_1_cse
      & butterFly1_15_f1_mux_2_cse & butterFly1_15_f1_mux_3_cse & butterFly1_15_f1_mux_4_cse
      & butterFly1_15_f1_mux_5_cse & butterFly1_15_f1_mux_6_cse & butterFly1_15_f1_mux_7_cse));
  z_out_37 <= MUX1HOT_v_32_8_2(xt_rsc_0_19_i_qa_d, xt_rsc_1_19_i_qa_d, xt_rsc_2_19_i_qa_d,
      xt_rsc_3_19_i_qa_d, xt_rsc_4_19_i_qa_d, xt_rsc_5_19_i_qa_d, xt_rsc_6_19_i_qa_d,
      xt_rsc_7_19_i_qa_d, STD_LOGIC_VECTOR'( butterFly1_15_f1_mux_cse & butterFly1_15_f1_mux_1_cse
      & butterFly1_15_f1_mux_2_cse & butterFly1_15_f1_mux_3_cse & butterFly1_15_f1_mux_4_cse
      & butterFly1_15_f1_mux_5_cse & butterFly1_15_f1_mux_6_cse & butterFly1_15_f1_mux_7_cse));
  z_out_38 <= MUX1HOT_v_32_8_2(xt_rsc_0_21_i_qa_d, xt_rsc_1_21_i_qa_d, xt_rsc_2_21_i_qa_d,
      xt_rsc_3_21_i_qa_d, xt_rsc_4_21_i_qa_d, xt_rsc_5_21_i_qa_d, xt_rsc_6_21_i_qa_d,
      xt_rsc_7_21_i_qa_d, STD_LOGIC_VECTOR'( butterFly1_15_f1_mux_cse & butterFly1_15_f1_mux_1_cse
      & butterFly1_15_f1_mux_2_cse & butterFly1_15_f1_mux_3_cse & butterFly1_15_f1_mux_4_cse
      & butterFly1_15_f1_mux_5_cse & butterFly1_15_f1_mux_6_cse & butterFly1_15_f1_mux_7_cse));
  z_out_39 <= MUX1HOT_v_32_8_2(xt_rsc_0_23_i_qa_d, xt_rsc_1_23_i_qa_d, xt_rsc_2_23_i_qa_d,
      xt_rsc_3_23_i_qa_d, xt_rsc_4_23_i_qa_d, xt_rsc_5_23_i_qa_d, xt_rsc_6_23_i_qa_d,
      xt_rsc_7_23_i_qa_d, STD_LOGIC_VECTOR'( butterFly1_15_f1_mux_cse & butterFly1_15_f1_mux_1_cse
      & butterFly1_15_f1_mux_2_cse & butterFly1_15_f1_mux_3_cse & butterFly1_15_f1_mux_4_cse
      & butterFly1_15_f1_mux_5_cse & butterFly1_15_f1_mux_6_cse & butterFly1_15_f1_mux_7_cse));
  z_out_40 <= MUX1HOT_v_32_8_2(xt_rsc_0_25_i_qa_d, xt_rsc_1_25_i_qa_d, xt_rsc_2_25_i_qa_d,
      xt_rsc_3_25_i_qa_d, xt_rsc_4_25_i_qa_d, xt_rsc_5_25_i_qa_d, xt_rsc_6_25_i_qa_d,
      xt_rsc_7_25_i_qa_d, STD_LOGIC_VECTOR'( butterFly1_15_f1_mux_cse & butterFly1_15_f1_mux_1_cse
      & butterFly1_15_f1_mux_2_cse & butterFly1_15_f1_mux_3_cse & butterFly1_15_f1_mux_4_cse
      & butterFly1_15_f1_mux_5_cse & butterFly1_15_f1_mux_6_cse & butterFly1_15_f1_mux_7_cse));
  z_out_41 <= MUX1HOT_v_32_8_2(xt_rsc_0_27_i_qa_d, xt_rsc_1_27_i_qa_d, xt_rsc_2_27_i_qa_d,
      xt_rsc_3_27_i_qa_d, xt_rsc_4_27_i_qa_d, xt_rsc_5_27_i_qa_d, xt_rsc_6_27_i_qa_d,
      xt_rsc_7_27_i_qa_d, STD_LOGIC_VECTOR'( butterFly1_15_f1_mux_cse & butterFly1_15_f1_mux_1_cse
      & butterFly1_15_f1_mux_2_cse & butterFly1_15_f1_mux_3_cse & butterFly1_15_f1_mux_4_cse
      & butterFly1_15_f1_mux_5_cse & butterFly1_15_f1_mux_6_cse & butterFly1_15_f1_mux_7_cse));
  z_out_42 <= MUX1HOT_v_32_8_2(xt_rsc_0_29_i_qa_d, xt_rsc_1_29_i_qa_d, xt_rsc_2_29_i_qa_d,
      xt_rsc_3_29_i_qa_d, xt_rsc_4_29_i_qa_d, xt_rsc_5_29_i_qa_d, xt_rsc_6_29_i_qa_d,
      xt_rsc_7_29_i_qa_d, STD_LOGIC_VECTOR'( butterFly1_15_f1_mux_cse & butterFly1_15_f1_mux_1_cse
      & butterFly1_15_f1_mux_2_cse & butterFly1_15_f1_mux_3_cse & butterFly1_15_f1_mux_4_cse
      & butterFly1_15_f1_mux_5_cse & butterFly1_15_f1_mux_6_cse & butterFly1_15_f1_mux_7_cse));
  z_out_43 <= MUX1HOT_v_32_8_2(xt_rsc_0_1_i_qa_d, xt_rsc_1_1_i_qa_d, xt_rsc_2_1_i_qa_d,
      xt_rsc_3_1_i_qa_d, xt_rsc_4_1_i_qa_d, xt_rsc_5_1_i_qa_d, xt_rsc_6_1_i_qa_d,
      xt_rsc_7_1_i_qa_d, STD_LOGIC_VECTOR'( butterFly2_f1_mux_cse & butterFly2_f1_mux_1_cse
      & butterFly2_f1_mux_2_cse & butterFly2_f1_mux_3_cse & butterFly2_f1_mux_4_cse
      & butterFly2_f1_mux_5_cse & butterFly2_f1_mux_6_cse & butterFly2_f1_mux_7_cse));
  z_out_44 <= MUX1HOT_v_32_8_2(xt_rsc_0_3_i_qa_d, xt_rsc_1_3_i_qa_d, xt_rsc_2_3_i_qa_d,
      xt_rsc_3_3_i_qa_d, xt_rsc_4_3_i_qa_d, xt_rsc_5_3_i_qa_d, xt_rsc_6_3_i_qa_d,
      xt_rsc_7_3_i_qa_d, STD_LOGIC_VECTOR'( butterFly2_f1_mux_cse & butterFly2_f1_mux_1_cse
      & butterFly2_f1_mux_2_cse & butterFly2_f1_mux_3_cse & butterFly2_f1_mux_4_cse
      & butterFly2_f1_mux_5_cse & butterFly2_f1_mux_6_cse & butterFly2_f1_mux_7_cse));
  z_out_45 <= MUX1HOT_v_32_8_2(xt_rsc_0_5_i_qa_d, xt_rsc_1_5_i_qa_d, xt_rsc_2_5_i_qa_d,
      xt_rsc_3_5_i_qa_d, xt_rsc_4_5_i_qa_d, xt_rsc_5_5_i_qa_d, xt_rsc_6_5_i_qa_d,
      xt_rsc_7_5_i_qa_d, STD_LOGIC_VECTOR'( butterFly2_f1_mux_cse & butterFly2_f1_mux_1_cse
      & butterFly2_f1_mux_2_cse & butterFly2_f1_mux_3_cse & butterFly2_f1_mux_4_cse
      & butterFly2_f1_mux_5_cse & butterFly2_f1_mux_6_cse & butterFly2_f1_mux_7_cse));
  z_out_46 <= MUX1HOT_v_32_8_2(xt_rsc_0_13_i_qa_d, xt_rsc_1_13_i_qa_d, xt_rsc_2_13_i_qa_d,
      xt_rsc_3_13_i_qa_d, xt_rsc_4_13_i_qa_d, xt_rsc_5_13_i_qa_d, xt_rsc_6_13_i_qa_d,
      xt_rsc_7_13_i_qa_d, STD_LOGIC_VECTOR'( butterFly2_f1_mux_cse & butterFly2_f1_mux_1_cse
      & butterFly2_f1_mux_2_cse & butterFly2_f1_mux_3_cse & butterFly2_f1_mux_4_cse
      & butterFly2_f1_mux_5_cse & butterFly2_f1_mux_6_cse & butterFly2_f1_mux_7_cse));
  z_out_47 <= MUX1HOT_v_32_8_2(xt_rsc_0_15_i_qa_d, xt_rsc_1_15_i_qa_d, xt_rsc_2_15_i_qa_d,
      xt_rsc_3_15_i_qa_d, xt_rsc_4_15_i_qa_d, xt_rsc_5_15_i_qa_d, xt_rsc_6_15_i_qa_d,
      xt_rsc_7_15_i_qa_d, STD_LOGIC_VECTOR'( butterFly2_f1_mux_cse & butterFly2_f1_mux_1_cse
      & butterFly2_f1_mux_2_cse & butterFly2_f1_mux_3_cse & butterFly2_f1_mux_4_cse
      & butterFly2_f1_mux_5_cse & butterFly2_f1_mux_6_cse & butterFly2_f1_mux_7_cse));
  z_out_48 <= MUX1HOT_v_32_8_2(xt_rsc_0_17_i_qa_d, xt_rsc_1_17_i_qa_d, xt_rsc_2_17_i_qa_d,
      xt_rsc_3_17_i_qa_d, xt_rsc_4_17_i_qa_d, xt_rsc_5_17_i_qa_d, xt_rsc_6_17_i_qa_d,
      xt_rsc_7_17_i_qa_d, STD_LOGIC_VECTOR'( butterFly2_f1_mux_cse & butterFly2_f1_mux_1_cse
      & butterFly2_f1_mux_2_cse & butterFly2_f1_mux_3_cse & butterFly2_f1_mux_4_cse
      & butterFly2_f1_mux_5_cse & butterFly2_f1_mux_6_cse & butterFly2_f1_mux_7_cse));
  z_out_49 <= MUX1HOT_v_32_8_2(xt_rsc_0_31_i_qa_d, xt_rsc_1_31_i_qa_d, xt_rsc_2_31_i_qa_d,
      xt_rsc_3_31_i_qa_d, xt_rsc_4_31_i_qa_d, xt_rsc_5_31_i_qa_d, xt_rsc_6_31_i_qa_d,
      xt_rsc_7_31_i_qa_d, STD_LOGIC_VECTOR'( butterFly2_f1_mux_cse & butterFly2_f1_mux_1_cse
      & butterFly2_f1_mux_2_cse & butterFly2_f1_mux_3_cse & butterFly2_f1_mux_4_cse
      & butterFly2_f1_mux_5_cse & butterFly2_f1_mux_6_cse & butterFly2_f1_mux_7_cse));
  z_out_50 <= MUX1HOT_v_32_8_2(yt_rsc_0_29_i_q_d, yt_rsc_1_29_i_q_d, yt_rsc_2_29_i_q_d,
      yt_rsc_3_29_i_q_d, yt_rsc_4_29_i_q_d, yt_rsc_5_29_i_q_d, yt_rsc_6_29_i_q_d,
      yt_rsc_7_29_i_q_d, STD_LOGIC_VECTOR'( butterFly1_31_f1_mux_cse & butterFly1_31_f1_mux_1_cse
      & butterFly1_31_f1_mux_2_cse & butterFly1_31_f1_mux_3_cse & butterFly1_31_f1_mux_4_cse
      & butterFly1_31_f1_mux_5_cse & butterFly1_31_f1_mux_6_cse & butterFly1_31_f1_mux_7_cse));
  z_out_51 <= MUX1HOT_v_32_8_2(yt_rsc_0_27_i_q_d, yt_rsc_1_27_i_q_d, yt_rsc_2_27_i_q_d,
      yt_rsc_3_27_i_q_d, yt_rsc_4_27_i_q_d, yt_rsc_5_27_i_q_d, yt_rsc_6_27_i_q_d,
      yt_rsc_7_27_i_q_d, STD_LOGIC_VECTOR'( butterFly1_31_f1_mux_cse & butterFly1_31_f1_mux_1_cse
      & butterFly1_31_f1_mux_2_cse & butterFly1_31_f1_mux_3_cse & butterFly1_31_f1_mux_4_cse
      & butterFly1_31_f1_mux_5_cse & butterFly1_31_f1_mux_6_cse & butterFly1_31_f1_mux_7_cse));
  z_out_52 <= MUX1HOT_v_32_8_2(yt_rsc_0_25_i_q_d, yt_rsc_1_25_i_q_d, yt_rsc_2_25_i_q_d,
      yt_rsc_3_25_i_q_d, yt_rsc_4_25_i_q_d, yt_rsc_5_25_i_q_d, yt_rsc_6_25_i_q_d,
      yt_rsc_7_25_i_q_d, STD_LOGIC_VECTOR'( butterFly1_31_f1_mux_cse & butterFly1_31_f1_mux_1_cse
      & butterFly1_31_f1_mux_2_cse & butterFly1_31_f1_mux_3_cse & butterFly1_31_f1_mux_4_cse
      & butterFly1_31_f1_mux_5_cse & butterFly1_31_f1_mux_6_cse & butterFly1_31_f1_mux_7_cse));
  z_out_53 <= MUX1HOT_v_32_8_2(yt_rsc_0_21_i_q_d, yt_rsc_1_21_i_q_d, yt_rsc_2_21_i_q_d,
      yt_rsc_3_21_i_q_d, yt_rsc_4_21_i_q_d, yt_rsc_5_21_i_q_d, yt_rsc_6_21_i_q_d,
      yt_rsc_7_21_i_q_d, STD_LOGIC_VECTOR'( butterFly1_31_f1_mux_cse & butterFly1_31_f1_mux_1_cse
      & butterFly1_31_f1_mux_2_cse & butterFly1_31_f1_mux_3_cse & butterFly1_31_f1_mux_4_cse
      & butterFly1_31_f1_mux_5_cse & butterFly1_31_f1_mux_6_cse & butterFly1_31_f1_mux_7_cse));
  z_out_54 <= MUX1HOT_v_32_8_2(yt_rsc_0_11_i_q_d, yt_rsc_1_11_i_q_d, yt_rsc_2_11_i_q_d,
      yt_rsc_3_11_i_q_d, yt_rsc_4_11_i_q_d, yt_rsc_5_11_i_q_d, yt_rsc_6_11_i_q_d,
      yt_rsc_7_11_i_q_d, STD_LOGIC_VECTOR'( butterFly2_21_f1_mux_cse & butterFly2_21_f1_mux_1_cse
      & butterFly2_21_f1_mux_2_cse & butterFly2_21_f1_mux_3_cse & butterFly2_21_f1_mux_4_cse
      & butterFly2_21_f1_mux_5_cse & butterFly2_21_f1_mux_6_cse & butterFly2_21_f1_mux_7_cse));
  z_out_55 <= MUX1HOT_v_32_8_2(yt_rsc_0_19_i_q_d, yt_rsc_1_19_i_q_d, yt_rsc_2_19_i_q_d,
      yt_rsc_3_19_i_q_d, yt_rsc_4_19_i_q_d, yt_rsc_5_19_i_q_d, yt_rsc_6_19_i_q_d,
      yt_rsc_7_19_i_q_d, STD_LOGIC_VECTOR'( butterFly1_31_f1_mux_cse & butterFly1_31_f1_mux_1_cse
      & butterFly1_31_f1_mux_2_cse & butterFly1_31_f1_mux_3_cse & butterFly1_31_f1_mux_4_cse
      & butterFly1_31_f1_mux_5_cse & butterFly1_31_f1_mux_6_cse & butterFly1_31_f1_mux_7_cse));
  z_out_56 <= MUX1HOT_v_32_8_2(yt_rsc_0_13_i_q_d, yt_rsc_1_13_i_q_d, yt_rsc_2_13_i_q_d,
      yt_rsc_3_13_i_q_d, yt_rsc_4_13_i_q_d, yt_rsc_5_13_i_q_d, yt_rsc_6_13_i_q_d,
      yt_rsc_7_13_i_q_d, STD_LOGIC_VECTOR'( butterFly2_21_f1_mux_cse & butterFly2_21_f1_mux_1_cse
      & butterFly2_21_f1_mux_2_cse & butterFly2_21_f1_mux_3_cse & butterFly2_21_f1_mux_4_cse
      & butterFly2_21_f1_mux_5_cse & butterFly2_21_f1_mux_6_cse & butterFly2_21_f1_mux_7_cse));
  z_out_57 <= MUX1HOT_v_32_8_2(yt_rsc_0_17_i_q_d, yt_rsc_1_17_i_q_d, yt_rsc_2_17_i_q_d,
      yt_rsc_3_17_i_q_d, yt_rsc_4_17_i_q_d, yt_rsc_5_17_i_q_d, yt_rsc_6_17_i_q_d,
      yt_rsc_7_17_i_q_d, STD_LOGIC_VECTOR'( butterFly1_31_f1_mux_cse & butterFly1_31_f1_mux_1_cse
      & butterFly1_31_f1_mux_2_cse & butterFly1_31_f1_mux_3_cse & butterFly1_31_f1_mux_4_cse
      & butterFly1_31_f1_mux_5_cse & butterFly1_31_f1_mux_6_cse & butterFly1_31_f1_mux_7_cse));
  z_out_58 <= MUX1HOT_v_32_8_2(yt_rsc_0_15_i_q_d, yt_rsc_1_15_i_q_d, yt_rsc_2_15_i_q_d,
      yt_rsc_3_15_i_q_d, yt_rsc_4_15_i_q_d, yt_rsc_5_15_i_q_d, yt_rsc_6_15_i_q_d,
      yt_rsc_7_15_i_q_d, STD_LOGIC_VECTOR'( butterFly2_21_f1_mux_cse & butterFly2_21_f1_mux_1_cse
      & butterFly2_21_f1_mux_2_cse & butterFly2_21_f1_mux_3_cse & butterFly2_21_f1_mux_4_cse
      & butterFly2_21_f1_mux_5_cse & butterFly2_21_f1_mux_6_cse & butterFly2_21_f1_mux_7_cse));
  z_out_59 <= MUX1HOT_v_32_8_2(yt_rsc_0_1_i_q_d, yt_rsc_1_1_i_q_d, yt_rsc_2_1_i_q_d,
      yt_rsc_3_1_i_q_d, yt_rsc_4_1_i_q_d, yt_rsc_5_1_i_q_d, yt_rsc_6_1_i_q_d, yt_rsc_7_1_i_q_d,
      STD_LOGIC_VECTOR'( butterFly1_31_f1_mux_cse & butterFly1_31_f1_mux_1_cse &
      butterFly1_31_f1_mux_2_cse & butterFly1_31_f1_mux_3_cse & butterFly1_31_f1_mux_4_cse
      & butterFly1_31_f1_mux_5_cse & butterFly1_31_f1_mux_6_cse & butterFly1_31_f1_mux_7_cse));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_1R1W_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_0_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_0_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_0_wea : OUT STD_LOGIC;
    xt_rsc_0_0_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_0_lz : OUT STD_LOGIC;
    xt_rsc_0_1_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_1_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_1_wea : OUT STD_LOGIC;
    xt_rsc_0_1_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_1_lz : OUT STD_LOGIC;
    xt_rsc_0_2_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_2_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_2_wea : OUT STD_LOGIC;
    xt_rsc_0_2_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_2_lz : OUT STD_LOGIC;
    xt_rsc_0_3_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_3_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_3_wea : OUT STD_LOGIC;
    xt_rsc_0_3_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_3_lz : OUT STD_LOGIC;
    xt_rsc_0_4_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_4_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_4_wea : OUT STD_LOGIC;
    xt_rsc_0_4_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_4_lz : OUT STD_LOGIC;
    xt_rsc_0_5_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_5_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_5_wea : OUT STD_LOGIC;
    xt_rsc_0_5_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_5_lz : OUT STD_LOGIC;
    xt_rsc_0_6_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_6_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_6_wea : OUT STD_LOGIC;
    xt_rsc_0_6_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_6_lz : OUT STD_LOGIC;
    xt_rsc_0_7_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_7_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_7_wea : OUT STD_LOGIC;
    xt_rsc_0_7_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_7_lz : OUT STD_LOGIC;
    xt_rsc_0_8_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_8_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_8_wea : OUT STD_LOGIC;
    xt_rsc_0_8_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_8_lz : OUT STD_LOGIC;
    xt_rsc_0_9_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_9_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_9_wea : OUT STD_LOGIC;
    xt_rsc_0_9_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_9_lz : OUT STD_LOGIC;
    xt_rsc_0_10_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_10_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_10_wea : OUT STD_LOGIC;
    xt_rsc_0_10_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_10_lz : OUT STD_LOGIC;
    xt_rsc_0_11_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_11_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_11_wea : OUT STD_LOGIC;
    xt_rsc_0_11_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_11_lz : OUT STD_LOGIC;
    xt_rsc_0_12_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_12_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_12_wea : OUT STD_LOGIC;
    xt_rsc_0_12_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_12_lz : OUT STD_LOGIC;
    xt_rsc_0_13_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_13_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_13_wea : OUT STD_LOGIC;
    xt_rsc_0_13_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_13_lz : OUT STD_LOGIC;
    xt_rsc_0_14_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_14_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_14_wea : OUT STD_LOGIC;
    xt_rsc_0_14_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_14_lz : OUT STD_LOGIC;
    xt_rsc_0_15_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_15_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_15_wea : OUT STD_LOGIC;
    xt_rsc_0_15_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_15_lz : OUT STD_LOGIC;
    xt_rsc_0_16_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_16_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_16_wea : OUT STD_LOGIC;
    xt_rsc_0_16_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_16_lz : OUT STD_LOGIC;
    xt_rsc_0_17_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_17_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_17_wea : OUT STD_LOGIC;
    xt_rsc_0_17_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_17_lz : OUT STD_LOGIC;
    xt_rsc_0_18_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_18_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_18_wea : OUT STD_LOGIC;
    xt_rsc_0_18_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_18_lz : OUT STD_LOGIC;
    xt_rsc_0_19_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_19_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_19_wea : OUT STD_LOGIC;
    xt_rsc_0_19_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_19_lz : OUT STD_LOGIC;
    xt_rsc_0_20_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_20_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_20_wea : OUT STD_LOGIC;
    xt_rsc_0_20_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_20_lz : OUT STD_LOGIC;
    xt_rsc_0_21_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_21_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_21_wea : OUT STD_LOGIC;
    xt_rsc_0_21_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_21_lz : OUT STD_LOGIC;
    xt_rsc_0_22_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_22_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_22_wea : OUT STD_LOGIC;
    xt_rsc_0_22_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_22_lz : OUT STD_LOGIC;
    xt_rsc_0_23_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_23_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_23_wea : OUT STD_LOGIC;
    xt_rsc_0_23_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_23_lz : OUT STD_LOGIC;
    xt_rsc_0_24_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_24_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_24_wea : OUT STD_LOGIC;
    xt_rsc_0_24_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_24_lz : OUT STD_LOGIC;
    xt_rsc_0_25_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_25_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_25_wea : OUT STD_LOGIC;
    xt_rsc_0_25_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_25_lz : OUT STD_LOGIC;
    xt_rsc_0_26_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_26_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_26_wea : OUT STD_LOGIC;
    xt_rsc_0_26_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_26_lz : OUT STD_LOGIC;
    xt_rsc_0_27_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_27_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_27_wea : OUT STD_LOGIC;
    xt_rsc_0_27_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_27_lz : OUT STD_LOGIC;
    xt_rsc_0_28_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_28_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_28_wea : OUT STD_LOGIC;
    xt_rsc_0_28_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_28_lz : OUT STD_LOGIC;
    xt_rsc_0_29_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_29_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_29_wea : OUT STD_LOGIC;
    xt_rsc_0_29_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_29_lz : OUT STD_LOGIC;
    xt_rsc_0_30_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_30_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_30_wea : OUT STD_LOGIC;
    xt_rsc_0_30_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_30_lz : OUT STD_LOGIC;
    xt_rsc_0_31_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_31_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_31_wea : OUT STD_LOGIC;
    xt_rsc_0_31_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_31_lz : OUT STD_LOGIC;
    xt_rsc_1_0_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_1_0_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_0_wea : OUT STD_LOGIC;
    xt_rsc_1_0_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_1_0_lz : OUT STD_LOGIC;
    xt_rsc_1_1_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_1_1_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_1_wea : OUT STD_LOGIC;
    xt_rsc_1_1_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_1_1_lz : OUT STD_LOGIC;
    xt_rsc_1_2_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_1_2_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_2_wea : OUT STD_LOGIC;
    xt_rsc_1_2_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_1_2_lz : OUT STD_LOGIC;
    xt_rsc_1_3_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_1_3_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_3_wea : OUT STD_LOGIC;
    xt_rsc_1_3_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_1_3_lz : OUT STD_LOGIC;
    xt_rsc_1_4_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_1_4_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_4_wea : OUT STD_LOGIC;
    xt_rsc_1_4_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_1_4_lz : OUT STD_LOGIC;
    xt_rsc_1_5_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_1_5_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_5_wea : OUT STD_LOGIC;
    xt_rsc_1_5_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_1_5_lz : OUT STD_LOGIC;
    xt_rsc_1_6_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_1_6_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_6_wea : OUT STD_LOGIC;
    xt_rsc_1_6_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_1_6_lz : OUT STD_LOGIC;
    xt_rsc_1_7_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_1_7_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_7_wea : OUT STD_LOGIC;
    xt_rsc_1_7_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_1_7_lz : OUT STD_LOGIC;
    xt_rsc_1_8_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_1_8_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_8_wea : OUT STD_LOGIC;
    xt_rsc_1_8_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_1_8_lz : OUT STD_LOGIC;
    xt_rsc_1_9_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_1_9_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_9_wea : OUT STD_LOGIC;
    xt_rsc_1_9_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_1_9_lz : OUT STD_LOGIC;
    xt_rsc_1_10_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_1_10_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_10_wea : OUT STD_LOGIC;
    xt_rsc_1_10_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_1_10_lz : OUT STD_LOGIC;
    xt_rsc_1_11_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_1_11_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_11_wea : OUT STD_LOGIC;
    xt_rsc_1_11_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_1_11_lz : OUT STD_LOGIC;
    xt_rsc_1_12_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_1_12_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_12_wea : OUT STD_LOGIC;
    xt_rsc_1_12_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_1_12_lz : OUT STD_LOGIC;
    xt_rsc_1_13_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_1_13_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_13_wea : OUT STD_LOGIC;
    xt_rsc_1_13_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_1_13_lz : OUT STD_LOGIC;
    xt_rsc_1_14_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_1_14_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_14_wea : OUT STD_LOGIC;
    xt_rsc_1_14_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_1_14_lz : OUT STD_LOGIC;
    xt_rsc_1_15_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_1_15_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_15_wea : OUT STD_LOGIC;
    xt_rsc_1_15_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_1_15_lz : OUT STD_LOGIC;
    xt_rsc_1_16_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_1_16_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_16_wea : OUT STD_LOGIC;
    xt_rsc_1_16_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_1_16_lz : OUT STD_LOGIC;
    xt_rsc_1_17_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_1_17_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_17_wea : OUT STD_LOGIC;
    xt_rsc_1_17_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_1_17_lz : OUT STD_LOGIC;
    xt_rsc_1_18_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_1_18_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_18_wea : OUT STD_LOGIC;
    xt_rsc_1_18_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_1_18_lz : OUT STD_LOGIC;
    xt_rsc_1_19_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_1_19_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_19_wea : OUT STD_LOGIC;
    xt_rsc_1_19_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_1_19_lz : OUT STD_LOGIC;
    xt_rsc_1_20_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_1_20_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_20_wea : OUT STD_LOGIC;
    xt_rsc_1_20_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_1_20_lz : OUT STD_LOGIC;
    xt_rsc_1_21_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_1_21_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_21_wea : OUT STD_LOGIC;
    xt_rsc_1_21_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_1_21_lz : OUT STD_LOGIC;
    xt_rsc_1_22_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_1_22_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_22_wea : OUT STD_LOGIC;
    xt_rsc_1_22_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_1_22_lz : OUT STD_LOGIC;
    xt_rsc_1_23_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_1_23_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_23_wea : OUT STD_LOGIC;
    xt_rsc_1_23_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_1_23_lz : OUT STD_LOGIC;
    xt_rsc_1_24_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_1_24_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_24_wea : OUT STD_LOGIC;
    xt_rsc_1_24_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_1_24_lz : OUT STD_LOGIC;
    xt_rsc_1_25_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_1_25_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_25_wea : OUT STD_LOGIC;
    xt_rsc_1_25_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_1_25_lz : OUT STD_LOGIC;
    xt_rsc_1_26_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_1_26_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_26_wea : OUT STD_LOGIC;
    xt_rsc_1_26_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_1_26_lz : OUT STD_LOGIC;
    xt_rsc_1_27_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_1_27_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_27_wea : OUT STD_LOGIC;
    xt_rsc_1_27_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_1_27_lz : OUT STD_LOGIC;
    xt_rsc_1_28_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_1_28_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_28_wea : OUT STD_LOGIC;
    xt_rsc_1_28_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_1_28_lz : OUT STD_LOGIC;
    xt_rsc_1_29_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_1_29_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_29_wea : OUT STD_LOGIC;
    xt_rsc_1_29_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_1_29_lz : OUT STD_LOGIC;
    xt_rsc_1_30_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_1_30_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_30_wea : OUT STD_LOGIC;
    xt_rsc_1_30_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_1_30_lz : OUT STD_LOGIC;
    xt_rsc_1_31_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_1_31_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_31_wea : OUT STD_LOGIC;
    xt_rsc_1_31_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_1_31_lz : OUT STD_LOGIC;
    xt_rsc_2_0_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_2_0_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_2_0_wea : OUT STD_LOGIC;
    xt_rsc_2_0_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_2_0_lz : OUT STD_LOGIC;
    xt_rsc_2_1_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_2_1_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_2_1_wea : OUT STD_LOGIC;
    xt_rsc_2_1_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_2_1_lz : OUT STD_LOGIC;
    xt_rsc_2_2_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_2_2_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_2_2_wea : OUT STD_LOGIC;
    xt_rsc_2_2_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_2_2_lz : OUT STD_LOGIC;
    xt_rsc_2_3_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_2_3_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_2_3_wea : OUT STD_LOGIC;
    xt_rsc_2_3_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_2_3_lz : OUT STD_LOGIC;
    xt_rsc_2_4_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_2_4_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_2_4_wea : OUT STD_LOGIC;
    xt_rsc_2_4_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_2_4_lz : OUT STD_LOGIC;
    xt_rsc_2_5_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_2_5_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_2_5_wea : OUT STD_LOGIC;
    xt_rsc_2_5_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_2_5_lz : OUT STD_LOGIC;
    xt_rsc_2_6_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_2_6_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_2_6_wea : OUT STD_LOGIC;
    xt_rsc_2_6_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_2_6_lz : OUT STD_LOGIC;
    xt_rsc_2_7_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_2_7_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_2_7_wea : OUT STD_LOGIC;
    xt_rsc_2_7_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_2_7_lz : OUT STD_LOGIC;
    xt_rsc_2_8_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_2_8_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_2_8_wea : OUT STD_LOGIC;
    xt_rsc_2_8_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_2_8_lz : OUT STD_LOGIC;
    xt_rsc_2_9_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_2_9_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_2_9_wea : OUT STD_LOGIC;
    xt_rsc_2_9_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_2_9_lz : OUT STD_LOGIC;
    xt_rsc_2_10_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_2_10_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_2_10_wea : OUT STD_LOGIC;
    xt_rsc_2_10_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_2_10_lz : OUT STD_LOGIC;
    xt_rsc_2_11_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_2_11_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_2_11_wea : OUT STD_LOGIC;
    xt_rsc_2_11_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_2_11_lz : OUT STD_LOGIC;
    xt_rsc_2_12_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_2_12_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_2_12_wea : OUT STD_LOGIC;
    xt_rsc_2_12_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_2_12_lz : OUT STD_LOGIC;
    xt_rsc_2_13_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_2_13_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_2_13_wea : OUT STD_LOGIC;
    xt_rsc_2_13_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_2_13_lz : OUT STD_LOGIC;
    xt_rsc_2_14_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_2_14_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_2_14_wea : OUT STD_LOGIC;
    xt_rsc_2_14_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_2_14_lz : OUT STD_LOGIC;
    xt_rsc_2_15_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_2_15_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_2_15_wea : OUT STD_LOGIC;
    xt_rsc_2_15_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_2_15_lz : OUT STD_LOGIC;
    xt_rsc_2_16_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_2_16_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_2_16_wea : OUT STD_LOGIC;
    xt_rsc_2_16_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_2_16_lz : OUT STD_LOGIC;
    xt_rsc_2_17_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_2_17_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_2_17_wea : OUT STD_LOGIC;
    xt_rsc_2_17_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_2_17_lz : OUT STD_LOGIC;
    xt_rsc_2_18_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_2_18_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_2_18_wea : OUT STD_LOGIC;
    xt_rsc_2_18_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_2_18_lz : OUT STD_LOGIC;
    xt_rsc_2_19_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_2_19_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_2_19_wea : OUT STD_LOGIC;
    xt_rsc_2_19_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_2_19_lz : OUT STD_LOGIC;
    xt_rsc_2_20_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_2_20_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_2_20_wea : OUT STD_LOGIC;
    xt_rsc_2_20_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_2_20_lz : OUT STD_LOGIC;
    xt_rsc_2_21_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_2_21_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_2_21_wea : OUT STD_LOGIC;
    xt_rsc_2_21_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_2_21_lz : OUT STD_LOGIC;
    xt_rsc_2_22_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_2_22_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_2_22_wea : OUT STD_LOGIC;
    xt_rsc_2_22_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_2_22_lz : OUT STD_LOGIC;
    xt_rsc_2_23_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_2_23_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_2_23_wea : OUT STD_LOGIC;
    xt_rsc_2_23_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_2_23_lz : OUT STD_LOGIC;
    xt_rsc_2_24_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_2_24_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_2_24_wea : OUT STD_LOGIC;
    xt_rsc_2_24_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_2_24_lz : OUT STD_LOGIC;
    xt_rsc_2_25_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_2_25_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_2_25_wea : OUT STD_LOGIC;
    xt_rsc_2_25_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_2_25_lz : OUT STD_LOGIC;
    xt_rsc_2_26_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_2_26_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_2_26_wea : OUT STD_LOGIC;
    xt_rsc_2_26_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_2_26_lz : OUT STD_LOGIC;
    xt_rsc_2_27_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_2_27_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_2_27_wea : OUT STD_LOGIC;
    xt_rsc_2_27_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_2_27_lz : OUT STD_LOGIC;
    xt_rsc_2_28_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_2_28_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_2_28_wea : OUT STD_LOGIC;
    xt_rsc_2_28_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_2_28_lz : OUT STD_LOGIC;
    xt_rsc_2_29_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_2_29_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_2_29_wea : OUT STD_LOGIC;
    xt_rsc_2_29_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_2_29_lz : OUT STD_LOGIC;
    xt_rsc_2_30_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_2_30_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_2_30_wea : OUT STD_LOGIC;
    xt_rsc_2_30_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_2_30_lz : OUT STD_LOGIC;
    xt_rsc_2_31_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_2_31_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_2_31_wea : OUT STD_LOGIC;
    xt_rsc_2_31_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_2_31_lz : OUT STD_LOGIC;
    xt_rsc_3_0_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_3_0_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_3_0_wea : OUT STD_LOGIC;
    xt_rsc_3_0_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_3_0_lz : OUT STD_LOGIC;
    xt_rsc_3_1_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_3_1_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_3_1_wea : OUT STD_LOGIC;
    xt_rsc_3_1_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_3_1_lz : OUT STD_LOGIC;
    xt_rsc_3_2_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_3_2_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_3_2_wea : OUT STD_LOGIC;
    xt_rsc_3_2_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_3_2_lz : OUT STD_LOGIC;
    xt_rsc_3_3_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_3_3_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_3_3_wea : OUT STD_LOGIC;
    xt_rsc_3_3_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_3_3_lz : OUT STD_LOGIC;
    xt_rsc_3_4_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_3_4_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_3_4_wea : OUT STD_LOGIC;
    xt_rsc_3_4_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_3_4_lz : OUT STD_LOGIC;
    xt_rsc_3_5_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_3_5_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_3_5_wea : OUT STD_LOGIC;
    xt_rsc_3_5_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_3_5_lz : OUT STD_LOGIC;
    xt_rsc_3_6_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_3_6_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_3_6_wea : OUT STD_LOGIC;
    xt_rsc_3_6_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_3_6_lz : OUT STD_LOGIC;
    xt_rsc_3_7_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_3_7_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_3_7_wea : OUT STD_LOGIC;
    xt_rsc_3_7_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_3_7_lz : OUT STD_LOGIC;
    xt_rsc_3_8_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_3_8_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_3_8_wea : OUT STD_LOGIC;
    xt_rsc_3_8_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_3_8_lz : OUT STD_LOGIC;
    xt_rsc_3_9_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_3_9_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_3_9_wea : OUT STD_LOGIC;
    xt_rsc_3_9_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_3_9_lz : OUT STD_LOGIC;
    xt_rsc_3_10_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_3_10_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_3_10_wea : OUT STD_LOGIC;
    xt_rsc_3_10_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_3_10_lz : OUT STD_LOGIC;
    xt_rsc_3_11_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_3_11_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_3_11_wea : OUT STD_LOGIC;
    xt_rsc_3_11_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_3_11_lz : OUT STD_LOGIC;
    xt_rsc_3_12_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_3_12_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_3_12_wea : OUT STD_LOGIC;
    xt_rsc_3_12_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_3_12_lz : OUT STD_LOGIC;
    xt_rsc_3_13_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_3_13_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_3_13_wea : OUT STD_LOGIC;
    xt_rsc_3_13_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_3_13_lz : OUT STD_LOGIC;
    xt_rsc_3_14_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_3_14_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_3_14_wea : OUT STD_LOGIC;
    xt_rsc_3_14_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_3_14_lz : OUT STD_LOGIC;
    xt_rsc_3_15_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_3_15_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_3_15_wea : OUT STD_LOGIC;
    xt_rsc_3_15_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_3_15_lz : OUT STD_LOGIC;
    xt_rsc_3_16_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_3_16_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_3_16_wea : OUT STD_LOGIC;
    xt_rsc_3_16_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_3_16_lz : OUT STD_LOGIC;
    xt_rsc_3_17_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_3_17_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_3_17_wea : OUT STD_LOGIC;
    xt_rsc_3_17_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_3_17_lz : OUT STD_LOGIC;
    xt_rsc_3_18_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_3_18_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_3_18_wea : OUT STD_LOGIC;
    xt_rsc_3_18_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_3_18_lz : OUT STD_LOGIC;
    xt_rsc_3_19_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_3_19_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_3_19_wea : OUT STD_LOGIC;
    xt_rsc_3_19_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_3_19_lz : OUT STD_LOGIC;
    xt_rsc_3_20_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_3_20_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_3_20_wea : OUT STD_LOGIC;
    xt_rsc_3_20_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_3_20_lz : OUT STD_LOGIC;
    xt_rsc_3_21_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_3_21_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_3_21_wea : OUT STD_LOGIC;
    xt_rsc_3_21_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_3_21_lz : OUT STD_LOGIC;
    xt_rsc_3_22_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_3_22_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_3_22_wea : OUT STD_LOGIC;
    xt_rsc_3_22_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_3_22_lz : OUT STD_LOGIC;
    xt_rsc_3_23_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_3_23_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_3_23_wea : OUT STD_LOGIC;
    xt_rsc_3_23_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_3_23_lz : OUT STD_LOGIC;
    xt_rsc_3_24_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_3_24_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_3_24_wea : OUT STD_LOGIC;
    xt_rsc_3_24_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_3_24_lz : OUT STD_LOGIC;
    xt_rsc_3_25_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_3_25_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_3_25_wea : OUT STD_LOGIC;
    xt_rsc_3_25_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_3_25_lz : OUT STD_LOGIC;
    xt_rsc_3_26_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_3_26_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_3_26_wea : OUT STD_LOGIC;
    xt_rsc_3_26_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_3_26_lz : OUT STD_LOGIC;
    xt_rsc_3_27_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_3_27_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_3_27_wea : OUT STD_LOGIC;
    xt_rsc_3_27_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_3_27_lz : OUT STD_LOGIC;
    xt_rsc_3_28_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_3_28_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_3_28_wea : OUT STD_LOGIC;
    xt_rsc_3_28_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_3_28_lz : OUT STD_LOGIC;
    xt_rsc_3_29_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_3_29_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_3_29_wea : OUT STD_LOGIC;
    xt_rsc_3_29_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_3_29_lz : OUT STD_LOGIC;
    xt_rsc_3_30_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_3_30_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_3_30_wea : OUT STD_LOGIC;
    xt_rsc_3_30_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_3_30_lz : OUT STD_LOGIC;
    xt_rsc_3_31_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_3_31_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_3_31_wea : OUT STD_LOGIC;
    xt_rsc_3_31_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_3_31_lz : OUT STD_LOGIC;
    xt_rsc_4_0_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_4_0_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_0_wea : OUT STD_LOGIC;
    xt_rsc_4_0_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_4_0_lz : OUT STD_LOGIC;
    xt_rsc_4_1_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_4_1_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_1_wea : OUT STD_LOGIC;
    xt_rsc_4_1_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_4_1_lz : OUT STD_LOGIC;
    xt_rsc_4_2_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_4_2_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_2_wea : OUT STD_LOGIC;
    xt_rsc_4_2_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_4_2_lz : OUT STD_LOGIC;
    xt_rsc_4_3_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_4_3_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_3_wea : OUT STD_LOGIC;
    xt_rsc_4_3_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_4_3_lz : OUT STD_LOGIC;
    xt_rsc_4_4_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_4_4_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_4_wea : OUT STD_LOGIC;
    xt_rsc_4_4_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_4_4_lz : OUT STD_LOGIC;
    xt_rsc_4_5_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_4_5_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_5_wea : OUT STD_LOGIC;
    xt_rsc_4_5_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_4_5_lz : OUT STD_LOGIC;
    xt_rsc_4_6_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_4_6_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_6_wea : OUT STD_LOGIC;
    xt_rsc_4_6_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_4_6_lz : OUT STD_LOGIC;
    xt_rsc_4_7_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_4_7_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_7_wea : OUT STD_LOGIC;
    xt_rsc_4_7_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_4_7_lz : OUT STD_LOGIC;
    xt_rsc_4_8_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_4_8_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_8_wea : OUT STD_LOGIC;
    xt_rsc_4_8_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_4_8_lz : OUT STD_LOGIC;
    xt_rsc_4_9_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_4_9_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_9_wea : OUT STD_LOGIC;
    xt_rsc_4_9_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_4_9_lz : OUT STD_LOGIC;
    xt_rsc_4_10_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_4_10_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_10_wea : OUT STD_LOGIC;
    xt_rsc_4_10_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_4_10_lz : OUT STD_LOGIC;
    xt_rsc_4_11_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_4_11_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_11_wea : OUT STD_LOGIC;
    xt_rsc_4_11_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_4_11_lz : OUT STD_LOGIC;
    xt_rsc_4_12_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_4_12_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_12_wea : OUT STD_LOGIC;
    xt_rsc_4_12_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_4_12_lz : OUT STD_LOGIC;
    xt_rsc_4_13_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_4_13_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_13_wea : OUT STD_LOGIC;
    xt_rsc_4_13_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_4_13_lz : OUT STD_LOGIC;
    xt_rsc_4_14_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_4_14_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_14_wea : OUT STD_LOGIC;
    xt_rsc_4_14_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_4_14_lz : OUT STD_LOGIC;
    xt_rsc_4_15_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_4_15_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_15_wea : OUT STD_LOGIC;
    xt_rsc_4_15_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_4_15_lz : OUT STD_LOGIC;
    xt_rsc_4_16_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_4_16_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_16_wea : OUT STD_LOGIC;
    xt_rsc_4_16_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_4_16_lz : OUT STD_LOGIC;
    xt_rsc_4_17_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_4_17_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_17_wea : OUT STD_LOGIC;
    xt_rsc_4_17_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_4_17_lz : OUT STD_LOGIC;
    xt_rsc_4_18_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_4_18_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_18_wea : OUT STD_LOGIC;
    xt_rsc_4_18_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_4_18_lz : OUT STD_LOGIC;
    xt_rsc_4_19_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_4_19_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_19_wea : OUT STD_LOGIC;
    xt_rsc_4_19_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_4_19_lz : OUT STD_LOGIC;
    xt_rsc_4_20_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_4_20_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_20_wea : OUT STD_LOGIC;
    xt_rsc_4_20_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_4_20_lz : OUT STD_LOGIC;
    xt_rsc_4_21_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_4_21_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_21_wea : OUT STD_LOGIC;
    xt_rsc_4_21_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_4_21_lz : OUT STD_LOGIC;
    xt_rsc_4_22_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_4_22_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_22_wea : OUT STD_LOGIC;
    xt_rsc_4_22_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_4_22_lz : OUT STD_LOGIC;
    xt_rsc_4_23_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_4_23_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_23_wea : OUT STD_LOGIC;
    xt_rsc_4_23_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_4_23_lz : OUT STD_LOGIC;
    xt_rsc_4_24_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_4_24_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_24_wea : OUT STD_LOGIC;
    xt_rsc_4_24_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_4_24_lz : OUT STD_LOGIC;
    xt_rsc_4_25_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_4_25_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_25_wea : OUT STD_LOGIC;
    xt_rsc_4_25_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_4_25_lz : OUT STD_LOGIC;
    xt_rsc_4_26_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_4_26_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_26_wea : OUT STD_LOGIC;
    xt_rsc_4_26_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_4_26_lz : OUT STD_LOGIC;
    xt_rsc_4_27_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_4_27_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_27_wea : OUT STD_LOGIC;
    xt_rsc_4_27_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_4_27_lz : OUT STD_LOGIC;
    xt_rsc_4_28_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_4_28_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_28_wea : OUT STD_LOGIC;
    xt_rsc_4_28_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_4_28_lz : OUT STD_LOGIC;
    xt_rsc_4_29_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_4_29_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_29_wea : OUT STD_LOGIC;
    xt_rsc_4_29_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_4_29_lz : OUT STD_LOGIC;
    xt_rsc_4_30_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_4_30_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_30_wea : OUT STD_LOGIC;
    xt_rsc_4_30_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_4_30_lz : OUT STD_LOGIC;
    xt_rsc_4_31_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_4_31_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_4_31_wea : OUT STD_LOGIC;
    xt_rsc_4_31_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_4_31_lz : OUT STD_LOGIC;
    xt_rsc_5_0_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_5_0_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_5_0_wea : OUT STD_LOGIC;
    xt_rsc_5_0_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_5_0_lz : OUT STD_LOGIC;
    xt_rsc_5_1_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_5_1_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_5_1_wea : OUT STD_LOGIC;
    xt_rsc_5_1_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_5_1_lz : OUT STD_LOGIC;
    xt_rsc_5_2_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_5_2_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_5_2_wea : OUT STD_LOGIC;
    xt_rsc_5_2_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_5_2_lz : OUT STD_LOGIC;
    xt_rsc_5_3_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_5_3_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_5_3_wea : OUT STD_LOGIC;
    xt_rsc_5_3_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_5_3_lz : OUT STD_LOGIC;
    xt_rsc_5_4_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_5_4_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_5_4_wea : OUT STD_LOGIC;
    xt_rsc_5_4_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_5_4_lz : OUT STD_LOGIC;
    xt_rsc_5_5_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_5_5_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_5_5_wea : OUT STD_LOGIC;
    xt_rsc_5_5_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_5_5_lz : OUT STD_LOGIC;
    xt_rsc_5_6_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_5_6_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_5_6_wea : OUT STD_LOGIC;
    xt_rsc_5_6_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_5_6_lz : OUT STD_LOGIC;
    xt_rsc_5_7_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_5_7_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_5_7_wea : OUT STD_LOGIC;
    xt_rsc_5_7_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_5_7_lz : OUT STD_LOGIC;
    xt_rsc_5_8_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_5_8_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_5_8_wea : OUT STD_LOGIC;
    xt_rsc_5_8_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_5_8_lz : OUT STD_LOGIC;
    xt_rsc_5_9_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_5_9_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_5_9_wea : OUT STD_LOGIC;
    xt_rsc_5_9_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_5_9_lz : OUT STD_LOGIC;
    xt_rsc_5_10_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_5_10_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_5_10_wea : OUT STD_LOGIC;
    xt_rsc_5_10_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_5_10_lz : OUT STD_LOGIC;
    xt_rsc_5_11_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_5_11_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_5_11_wea : OUT STD_LOGIC;
    xt_rsc_5_11_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_5_11_lz : OUT STD_LOGIC;
    xt_rsc_5_12_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_5_12_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_5_12_wea : OUT STD_LOGIC;
    xt_rsc_5_12_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_5_12_lz : OUT STD_LOGIC;
    xt_rsc_5_13_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_5_13_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_5_13_wea : OUT STD_LOGIC;
    xt_rsc_5_13_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_5_13_lz : OUT STD_LOGIC;
    xt_rsc_5_14_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_5_14_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_5_14_wea : OUT STD_LOGIC;
    xt_rsc_5_14_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_5_14_lz : OUT STD_LOGIC;
    xt_rsc_5_15_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_5_15_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_5_15_wea : OUT STD_LOGIC;
    xt_rsc_5_15_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_5_15_lz : OUT STD_LOGIC;
    xt_rsc_5_16_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_5_16_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_5_16_wea : OUT STD_LOGIC;
    xt_rsc_5_16_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_5_16_lz : OUT STD_LOGIC;
    xt_rsc_5_17_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_5_17_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_5_17_wea : OUT STD_LOGIC;
    xt_rsc_5_17_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_5_17_lz : OUT STD_LOGIC;
    xt_rsc_5_18_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_5_18_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_5_18_wea : OUT STD_LOGIC;
    xt_rsc_5_18_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_5_18_lz : OUT STD_LOGIC;
    xt_rsc_5_19_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_5_19_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_5_19_wea : OUT STD_LOGIC;
    xt_rsc_5_19_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_5_19_lz : OUT STD_LOGIC;
    xt_rsc_5_20_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_5_20_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_5_20_wea : OUT STD_LOGIC;
    xt_rsc_5_20_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_5_20_lz : OUT STD_LOGIC;
    xt_rsc_5_21_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_5_21_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_5_21_wea : OUT STD_LOGIC;
    xt_rsc_5_21_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_5_21_lz : OUT STD_LOGIC;
    xt_rsc_5_22_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_5_22_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_5_22_wea : OUT STD_LOGIC;
    xt_rsc_5_22_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_5_22_lz : OUT STD_LOGIC;
    xt_rsc_5_23_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_5_23_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_5_23_wea : OUT STD_LOGIC;
    xt_rsc_5_23_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_5_23_lz : OUT STD_LOGIC;
    xt_rsc_5_24_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_5_24_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_5_24_wea : OUT STD_LOGIC;
    xt_rsc_5_24_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_5_24_lz : OUT STD_LOGIC;
    xt_rsc_5_25_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_5_25_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_5_25_wea : OUT STD_LOGIC;
    xt_rsc_5_25_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_5_25_lz : OUT STD_LOGIC;
    xt_rsc_5_26_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_5_26_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_5_26_wea : OUT STD_LOGIC;
    xt_rsc_5_26_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_5_26_lz : OUT STD_LOGIC;
    xt_rsc_5_27_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_5_27_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_5_27_wea : OUT STD_LOGIC;
    xt_rsc_5_27_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_5_27_lz : OUT STD_LOGIC;
    xt_rsc_5_28_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_5_28_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_5_28_wea : OUT STD_LOGIC;
    xt_rsc_5_28_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_5_28_lz : OUT STD_LOGIC;
    xt_rsc_5_29_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_5_29_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_5_29_wea : OUT STD_LOGIC;
    xt_rsc_5_29_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_5_29_lz : OUT STD_LOGIC;
    xt_rsc_5_30_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_5_30_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_5_30_wea : OUT STD_LOGIC;
    xt_rsc_5_30_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_5_30_lz : OUT STD_LOGIC;
    xt_rsc_5_31_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_5_31_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_5_31_wea : OUT STD_LOGIC;
    xt_rsc_5_31_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_5_31_lz : OUT STD_LOGIC;
    xt_rsc_6_0_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_6_0_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_6_0_wea : OUT STD_LOGIC;
    xt_rsc_6_0_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_6_0_lz : OUT STD_LOGIC;
    xt_rsc_6_1_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_6_1_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_6_1_wea : OUT STD_LOGIC;
    xt_rsc_6_1_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_6_1_lz : OUT STD_LOGIC;
    xt_rsc_6_2_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_6_2_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_6_2_wea : OUT STD_LOGIC;
    xt_rsc_6_2_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_6_2_lz : OUT STD_LOGIC;
    xt_rsc_6_3_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_6_3_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_6_3_wea : OUT STD_LOGIC;
    xt_rsc_6_3_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_6_3_lz : OUT STD_LOGIC;
    xt_rsc_6_4_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_6_4_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_6_4_wea : OUT STD_LOGIC;
    xt_rsc_6_4_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_6_4_lz : OUT STD_LOGIC;
    xt_rsc_6_5_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_6_5_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_6_5_wea : OUT STD_LOGIC;
    xt_rsc_6_5_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_6_5_lz : OUT STD_LOGIC;
    xt_rsc_6_6_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_6_6_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_6_6_wea : OUT STD_LOGIC;
    xt_rsc_6_6_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_6_6_lz : OUT STD_LOGIC;
    xt_rsc_6_7_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_6_7_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_6_7_wea : OUT STD_LOGIC;
    xt_rsc_6_7_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_6_7_lz : OUT STD_LOGIC;
    xt_rsc_6_8_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_6_8_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_6_8_wea : OUT STD_LOGIC;
    xt_rsc_6_8_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_6_8_lz : OUT STD_LOGIC;
    xt_rsc_6_9_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_6_9_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_6_9_wea : OUT STD_LOGIC;
    xt_rsc_6_9_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_6_9_lz : OUT STD_LOGIC;
    xt_rsc_6_10_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_6_10_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_6_10_wea : OUT STD_LOGIC;
    xt_rsc_6_10_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_6_10_lz : OUT STD_LOGIC;
    xt_rsc_6_11_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_6_11_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_6_11_wea : OUT STD_LOGIC;
    xt_rsc_6_11_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_6_11_lz : OUT STD_LOGIC;
    xt_rsc_6_12_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_6_12_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_6_12_wea : OUT STD_LOGIC;
    xt_rsc_6_12_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_6_12_lz : OUT STD_LOGIC;
    xt_rsc_6_13_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_6_13_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_6_13_wea : OUT STD_LOGIC;
    xt_rsc_6_13_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_6_13_lz : OUT STD_LOGIC;
    xt_rsc_6_14_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_6_14_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_6_14_wea : OUT STD_LOGIC;
    xt_rsc_6_14_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_6_14_lz : OUT STD_LOGIC;
    xt_rsc_6_15_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_6_15_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_6_15_wea : OUT STD_LOGIC;
    xt_rsc_6_15_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_6_15_lz : OUT STD_LOGIC;
    xt_rsc_6_16_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_6_16_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_6_16_wea : OUT STD_LOGIC;
    xt_rsc_6_16_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_6_16_lz : OUT STD_LOGIC;
    xt_rsc_6_17_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_6_17_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_6_17_wea : OUT STD_LOGIC;
    xt_rsc_6_17_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_6_17_lz : OUT STD_LOGIC;
    xt_rsc_6_18_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_6_18_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_6_18_wea : OUT STD_LOGIC;
    xt_rsc_6_18_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_6_18_lz : OUT STD_LOGIC;
    xt_rsc_6_19_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_6_19_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_6_19_wea : OUT STD_LOGIC;
    xt_rsc_6_19_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_6_19_lz : OUT STD_LOGIC;
    xt_rsc_6_20_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_6_20_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_6_20_wea : OUT STD_LOGIC;
    xt_rsc_6_20_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_6_20_lz : OUT STD_LOGIC;
    xt_rsc_6_21_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_6_21_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_6_21_wea : OUT STD_LOGIC;
    xt_rsc_6_21_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_6_21_lz : OUT STD_LOGIC;
    xt_rsc_6_22_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_6_22_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_6_22_wea : OUT STD_LOGIC;
    xt_rsc_6_22_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_6_22_lz : OUT STD_LOGIC;
    xt_rsc_6_23_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_6_23_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_6_23_wea : OUT STD_LOGIC;
    xt_rsc_6_23_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_6_23_lz : OUT STD_LOGIC;
    xt_rsc_6_24_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_6_24_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_6_24_wea : OUT STD_LOGIC;
    xt_rsc_6_24_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_6_24_lz : OUT STD_LOGIC;
    xt_rsc_6_25_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_6_25_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_6_25_wea : OUT STD_LOGIC;
    xt_rsc_6_25_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_6_25_lz : OUT STD_LOGIC;
    xt_rsc_6_26_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_6_26_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_6_26_wea : OUT STD_LOGIC;
    xt_rsc_6_26_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_6_26_lz : OUT STD_LOGIC;
    xt_rsc_6_27_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_6_27_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_6_27_wea : OUT STD_LOGIC;
    xt_rsc_6_27_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_6_27_lz : OUT STD_LOGIC;
    xt_rsc_6_28_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_6_28_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_6_28_wea : OUT STD_LOGIC;
    xt_rsc_6_28_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_6_28_lz : OUT STD_LOGIC;
    xt_rsc_6_29_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_6_29_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_6_29_wea : OUT STD_LOGIC;
    xt_rsc_6_29_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_6_29_lz : OUT STD_LOGIC;
    xt_rsc_6_30_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_6_30_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_6_30_wea : OUT STD_LOGIC;
    xt_rsc_6_30_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_6_30_lz : OUT STD_LOGIC;
    xt_rsc_6_31_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_6_31_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_6_31_wea : OUT STD_LOGIC;
    xt_rsc_6_31_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_6_31_lz : OUT STD_LOGIC;
    xt_rsc_7_0_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_7_0_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_7_0_wea : OUT STD_LOGIC;
    xt_rsc_7_0_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_7_0_lz : OUT STD_LOGIC;
    xt_rsc_7_1_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_7_1_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_7_1_wea : OUT STD_LOGIC;
    xt_rsc_7_1_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_7_1_lz : OUT STD_LOGIC;
    xt_rsc_7_2_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_7_2_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_7_2_wea : OUT STD_LOGIC;
    xt_rsc_7_2_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_7_2_lz : OUT STD_LOGIC;
    xt_rsc_7_3_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_7_3_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_7_3_wea : OUT STD_LOGIC;
    xt_rsc_7_3_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_7_3_lz : OUT STD_LOGIC;
    xt_rsc_7_4_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_7_4_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_7_4_wea : OUT STD_LOGIC;
    xt_rsc_7_4_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_7_4_lz : OUT STD_LOGIC;
    xt_rsc_7_5_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_7_5_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_7_5_wea : OUT STD_LOGIC;
    xt_rsc_7_5_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_7_5_lz : OUT STD_LOGIC;
    xt_rsc_7_6_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_7_6_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_7_6_wea : OUT STD_LOGIC;
    xt_rsc_7_6_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_7_6_lz : OUT STD_LOGIC;
    xt_rsc_7_7_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_7_7_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_7_7_wea : OUT STD_LOGIC;
    xt_rsc_7_7_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_7_7_lz : OUT STD_LOGIC;
    xt_rsc_7_8_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_7_8_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_7_8_wea : OUT STD_LOGIC;
    xt_rsc_7_8_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_7_8_lz : OUT STD_LOGIC;
    xt_rsc_7_9_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_7_9_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_7_9_wea : OUT STD_LOGIC;
    xt_rsc_7_9_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_7_9_lz : OUT STD_LOGIC;
    xt_rsc_7_10_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_7_10_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_7_10_wea : OUT STD_LOGIC;
    xt_rsc_7_10_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_7_10_lz : OUT STD_LOGIC;
    xt_rsc_7_11_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_7_11_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_7_11_wea : OUT STD_LOGIC;
    xt_rsc_7_11_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_7_11_lz : OUT STD_LOGIC;
    xt_rsc_7_12_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_7_12_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_7_12_wea : OUT STD_LOGIC;
    xt_rsc_7_12_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_7_12_lz : OUT STD_LOGIC;
    xt_rsc_7_13_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_7_13_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_7_13_wea : OUT STD_LOGIC;
    xt_rsc_7_13_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_7_13_lz : OUT STD_LOGIC;
    xt_rsc_7_14_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_7_14_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_7_14_wea : OUT STD_LOGIC;
    xt_rsc_7_14_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_7_14_lz : OUT STD_LOGIC;
    xt_rsc_7_15_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_7_15_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_7_15_wea : OUT STD_LOGIC;
    xt_rsc_7_15_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_7_15_lz : OUT STD_LOGIC;
    xt_rsc_7_16_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_7_16_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_7_16_wea : OUT STD_LOGIC;
    xt_rsc_7_16_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_7_16_lz : OUT STD_LOGIC;
    xt_rsc_7_17_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_7_17_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_7_17_wea : OUT STD_LOGIC;
    xt_rsc_7_17_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_7_17_lz : OUT STD_LOGIC;
    xt_rsc_7_18_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_7_18_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_7_18_wea : OUT STD_LOGIC;
    xt_rsc_7_18_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_7_18_lz : OUT STD_LOGIC;
    xt_rsc_7_19_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_7_19_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_7_19_wea : OUT STD_LOGIC;
    xt_rsc_7_19_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_7_19_lz : OUT STD_LOGIC;
    xt_rsc_7_20_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_7_20_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_7_20_wea : OUT STD_LOGIC;
    xt_rsc_7_20_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_7_20_lz : OUT STD_LOGIC;
    xt_rsc_7_21_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_7_21_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_7_21_wea : OUT STD_LOGIC;
    xt_rsc_7_21_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_7_21_lz : OUT STD_LOGIC;
    xt_rsc_7_22_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_7_22_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_7_22_wea : OUT STD_LOGIC;
    xt_rsc_7_22_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_7_22_lz : OUT STD_LOGIC;
    xt_rsc_7_23_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_7_23_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_7_23_wea : OUT STD_LOGIC;
    xt_rsc_7_23_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_7_23_lz : OUT STD_LOGIC;
    xt_rsc_7_24_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_7_24_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_7_24_wea : OUT STD_LOGIC;
    xt_rsc_7_24_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_7_24_lz : OUT STD_LOGIC;
    xt_rsc_7_25_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_7_25_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_7_25_wea : OUT STD_LOGIC;
    xt_rsc_7_25_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_7_25_lz : OUT STD_LOGIC;
    xt_rsc_7_26_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_7_26_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_7_26_wea : OUT STD_LOGIC;
    xt_rsc_7_26_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_7_26_lz : OUT STD_LOGIC;
    xt_rsc_7_27_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_7_27_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_7_27_wea : OUT STD_LOGIC;
    xt_rsc_7_27_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_7_27_lz : OUT STD_LOGIC;
    xt_rsc_7_28_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_7_28_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_7_28_wea : OUT STD_LOGIC;
    xt_rsc_7_28_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_7_28_lz : OUT STD_LOGIC;
    xt_rsc_7_29_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_7_29_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_7_29_wea : OUT STD_LOGIC;
    xt_rsc_7_29_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_7_29_lz : OUT STD_LOGIC;
    xt_rsc_7_30_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_7_30_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_7_30_wea : OUT STD_LOGIC;
    xt_rsc_7_30_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_7_30_lz : OUT STD_LOGIC;
    xt_rsc_7_31_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_7_31_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_7_31_wea : OUT STD_LOGIC;
    xt_rsc_7_31_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_7_31_lz : OUT STD_LOGIC;
    p_rsc_dat : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    p_rsc_triosy_lz : OUT STD_LOGIC;
    r_rsc_dat : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    r_rsc_triosy_lz : OUT STD_LOGIC;
    twiddle_rsc_0_0_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_0_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_0_wea : OUT STD_LOGIC;
    twiddle_rsc_0_0_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_0_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_0_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_0_web : OUT STD_LOGIC;
    twiddle_rsc_0_0_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_triosy_0_0_lz : OUT STD_LOGIC;
    twiddle_rsc_0_1_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_1_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_1_wea : OUT STD_LOGIC;
    twiddle_rsc_0_1_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_1_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_1_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_1_web : OUT STD_LOGIC;
    twiddle_rsc_0_1_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_triosy_0_1_lz : OUT STD_LOGIC;
    twiddle_rsc_0_2_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_2_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_2_wea : OUT STD_LOGIC;
    twiddle_rsc_0_2_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_2_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_2_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_2_web : OUT STD_LOGIC;
    twiddle_rsc_0_2_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_triosy_0_2_lz : OUT STD_LOGIC;
    twiddle_rsc_0_3_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_3_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_3_wea : OUT STD_LOGIC;
    twiddle_rsc_0_3_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_3_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_3_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_3_web : OUT STD_LOGIC;
    twiddle_rsc_0_3_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_triosy_0_3_lz : OUT STD_LOGIC;
    twiddle_rsc_0_4_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_4_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_4_wea : OUT STD_LOGIC;
    twiddle_rsc_0_4_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_4_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_4_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_4_web : OUT STD_LOGIC;
    twiddle_rsc_0_4_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_triosy_0_4_lz : OUT STD_LOGIC;
    twiddle_rsc_0_5_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_5_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_5_wea : OUT STD_LOGIC;
    twiddle_rsc_0_5_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_5_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_5_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_5_web : OUT STD_LOGIC;
    twiddle_rsc_0_5_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_triosy_0_5_lz : OUT STD_LOGIC;
    twiddle_rsc_0_6_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_6_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_6_wea : OUT STD_LOGIC;
    twiddle_rsc_0_6_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_6_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_6_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_6_web : OUT STD_LOGIC;
    twiddle_rsc_0_6_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_triosy_0_6_lz : OUT STD_LOGIC;
    twiddle_rsc_0_7_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_7_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_7_wea : OUT STD_LOGIC;
    twiddle_rsc_0_7_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_7_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_7_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_7_web : OUT STD_LOGIC;
    twiddle_rsc_0_7_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_triosy_0_7_lz : OUT STD_LOGIC;
    twiddle_rsc_0_8_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_8_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_8_wea : OUT STD_LOGIC;
    twiddle_rsc_0_8_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_8_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_8_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_8_web : OUT STD_LOGIC;
    twiddle_rsc_0_8_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_triosy_0_8_lz : OUT STD_LOGIC;
    twiddle_rsc_0_9_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_9_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_9_wea : OUT STD_LOGIC;
    twiddle_rsc_0_9_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_9_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_9_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_9_web : OUT STD_LOGIC;
    twiddle_rsc_0_9_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_triosy_0_9_lz : OUT STD_LOGIC;
    twiddle_rsc_0_10_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_10_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_10_wea : OUT STD_LOGIC;
    twiddle_rsc_0_10_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_10_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_10_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_10_web : OUT STD_LOGIC;
    twiddle_rsc_0_10_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_triosy_0_10_lz : OUT STD_LOGIC;
    twiddle_rsc_0_11_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_11_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_11_wea : OUT STD_LOGIC;
    twiddle_rsc_0_11_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_11_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_11_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_11_web : OUT STD_LOGIC;
    twiddle_rsc_0_11_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_triosy_0_11_lz : OUT STD_LOGIC;
    twiddle_rsc_0_12_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_12_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_12_wea : OUT STD_LOGIC;
    twiddle_rsc_0_12_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_12_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_12_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_12_web : OUT STD_LOGIC;
    twiddle_rsc_0_12_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_triosy_0_12_lz : OUT STD_LOGIC;
    twiddle_rsc_0_13_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_13_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_13_wea : OUT STD_LOGIC;
    twiddle_rsc_0_13_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_13_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_13_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_13_web : OUT STD_LOGIC;
    twiddle_rsc_0_13_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_triosy_0_13_lz : OUT STD_LOGIC;
    twiddle_rsc_0_14_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_14_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_14_wea : OUT STD_LOGIC;
    twiddle_rsc_0_14_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_14_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_14_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_14_web : OUT STD_LOGIC;
    twiddle_rsc_0_14_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_triosy_0_14_lz : OUT STD_LOGIC;
    twiddle_rsc_0_15_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_15_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_15_wea : OUT STD_LOGIC;
    twiddle_rsc_0_15_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_15_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_15_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_15_web : OUT STD_LOGIC;
    twiddle_rsc_0_15_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_triosy_0_15_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_0_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_0_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_0_wea : OUT STD_LOGIC;
    twiddle_h_rsc_0_0_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_0_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_0_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_0_web : OUT STD_LOGIC;
    twiddle_h_rsc_0_0_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_triosy_0_0_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_1_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_1_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_1_wea : OUT STD_LOGIC;
    twiddle_h_rsc_0_1_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_1_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_1_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_1_web : OUT STD_LOGIC;
    twiddle_h_rsc_0_1_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_triosy_0_1_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_2_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_2_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_2_wea : OUT STD_LOGIC;
    twiddle_h_rsc_0_2_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_2_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_2_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_2_web : OUT STD_LOGIC;
    twiddle_h_rsc_0_2_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_triosy_0_2_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_3_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_3_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_3_wea : OUT STD_LOGIC;
    twiddle_h_rsc_0_3_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_3_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_3_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_3_web : OUT STD_LOGIC;
    twiddle_h_rsc_0_3_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_triosy_0_3_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_4_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_4_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_4_wea : OUT STD_LOGIC;
    twiddle_h_rsc_0_4_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_4_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_4_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_4_web : OUT STD_LOGIC;
    twiddle_h_rsc_0_4_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_triosy_0_4_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_5_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_5_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_5_wea : OUT STD_LOGIC;
    twiddle_h_rsc_0_5_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_5_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_5_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_5_web : OUT STD_LOGIC;
    twiddle_h_rsc_0_5_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_triosy_0_5_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_6_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_6_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_6_wea : OUT STD_LOGIC;
    twiddle_h_rsc_0_6_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_6_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_6_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_6_web : OUT STD_LOGIC;
    twiddle_h_rsc_0_6_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_triosy_0_6_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_7_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_7_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_7_wea : OUT STD_LOGIC;
    twiddle_h_rsc_0_7_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_7_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_7_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_7_web : OUT STD_LOGIC;
    twiddle_h_rsc_0_7_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_triosy_0_7_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_8_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_8_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_8_wea : OUT STD_LOGIC;
    twiddle_h_rsc_0_8_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_8_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_8_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_8_web : OUT STD_LOGIC;
    twiddle_h_rsc_0_8_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_triosy_0_8_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_9_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_9_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_9_wea : OUT STD_LOGIC;
    twiddle_h_rsc_0_9_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_9_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_9_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_9_web : OUT STD_LOGIC;
    twiddle_h_rsc_0_9_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_triosy_0_9_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_10_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_10_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_10_wea : OUT STD_LOGIC;
    twiddle_h_rsc_0_10_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_10_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_10_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_10_web : OUT STD_LOGIC;
    twiddle_h_rsc_0_10_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_triosy_0_10_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_11_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_11_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_11_wea : OUT STD_LOGIC;
    twiddle_h_rsc_0_11_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_11_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_11_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_11_web : OUT STD_LOGIC;
    twiddle_h_rsc_0_11_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_triosy_0_11_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_12_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_12_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_12_wea : OUT STD_LOGIC;
    twiddle_h_rsc_0_12_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_12_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_12_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_12_web : OUT STD_LOGIC;
    twiddle_h_rsc_0_12_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_triosy_0_12_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_13_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_13_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_13_wea : OUT STD_LOGIC;
    twiddle_h_rsc_0_13_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_13_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_13_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_13_web : OUT STD_LOGIC;
    twiddle_h_rsc_0_13_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_triosy_0_13_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_14_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_14_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_14_wea : OUT STD_LOGIC;
    twiddle_h_rsc_0_14_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_14_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_14_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_14_web : OUT STD_LOGIC;
    twiddle_h_rsc_0_14_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_triosy_0_14_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_15_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_15_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_15_wea : OUT STD_LOGIC;
    twiddle_h_rsc_0_15_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_15_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_15_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_15_web : OUT STD_LOGIC;
    twiddle_h_rsc_0_15_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_triosy_0_15_lz : OUT STD_LOGIC
  );
END peaseNTT;

ARCHITECTURE v14 OF peaseNTT IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';

  -- Interconnect Declarations
  SIGNAL yt_rsc_0_0_i_clkr_en_d : STD_LOGIC;
  SIGNAL yt_rsc_0_0_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_1_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_2_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_3_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_4_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_5_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_6_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_7_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_8_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_9_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_10_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_11_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_12_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_13_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_14_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_15_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_16_i_clkr_en_d : STD_LOGIC;
  SIGNAL yt_rsc_0_16_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_17_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_18_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_19_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_20_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_21_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_22_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_23_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_24_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_25_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_26_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_27_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_28_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_29_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_30_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_31_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_0_i_clkr_en_d : STD_LOGIC;
  SIGNAL yt_rsc_1_0_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_1_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_2_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_3_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_4_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_5_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_6_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_7_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_8_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_9_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_10_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_11_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_12_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_13_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_14_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_15_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_16_i_clkr_en_d : STD_LOGIC;
  SIGNAL yt_rsc_1_16_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_17_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_18_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_19_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_20_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_21_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_22_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_23_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_24_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_25_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_26_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_27_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_28_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_29_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_30_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_31_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_0_i_clkr_en_d : STD_LOGIC;
  SIGNAL yt_rsc_2_0_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_1_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_2_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_3_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_4_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_5_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_6_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_7_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_8_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_9_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_10_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_11_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_12_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_13_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_14_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_15_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_16_i_clkr_en_d : STD_LOGIC;
  SIGNAL yt_rsc_2_16_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_17_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_18_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_19_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_20_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_21_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_22_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_23_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_24_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_25_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_26_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_27_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_28_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_29_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_30_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_31_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_0_i_clkr_en_d : STD_LOGIC;
  SIGNAL yt_rsc_3_0_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_1_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_2_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_3_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_4_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_5_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_6_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_7_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_8_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_9_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_10_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_11_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_12_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_13_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_14_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_15_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_16_i_clkr_en_d : STD_LOGIC;
  SIGNAL yt_rsc_3_16_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_17_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_18_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_19_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_20_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_21_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_22_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_23_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_24_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_25_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_26_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_27_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_28_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_29_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_30_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_31_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_0_i_clkr_en_d : STD_LOGIC;
  SIGNAL yt_rsc_4_0_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_1_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_2_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_3_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_4_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_5_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_6_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_7_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_8_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_9_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_10_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_11_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_12_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_13_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_14_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_15_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_16_i_clkr_en_d : STD_LOGIC;
  SIGNAL yt_rsc_4_16_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_17_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_18_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_19_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_20_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_21_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_22_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_23_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_24_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_25_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_26_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_27_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_28_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_29_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_30_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_31_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_0_i_clkr_en_d : STD_LOGIC;
  SIGNAL yt_rsc_5_0_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_1_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_2_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_3_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_4_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_5_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_6_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_7_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_8_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_9_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_10_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_11_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_12_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_13_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_14_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_15_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_16_i_clkr_en_d : STD_LOGIC;
  SIGNAL yt_rsc_5_16_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_17_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_18_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_19_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_20_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_21_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_22_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_23_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_24_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_25_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_26_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_27_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_28_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_29_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_30_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_31_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_0_i_clkr_en_d : STD_LOGIC;
  SIGNAL yt_rsc_6_0_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_1_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_2_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_3_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_4_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_5_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_6_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_7_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_8_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_9_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_10_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_11_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_12_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_13_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_14_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_15_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_16_i_clkr_en_d : STD_LOGIC;
  SIGNAL yt_rsc_6_16_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_17_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_18_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_19_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_20_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_21_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_22_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_23_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_24_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_25_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_26_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_27_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_28_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_29_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_30_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_31_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_0_i_clkr_en_d : STD_LOGIC;
  SIGNAL yt_rsc_7_0_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_1_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_2_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_3_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_4_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_5_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_6_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_7_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_8_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_9_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_10_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_11_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_12_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_13_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_14_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_15_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_16_i_clkr_en_d : STD_LOGIC;
  SIGNAL yt_rsc_7_16_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_17_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_18_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_19_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_20_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_21_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_22_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_23_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_24_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_25_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_26_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_27_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_28_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_29_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_30_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_31_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_0_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_1_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_2_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_3_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_4_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_5_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_6_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_7_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_8_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_9_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_10_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_11_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_12_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_13_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_14_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_15_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_16_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_17_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_18_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_19_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_20_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_21_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_22_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_23_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_24_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_25_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_26_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_27_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_28_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_29_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_30_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_31_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_0_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_1_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_2_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_3_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_4_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_5_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_6_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_7_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_8_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_9_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_10_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_11_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_12_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_13_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_14_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_15_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_16_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_17_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_18_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_19_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_20_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_21_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_22_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_23_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_24_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_25_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_26_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_27_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_28_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_29_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_30_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_31_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_0_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_1_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_2_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_3_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_4_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_5_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_6_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_7_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_8_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_9_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_10_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_11_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_12_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_13_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_14_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_15_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_16_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_17_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_18_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_19_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_20_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_21_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_22_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_23_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_24_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_25_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_26_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_27_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_28_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_29_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_30_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_31_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_0_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_1_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_2_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_3_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_4_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_5_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_6_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_7_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_8_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_9_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_10_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_11_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_12_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_13_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_14_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_15_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_16_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_17_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_18_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_19_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_20_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_21_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_22_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_23_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_24_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_25_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_26_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_27_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_28_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_29_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_30_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_31_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_0_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_1_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_2_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_3_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_4_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_5_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_6_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_7_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_8_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_9_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_10_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_11_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_12_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_13_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_14_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_15_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_16_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_17_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_18_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_19_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_20_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_21_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_22_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_23_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_24_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_25_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_26_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_27_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_28_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_29_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_30_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_31_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_0_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_1_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_2_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_3_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_4_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_5_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_6_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_7_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_8_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_9_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_10_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_11_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_12_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_13_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_14_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_15_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_16_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_17_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_18_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_19_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_20_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_21_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_22_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_23_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_24_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_25_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_26_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_27_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_28_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_29_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_30_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_31_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_0_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_1_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_2_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_3_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_4_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_5_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_6_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_7_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_8_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_9_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_10_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_11_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_12_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_13_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_14_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_15_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_16_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_17_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_18_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_19_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_20_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_21_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_22_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_23_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_24_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_25_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_26_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_27_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_28_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_29_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_30_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_31_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_0_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_1_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_2_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_3_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_4_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_5_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_6_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_7_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_8_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_9_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_10_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_11_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_12_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_13_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_14_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_15_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_16_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_17_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_18_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_19_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_20_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_21_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_22_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_23_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_24_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_25_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_26_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_27_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_28_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_29_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_30_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_31_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1
      DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1
      DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1
      DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1
      DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1
      DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1
      DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1
      DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1
      DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1
      DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1
      DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1
      DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1
      DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1
      DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1
      DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1
      DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1
      DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_8_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_8_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_9_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_9_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_10_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_10_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_11_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_11_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_12_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_12_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_13_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_13_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_14_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_14_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_15_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_15_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL yt_rsc_0_0_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_0_0_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_0_0_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_0_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_0_we : STD_LOGIC;
  SIGNAL yt_rsc_0_0_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_0_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_1_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_0_1_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_0_1_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_1_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_1_we : STD_LOGIC;
  SIGNAL yt_rsc_0_1_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_1_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_2_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_0_2_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_0_2_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_2_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_2_we : STD_LOGIC;
  SIGNAL yt_rsc_0_2_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_2_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_3_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_0_3_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_0_3_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_3_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_3_we : STD_LOGIC;
  SIGNAL yt_rsc_0_3_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_3_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_4_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_0_4_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_0_4_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_4_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_4_we : STD_LOGIC;
  SIGNAL yt_rsc_0_4_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_4_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_5_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_0_5_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_0_5_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_5_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_5_we : STD_LOGIC;
  SIGNAL yt_rsc_0_5_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_5_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_6_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_0_6_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_0_6_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_6_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_6_we : STD_LOGIC;
  SIGNAL yt_rsc_0_6_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_6_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_7_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_0_7_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_0_7_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_7_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_7_we : STD_LOGIC;
  SIGNAL yt_rsc_0_7_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_7_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_8_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_0_8_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_0_8_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_8_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_8_we : STD_LOGIC;
  SIGNAL yt_rsc_0_8_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_8_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_9_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_0_9_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_0_9_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_9_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_9_we : STD_LOGIC;
  SIGNAL yt_rsc_0_9_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_9_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_10_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_0_10_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_0_10_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_10_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_10_we : STD_LOGIC;
  SIGNAL yt_rsc_0_10_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_10_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_11_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_0_11_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_0_11_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_11_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_11_we : STD_LOGIC;
  SIGNAL yt_rsc_0_11_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_11_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_12_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_0_12_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_0_12_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_12_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_12_we : STD_LOGIC;
  SIGNAL yt_rsc_0_12_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_12_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_13_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_0_13_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_0_13_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_13_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_13_we : STD_LOGIC;
  SIGNAL yt_rsc_0_13_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_13_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_14_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_0_14_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_0_14_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_14_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_14_we : STD_LOGIC;
  SIGNAL yt_rsc_0_14_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_14_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_15_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_0_15_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_0_15_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_15_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_15_we : STD_LOGIC;
  SIGNAL yt_rsc_0_15_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_15_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_16_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_0_16_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_0_16_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_16_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_16_we : STD_LOGIC;
  SIGNAL yt_rsc_0_16_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_16_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_17_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_0_17_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_0_17_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_17_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_17_we : STD_LOGIC;
  SIGNAL yt_rsc_0_17_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_17_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_18_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_0_18_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_0_18_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_18_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_18_we : STD_LOGIC;
  SIGNAL yt_rsc_0_18_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_18_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_19_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_0_19_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_0_19_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_19_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_19_we : STD_LOGIC;
  SIGNAL yt_rsc_0_19_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_19_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_20_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_0_20_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_0_20_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_20_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_20_we : STD_LOGIC;
  SIGNAL yt_rsc_0_20_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_20_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_21_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_0_21_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_0_21_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_21_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_21_we : STD_LOGIC;
  SIGNAL yt_rsc_0_21_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_21_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_22_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_0_22_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_0_22_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_22_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_22_we : STD_LOGIC;
  SIGNAL yt_rsc_0_22_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_22_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_23_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_0_23_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_0_23_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_23_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_23_we : STD_LOGIC;
  SIGNAL yt_rsc_0_23_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_23_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_24_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_0_24_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_0_24_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_24_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_24_we : STD_LOGIC;
  SIGNAL yt_rsc_0_24_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_24_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_25_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_0_25_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_0_25_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_25_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_25_we : STD_LOGIC;
  SIGNAL yt_rsc_0_25_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_25_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_26_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_0_26_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_0_26_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_26_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_26_we : STD_LOGIC;
  SIGNAL yt_rsc_0_26_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_26_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_27_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_0_27_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_0_27_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_27_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_27_we : STD_LOGIC;
  SIGNAL yt_rsc_0_27_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_27_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_28_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_0_28_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_0_28_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_28_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_28_we : STD_LOGIC;
  SIGNAL yt_rsc_0_28_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_28_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_29_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_0_29_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_0_29_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_29_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_29_we : STD_LOGIC;
  SIGNAL yt_rsc_0_29_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_29_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_30_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_0_30_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_0_30_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_30_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_30_we : STD_LOGIC;
  SIGNAL yt_rsc_0_30_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_30_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_31_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_0_31_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_0_31_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_31_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_31_we : STD_LOGIC;
  SIGNAL yt_rsc_0_31_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_31_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_0_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_1_0_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_1_0_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_0_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_0_we : STD_LOGIC;
  SIGNAL yt_rsc_1_0_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_0_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_1_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_1_1_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_1_1_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_1_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_1_we : STD_LOGIC;
  SIGNAL yt_rsc_1_1_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_1_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_2_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_1_2_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_1_2_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_2_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_2_we : STD_LOGIC;
  SIGNAL yt_rsc_1_2_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_2_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_3_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_1_3_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_1_3_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_3_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_3_we : STD_LOGIC;
  SIGNAL yt_rsc_1_3_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_3_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_4_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_1_4_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_1_4_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_4_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_4_we : STD_LOGIC;
  SIGNAL yt_rsc_1_4_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_4_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_5_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_1_5_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_1_5_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_5_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_5_we : STD_LOGIC;
  SIGNAL yt_rsc_1_5_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_5_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_6_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_1_6_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_1_6_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_6_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_6_we : STD_LOGIC;
  SIGNAL yt_rsc_1_6_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_6_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_7_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_1_7_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_1_7_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_7_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_7_we : STD_LOGIC;
  SIGNAL yt_rsc_1_7_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_7_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_8_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_1_8_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_1_8_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_8_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_8_we : STD_LOGIC;
  SIGNAL yt_rsc_1_8_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_8_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_9_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_1_9_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_1_9_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_9_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_9_we : STD_LOGIC;
  SIGNAL yt_rsc_1_9_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_9_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_10_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_1_10_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_1_10_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_10_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_10_we : STD_LOGIC;
  SIGNAL yt_rsc_1_10_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_10_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_11_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_1_11_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_1_11_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_11_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_11_we : STD_LOGIC;
  SIGNAL yt_rsc_1_11_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_11_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_12_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_1_12_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_1_12_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_12_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_12_we : STD_LOGIC;
  SIGNAL yt_rsc_1_12_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_12_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_13_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_1_13_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_1_13_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_13_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_13_we : STD_LOGIC;
  SIGNAL yt_rsc_1_13_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_13_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_14_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_1_14_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_1_14_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_14_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_14_we : STD_LOGIC;
  SIGNAL yt_rsc_1_14_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_14_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_15_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_1_15_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_1_15_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_15_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_15_we : STD_LOGIC;
  SIGNAL yt_rsc_1_15_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_15_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_16_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_1_16_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_1_16_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_16_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_16_we : STD_LOGIC;
  SIGNAL yt_rsc_1_16_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_16_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_17_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_1_17_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_1_17_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_17_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_17_we : STD_LOGIC;
  SIGNAL yt_rsc_1_17_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_17_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_18_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_1_18_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_1_18_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_18_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_18_we : STD_LOGIC;
  SIGNAL yt_rsc_1_18_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_18_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_19_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_1_19_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_1_19_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_19_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_19_we : STD_LOGIC;
  SIGNAL yt_rsc_1_19_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_19_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_20_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_1_20_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_1_20_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_20_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_20_we : STD_LOGIC;
  SIGNAL yt_rsc_1_20_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_20_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_21_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_1_21_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_1_21_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_21_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_21_we : STD_LOGIC;
  SIGNAL yt_rsc_1_21_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_21_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_22_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_1_22_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_1_22_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_22_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_22_we : STD_LOGIC;
  SIGNAL yt_rsc_1_22_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_22_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_23_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_1_23_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_1_23_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_23_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_23_we : STD_LOGIC;
  SIGNAL yt_rsc_1_23_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_23_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_24_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_1_24_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_1_24_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_24_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_24_we : STD_LOGIC;
  SIGNAL yt_rsc_1_24_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_24_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_25_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_1_25_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_1_25_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_25_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_25_we : STD_LOGIC;
  SIGNAL yt_rsc_1_25_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_25_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_26_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_1_26_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_1_26_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_26_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_26_we : STD_LOGIC;
  SIGNAL yt_rsc_1_26_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_26_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_27_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_1_27_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_1_27_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_27_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_27_we : STD_LOGIC;
  SIGNAL yt_rsc_1_27_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_27_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_28_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_1_28_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_1_28_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_28_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_28_we : STD_LOGIC;
  SIGNAL yt_rsc_1_28_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_28_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_29_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_1_29_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_1_29_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_29_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_29_we : STD_LOGIC;
  SIGNAL yt_rsc_1_29_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_29_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_30_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_1_30_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_1_30_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_30_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_30_we : STD_LOGIC;
  SIGNAL yt_rsc_1_30_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_30_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_31_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_1_31_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_1_31_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_31_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_31_we : STD_LOGIC;
  SIGNAL yt_rsc_1_31_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_31_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_0_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_2_0_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_2_0_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_0_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_0_we : STD_LOGIC;
  SIGNAL yt_rsc_2_0_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_0_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_1_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_2_1_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_2_1_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_1_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_1_we : STD_LOGIC;
  SIGNAL yt_rsc_2_1_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_1_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_2_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_2_2_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_2_2_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_2_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_2_we : STD_LOGIC;
  SIGNAL yt_rsc_2_2_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_2_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_3_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_2_3_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_2_3_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_3_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_3_we : STD_LOGIC;
  SIGNAL yt_rsc_2_3_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_3_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_4_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_2_4_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_2_4_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_4_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_4_we : STD_LOGIC;
  SIGNAL yt_rsc_2_4_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_4_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_5_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_2_5_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_2_5_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_5_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_5_we : STD_LOGIC;
  SIGNAL yt_rsc_2_5_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_5_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_6_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_2_6_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_2_6_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_6_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_6_we : STD_LOGIC;
  SIGNAL yt_rsc_2_6_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_6_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_7_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_2_7_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_2_7_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_7_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_7_we : STD_LOGIC;
  SIGNAL yt_rsc_2_7_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_7_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_8_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_2_8_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_2_8_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_8_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_8_we : STD_LOGIC;
  SIGNAL yt_rsc_2_8_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_8_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_9_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_2_9_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_2_9_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_9_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_9_we : STD_LOGIC;
  SIGNAL yt_rsc_2_9_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_9_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_10_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_2_10_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_2_10_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_10_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_10_we : STD_LOGIC;
  SIGNAL yt_rsc_2_10_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_10_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_11_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_2_11_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_2_11_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_11_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_11_we : STD_LOGIC;
  SIGNAL yt_rsc_2_11_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_11_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_12_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_2_12_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_2_12_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_12_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_12_we : STD_LOGIC;
  SIGNAL yt_rsc_2_12_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_12_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_13_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_2_13_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_2_13_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_13_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_13_we : STD_LOGIC;
  SIGNAL yt_rsc_2_13_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_13_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_14_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_2_14_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_2_14_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_14_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_14_we : STD_LOGIC;
  SIGNAL yt_rsc_2_14_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_14_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_15_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_2_15_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_2_15_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_15_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_15_we : STD_LOGIC;
  SIGNAL yt_rsc_2_15_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_15_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_16_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_2_16_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_2_16_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_16_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_16_we : STD_LOGIC;
  SIGNAL yt_rsc_2_16_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_16_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_17_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_2_17_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_2_17_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_17_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_17_we : STD_LOGIC;
  SIGNAL yt_rsc_2_17_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_17_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_18_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_2_18_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_2_18_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_18_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_18_we : STD_LOGIC;
  SIGNAL yt_rsc_2_18_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_18_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_19_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_2_19_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_2_19_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_19_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_19_we : STD_LOGIC;
  SIGNAL yt_rsc_2_19_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_19_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_20_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_2_20_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_2_20_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_20_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_20_we : STD_LOGIC;
  SIGNAL yt_rsc_2_20_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_20_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_21_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_2_21_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_2_21_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_21_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_21_we : STD_LOGIC;
  SIGNAL yt_rsc_2_21_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_21_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_22_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_2_22_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_2_22_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_22_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_22_we : STD_LOGIC;
  SIGNAL yt_rsc_2_22_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_22_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_23_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_2_23_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_2_23_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_23_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_23_we : STD_LOGIC;
  SIGNAL yt_rsc_2_23_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_23_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_24_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_2_24_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_2_24_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_24_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_24_we : STD_LOGIC;
  SIGNAL yt_rsc_2_24_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_24_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_25_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_2_25_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_2_25_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_25_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_25_we : STD_LOGIC;
  SIGNAL yt_rsc_2_25_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_25_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_26_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_2_26_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_2_26_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_26_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_26_we : STD_LOGIC;
  SIGNAL yt_rsc_2_26_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_26_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_27_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_2_27_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_2_27_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_27_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_27_we : STD_LOGIC;
  SIGNAL yt_rsc_2_27_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_27_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_28_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_2_28_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_2_28_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_28_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_28_we : STD_LOGIC;
  SIGNAL yt_rsc_2_28_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_28_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_29_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_2_29_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_2_29_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_29_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_29_we : STD_LOGIC;
  SIGNAL yt_rsc_2_29_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_29_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_30_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_2_30_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_2_30_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_30_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_30_we : STD_LOGIC;
  SIGNAL yt_rsc_2_30_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_30_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_31_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_2_31_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_2_31_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_31_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_31_we : STD_LOGIC;
  SIGNAL yt_rsc_2_31_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_31_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_0_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_3_0_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_3_0_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_0_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_0_we : STD_LOGIC;
  SIGNAL yt_rsc_3_0_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_0_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_1_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_3_1_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_3_1_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_1_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_1_we : STD_LOGIC;
  SIGNAL yt_rsc_3_1_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_1_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_2_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_3_2_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_3_2_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_2_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_2_we : STD_LOGIC;
  SIGNAL yt_rsc_3_2_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_2_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_3_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_3_3_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_3_3_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_3_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_3_we : STD_LOGIC;
  SIGNAL yt_rsc_3_3_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_3_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_4_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_3_4_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_3_4_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_4_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_4_we : STD_LOGIC;
  SIGNAL yt_rsc_3_4_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_4_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_5_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_3_5_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_3_5_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_5_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_5_we : STD_LOGIC;
  SIGNAL yt_rsc_3_5_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_5_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_6_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_3_6_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_3_6_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_6_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_6_we : STD_LOGIC;
  SIGNAL yt_rsc_3_6_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_6_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_7_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_3_7_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_3_7_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_7_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_7_we : STD_LOGIC;
  SIGNAL yt_rsc_3_7_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_7_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_8_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_3_8_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_3_8_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_8_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_8_we : STD_LOGIC;
  SIGNAL yt_rsc_3_8_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_8_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_9_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_3_9_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_3_9_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_9_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_9_we : STD_LOGIC;
  SIGNAL yt_rsc_3_9_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_9_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_10_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_3_10_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_3_10_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_10_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_10_we : STD_LOGIC;
  SIGNAL yt_rsc_3_10_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_10_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_11_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_3_11_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_3_11_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_11_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_11_we : STD_LOGIC;
  SIGNAL yt_rsc_3_11_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_11_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_12_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_3_12_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_3_12_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_12_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_12_we : STD_LOGIC;
  SIGNAL yt_rsc_3_12_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_12_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_13_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_3_13_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_3_13_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_13_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_13_we : STD_LOGIC;
  SIGNAL yt_rsc_3_13_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_13_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_14_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_3_14_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_3_14_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_14_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_14_we : STD_LOGIC;
  SIGNAL yt_rsc_3_14_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_14_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_15_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_3_15_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_3_15_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_15_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_15_we : STD_LOGIC;
  SIGNAL yt_rsc_3_15_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_15_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_16_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_3_16_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_3_16_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_16_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_16_we : STD_LOGIC;
  SIGNAL yt_rsc_3_16_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_16_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_17_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_3_17_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_3_17_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_17_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_17_we : STD_LOGIC;
  SIGNAL yt_rsc_3_17_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_17_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_18_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_3_18_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_3_18_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_18_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_18_we : STD_LOGIC;
  SIGNAL yt_rsc_3_18_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_18_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_19_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_3_19_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_3_19_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_19_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_19_we : STD_LOGIC;
  SIGNAL yt_rsc_3_19_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_19_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_20_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_3_20_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_3_20_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_20_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_20_we : STD_LOGIC;
  SIGNAL yt_rsc_3_20_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_20_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_21_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_3_21_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_3_21_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_21_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_21_we : STD_LOGIC;
  SIGNAL yt_rsc_3_21_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_21_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_22_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_3_22_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_3_22_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_22_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_22_we : STD_LOGIC;
  SIGNAL yt_rsc_3_22_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_22_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_23_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_3_23_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_3_23_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_23_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_23_we : STD_LOGIC;
  SIGNAL yt_rsc_3_23_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_23_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_24_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_3_24_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_3_24_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_24_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_24_we : STD_LOGIC;
  SIGNAL yt_rsc_3_24_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_24_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_25_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_3_25_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_3_25_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_25_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_25_we : STD_LOGIC;
  SIGNAL yt_rsc_3_25_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_25_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_26_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_3_26_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_3_26_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_26_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_26_we : STD_LOGIC;
  SIGNAL yt_rsc_3_26_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_26_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_27_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_3_27_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_3_27_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_27_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_27_we : STD_LOGIC;
  SIGNAL yt_rsc_3_27_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_27_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_28_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_3_28_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_3_28_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_28_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_28_we : STD_LOGIC;
  SIGNAL yt_rsc_3_28_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_28_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_29_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_3_29_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_3_29_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_29_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_29_we : STD_LOGIC;
  SIGNAL yt_rsc_3_29_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_29_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_30_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_3_30_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_3_30_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_30_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_30_we : STD_LOGIC;
  SIGNAL yt_rsc_3_30_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_30_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_31_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_3_31_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_3_31_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_31_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_31_we : STD_LOGIC;
  SIGNAL yt_rsc_3_31_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_31_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_0_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_4_0_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_4_0_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_0_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_0_we : STD_LOGIC;
  SIGNAL yt_rsc_4_0_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_0_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_1_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_4_1_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_4_1_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_1_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_1_we : STD_LOGIC;
  SIGNAL yt_rsc_4_1_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_1_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_2_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_4_2_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_4_2_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_2_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_2_we : STD_LOGIC;
  SIGNAL yt_rsc_4_2_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_2_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_3_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_4_3_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_4_3_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_3_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_3_we : STD_LOGIC;
  SIGNAL yt_rsc_4_3_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_3_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_4_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_4_4_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_4_4_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_4_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_4_we : STD_LOGIC;
  SIGNAL yt_rsc_4_4_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_4_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_5_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_4_5_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_4_5_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_5_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_5_we : STD_LOGIC;
  SIGNAL yt_rsc_4_5_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_5_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_6_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_4_6_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_4_6_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_6_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_6_we : STD_LOGIC;
  SIGNAL yt_rsc_4_6_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_6_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_7_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_4_7_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_4_7_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_7_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_7_we : STD_LOGIC;
  SIGNAL yt_rsc_4_7_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_7_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_8_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_4_8_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_4_8_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_8_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_8_we : STD_LOGIC;
  SIGNAL yt_rsc_4_8_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_8_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_9_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_4_9_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_4_9_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_9_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_9_we : STD_LOGIC;
  SIGNAL yt_rsc_4_9_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_9_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_10_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_4_10_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_4_10_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_10_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_10_we : STD_LOGIC;
  SIGNAL yt_rsc_4_10_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_10_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_11_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_4_11_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_4_11_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_11_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_11_we : STD_LOGIC;
  SIGNAL yt_rsc_4_11_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_11_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_12_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_4_12_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_4_12_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_12_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_12_we : STD_LOGIC;
  SIGNAL yt_rsc_4_12_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_12_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_13_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_4_13_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_4_13_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_13_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_13_we : STD_LOGIC;
  SIGNAL yt_rsc_4_13_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_13_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_14_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_4_14_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_4_14_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_14_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_14_we : STD_LOGIC;
  SIGNAL yt_rsc_4_14_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_14_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_15_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_4_15_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_4_15_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_15_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_15_we : STD_LOGIC;
  SIGNAL yt_rsc_4_15_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_15_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_16_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_4_16_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_4_16_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_16_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_16_we : STD_LOGIC;
  SIGNAL yt_rsc_4_16_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_16_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_17_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_4_17_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_4_17_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_17_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_17_we : STD_LOGIC;
  SIGNAL yt_rsc_4_17_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_17_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_18_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_4_18_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_4_18_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_18_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_18_we : STD_LOGIC;
  SIGNAL yt_rsc_4_18_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_18_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_19_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_4_19_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_4_19_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_19_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_19_we : STD_LOGIC;
  SIGNAL yt_rsc_4_19_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_19_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_20_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_4_20_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_4_20_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_20_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_20_we : STD_LOGIC;
  SIGNAL yt_rsc_4_20_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_20_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_21_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_4_21_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_4_21_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_21_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_21_we : STD_LOGIC;
  SIGNAL yt_rsc_4_21_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_21_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_22_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_4_22_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_4_22_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_22_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_22_we : STD_LOGIC;
  SIGNAL yt_rsc_4_22_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_22_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_23_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_4_23_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_4_23_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_23_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_23_we : STD_LOGIC;
  SIGNAL yt_rsc_4_23_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_23_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_24_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_4_24_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_4_24_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_24_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_24_we : STD_LOGIC;
  SIGNAL yt_rsc_4_24_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_24_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_25_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_4_25_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_4_25_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_25_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_25_we : STD_LOGIC;
  SIGNAL yt_rsc_4_25_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_25_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_26_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_4_26_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_4_26_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_26_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_26_we : STD_LOGIC;
  SIGNAL yt_rsc_4_26_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_26_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_27_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_4_27_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_4_27_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_27_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_27_we : STD_LOGIC;
  SIGNAL yt_rsc_4_27_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_27_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_28_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_4_28_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_4_28_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_28_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_28_we : STD_LOGIC;
  SIGNAL yt_rsc_4_28_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_28_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_29_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_4_29_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_4_29_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_29_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_29_we : STD_LOGIC;
  SIGNAL yt_rsc_4_29_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_29_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_30_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_4_30_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_4_30_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_30_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_30_we : STD_LOGIC;
  SIGNAL yt_rsc_4_30_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_30_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_31_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_4_31_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_4_31_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_31_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_31_we : STD_LOGIC;
  SIGNAL yt_rsc_4_31_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_31_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_0_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_5_0_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_5_0_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_0_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_0_we : STD_LOGIC;
  SIGNAL yt_rsc_5_0_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_0_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_1_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_5_1_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_5_1_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_1_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_1_we : STD_LOGIC;
  SIGNAL yt_rsc_5_1_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_1_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_2_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_5_2_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_5_2_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_2_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_2_we : STD_LOGIC;
  SIGNAL yt_rsc_5_2_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_2_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_3_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_5_3_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_5_3_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_3_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_3_we : STD_LOGIC;
  SIGNAL yt_rsc_5_3_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_3_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_4_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_5_4_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_5_4_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_4_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_4_we : STD_LOGIC;
  SIGNAL yt_rsc_5_4_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_4_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_5_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_5_5_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_5_5_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_5_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_5_we : STD_LOGIC;
  SIGNAL yt_rsc_5_5_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_5_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_6_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_5_6_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_5_6_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_6_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_6_we : STD_LOGIC;
  SIGNAL yt_rsc_5_6_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_6_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_7_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_5_7_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_5_7_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_7_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_7_we : STD_LOGIC;
  SIGNAL yt_rsc_5_7_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_7_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_8_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_5_8_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_5_8_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_8_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_8_we : STD_LOGIC;
  SIGNAL yt_rsc_5_8_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_8_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_9_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_5_9_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_5_9_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_9_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_9_we : STD_LOGIC;
  SIGNAL yt_rsc_5_9_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_9_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_10_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_5_10_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_5_10_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_10_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_10_we : STD_LOGIC;
  SIGNAL yt_rsc_5_10_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_10_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_11_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_5_11_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_5_11_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_11_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_11_we : STD_LOGIC;
  SIGNAL yt_rsc_5_11_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_11_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_12_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_5_12_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_5_12_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_12_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_12_we : STD_LOGIC;
  SIGNAL yt_rsc_5_12_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_12_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_13_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_5_13_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_5_13_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_13_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_13_we : STD_LOGIC;
  SIGNAL yt_rsc_5_13_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_13_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_14_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_5_14_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_5_14_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_14_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_14_we : STD_LOGIC;
  SIGNAL yt_rsc_5_14_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_14_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_15_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_5_15_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_5_15_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_15_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_15_we : STD_LOGIC;
  SIGNAL yt_rsc_5_15_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_15_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_16_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_5_16_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_5_16_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_16_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_16_we : STD_LOGIC;
  SIGNAL yt_rsc_5_16_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_16_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_17_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_5_17_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_5_17_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_17_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_17_we : STD_LOGIC;
  SIGNAL yt_rsc_5_17_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_17_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_18_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_5_18_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_5_18_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_18_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_18_we : STD_LOGIC;
  SIGNAL yt_rsc_5_18_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_18_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_19_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_5_19_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_5_19_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_19_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_19_we : STD_LOGIC;
  SIGNAL yt_rsc_5_19_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_19_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_20_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_5_20_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_5_20_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_20_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_20_we : STD_LOGIC;
  SIGNAL yt_rsc_5_20_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_20_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_21_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_5_21_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_5_21_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_21_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_21_we : STD_LOGIC;
  SIGNAL yt_rsc_5_21_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_21_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_22_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_5_22_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_5_22_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_22_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_22_we : STD_LOGIC;
  SIGNAL yt_rsc_5_22_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_22_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_23_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_5_23_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_5_23_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_23_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_23_we : STD_LOGIC;
  SIGNAL yt_rsc_5_23_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_23_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_24_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_5_24_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_5_24_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_24_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_24_we : STD_LOGIC;
  SIGNAL yt_rsc_5_24_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_24_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_25_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_5_25_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_5_25_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_25_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_25_we : STD_LOGIC;
  SIGNAL yt_rsc_5_25_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_25_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_26_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_5_26_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_5_26_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_26_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_26_we : STD_LOGIC;
  SIGNAL yt_rsc_5_26_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_26_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_27_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_5_27_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_5_27_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_27_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_27_we : STD_LOGIC;
  SIGNAL yt_rsc_5_27_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_27_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_28_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_5_28_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_5_28_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_28_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_28_we : STD_LOGIC;
  SIGNAL yt_rsc_5_28_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_28_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_29_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_5_29_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_5_29_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_29_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_29_we : STD_LOGIC;
  SIGNAL yt_rsc_5_29_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_29_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_30_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_5_30_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_5_30_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_30_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_30_we : STD_LOGIC;
  SIGNAL yt_rsc_5_30_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_30_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_31_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_5_31_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_5_31_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_31_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_31_we : STD_LOGIC;
  SIGNAL yt_rsc_5_31_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_31_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_0_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_6_0_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_6_0_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_0_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_0_we : STD_LOGIC;
  SIGNAL yt_rsc_6_0_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_0_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_1_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_6_1_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_6_1_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_1_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_1_we : STD_LOGIC;
  SIGNAL yt_rsc_6_1_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_1_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_2_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_6_2_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_6_2_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_2_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_2_we : STD_LOGIC;
  SIGNAL yt_rsc_6_2_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_2_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_3_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_6_3_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_6_3_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_3_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_3_we : STD_LOGIC;
  SIGNAL yt_rsc_6_3_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_3_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_4_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_6_4_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_6_4_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_4_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_4_we : STD_LOGIC;
  SIGNAL yt_rsc_6_4_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_4_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_5_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_6_5_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_6_5_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_5_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_5_we : STD_LOGIC;
  SIGNAL yt_rsc_6_5_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_5_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_6_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_6_6_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_6_6_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_6_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_6_we : STD_LOGIC;
  SIGNAL yt_rsc_6_6_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_6_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_7_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_6_7_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_6_7_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_7_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_7_we : STD_LOGIC;
  SIGNAL yt_rsc_6_7_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_7_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_8_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_6_8_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_6_8_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_8_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_8_we : STD_LOGIC;
  SIGNAL yt_rsc_6_8_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_8_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_9_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_6_9_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_6_9_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_9_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_9_we : STD_LOGIC;
  SIGNAL yt_rsc_6_9_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_9_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_10_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_6_10_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_6_10_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_10_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_10_we : STD_LOGIC;
  SIGNAL yt_rsc_6_10_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_10_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_11_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_6_11_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_6_11_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_11_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_11_we : STD_LOGIC;
  SIGNAL yt_rsc_6_11_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_11_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_12_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_6_12_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_6_12_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_12_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_12_we : STD_LOGIC;
  SIGNAL yt_rsc_6_12_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_12_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_13_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_6_13_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_6_13_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_13_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_13_we : STD_LOGIC;
  SIGNAL yt_rsc_6_13_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_13_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_14_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_6_14_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_6_14_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_14_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_14_we : STD_LOGIC;
  SIGNAL yt_rsc_6_14_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_14_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_15_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_6_15_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_6_15_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_15_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_15_we : STD_LOGIC;
  SIGNAL yt_rsc_6_15_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_15_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_16_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_6_16_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_6_16_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_16_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_16_we : STD_LOGIC;
  SIGNAL yt_rsc_6_16_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_16_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_17_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_6_17_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_6_17_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_17_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_17_we : STD_LOGIC;
  SIGNAL yt_rsc_6_17_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_17_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_18_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_6_18_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_6_18_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_18_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_18_we : STD_LOGIC;
  SIGNAL yt_rsc_6_18_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_18_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_19_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_6_19_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_6_19_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_19_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_19_we : STD_LOGIC;
  SIGNAL yt_rsc_6_19_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_19_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_20_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_6_20_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_6_20_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_20_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_20_we : STD_LOGIC;
  SIGNAL yt_rsc_6_20_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_20_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_21_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_6_21_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_6_21_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_21_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_21_we : STD_LOGIC;
  SIGNAL yt_rsc_6_21_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_21_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_22_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_6_22_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_6_22_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_22_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_22_we : STD_LOGIC;
  SIGNAL yt_rsc_6_22_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_22_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_23_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_6_23_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_6_23_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_23_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_23_we : STD_LOGIC;
  SIGNAL yt_rsc_6_23_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_23_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_24_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_6_24_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_6_24_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_24_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_24_we : STD_LOGIC;
  SIGNAL yt_rsc_6_24_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_24_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_25_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_6_25_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_6_25_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_25_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_25_we : STD_LOGIC;
  SIGNAL yt_rsc_6_25_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_25_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_26_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_6_26_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_6_26_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_26_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_26_we : STD_LOGIC;
  SIGNAL yt_rsc_6_26_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_26_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_27_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_6_27_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_6_27_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_27_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_27_we : STD_LOGIC;
  SIGNAL yt_rsc_6_27_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_27_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_28_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_6_28_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_6_28_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_28_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_28_we : STD_LOGIC;
  SIGNAL yt_rsc_6_28_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_28_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_29_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_6_29_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_6_29_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_29_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_29_we : STD_LOGIC;
  SIGNAL yt_rsc_6_29_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_29_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_30_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_6_30_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_6_30_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_30_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_30_we : STD_LOGIC;
  SIGNAL yt_rsc_6_30_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_30_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_31_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_6_31_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_6_31_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_31_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_31_we : STD_LOGIC;
  SIGNAL yt_rsc_6_31_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_31_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_0_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_7_0_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_7_0_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_0_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_0_we : STD_LOGIC;
  SIGNAL yt_rsc_7_0_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_0_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_1_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_7_1_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_7_1_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_1_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_1_we : STD_LOGIC;
  SIGNAL yt_rsc_7_1_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_1_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_2_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_7_2_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_7_2_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_2_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_2_we : STD_LOGIC;
  SIGNAL yt_rsc_7_2_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_2_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_3_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_7_3_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_7_3_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_3_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_3_we : STD_LOGIC;
  SIGNAL yt_rsc_7_3_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_3_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_4_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_7_4_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_7_4_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_4_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_4_we : STD_LOGIC;
  SIGNAL yt_rsc_7_4_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_4_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_5_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_7_5_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_7_5_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_5_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_5_we : STD_LOGIC;
  SIGNAL yt_rsc_7_5_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_5_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_6_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_7_6_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_7_6_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_6_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_6_we : STD_LOGIC;
  SIGNAL yt_rsc_7_6_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_6_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_7_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_7_7_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_7_7_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_7_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_7_we : STD_LOGIC;
  SIGNAL yt_rsc_7_7_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_7_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_8_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_7_8_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_7_8_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_8_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_8_we : STD_LOGIC;
  SIGNAL yt_rsc_7_8_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_8_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_9_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_7_9_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_7_9_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_9_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_9_we : STD_LOGIC;
  SIGNAL yt_rsc_7_9_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_9_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_10_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_7_10_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_7_10_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_10_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_10_we : STD_LOGIC;
  SIGNAL yt_rsc_7_10_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_10_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_11_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_7_11_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_7_11_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_11_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_11_we : STD_LOGIC;
  SIGNAL yt_rsc_7_11_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_11_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_12_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_7_12_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_7_12_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_12_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_12_we : STD_LOGIC;
  SIGNAL yt_rsc_7_12_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_12_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_13_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_7_13_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_7_13_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_13_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_13_we : STD_LOGIC;
  SIGNAL yt_rsc_7_13_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_13_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_14_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_7_14_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_7_14_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_14_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_14_we : STD_LOGIC;
  SIGNAL yt_rsc_7_14_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_14_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_15_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_7_15_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_7_15_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_15_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_15_we : STD_LOGIC;
  SIGNAL yt_rsc_7_15_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_15_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_16_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_7_16_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_7_16_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_16_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_16_we : STD_LOGIC;
  SIGNAL yt_rsc_7_16_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_16_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_17_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_7_17_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_7_17_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_17_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_17_we : STD_LOGIC;
  SIGNAL yt_rsc_7_17_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_17_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_18_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_7_18_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_7_18_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_18_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_18_we : STD_LOGIC;
  SIGNAL yt_rsc_7_18_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_18_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_19_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_7_19_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_7_19_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_19_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_19_we : STD_LOGIC;
  SIGNAL yt_rsc_7_19_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_19_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_20_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_7_20_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_7_20_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_20_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_20_we : STD_LOGIC;
  SIGNAL yt_rsc_7_20_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_20_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_21_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_7_21_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_7_21_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_21_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_21_we : STD_LOGIC;
  SIGNAL yt_rsc_7_21_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_21_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_22_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_7_22_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_7_22_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_22_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_22_we : STD_LOGIC;
  SIGNAL yt_rsc_7_22_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_22_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_23_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_7_23_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_7_23_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_23_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_23_we : STD_LOGIC;
  SIGNAL yt_rsc_7_23_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_23_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_24_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_7_24_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_7_24_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_24_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_24_we : STD_LOGIC;
  SIGNAL yt_rsc_7_24_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_24_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_25_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_7_25_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_7_25_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_25_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_25_we : STD_LOGIC;
  SIGNAL yt_rsc_7_25_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_25_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_26_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_7_26_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_7_26_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_26_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_26_we : STD_LOGIC;
  SIGNAL yt_rsc_7_26_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_26_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_27_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_7_27_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_7_27_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_27_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_27_we : STD_LOGIC;
  SIGNAL yt_rsc_7_27_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_27_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_28_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_7_28_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_7_28_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_28_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_28_we : STD_LOGIC;
  SIGNAL yt_rsc_7_28_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_28_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_29_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_7_29_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_7_29_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_29_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_29_we : STD_LOGIC;
  SIGNAL yt_rsc_7_29_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_29_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_30_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_7_30_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_7_30_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_30_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_30_we : STD_LOGIC;
  SIGNAL yt_rsc_7_30_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_30_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_31_clkr_en : STD_LOGIC;
  SIGNAL yt_rsc_7_31_clkw_en : STD_LOGIC;
  SIGNAL yt_rsc_7_31_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_31_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_31_we : STD_LOGIC;
  SIGNAL yt_rsc_7_31_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_31_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_0_i_d_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_0_i_radr_d_iff : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_0_i_wadr_d_iff : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_0_i_we_d_iff : STD_LOGIC;
  SIGNAL yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff : STD_LOGIC;
  SIGNAL yt_rsc_0_1_i_d_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_1_i_wadr_d_iff : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_2_i_d_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_2_i_wadr_d_iff : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_3_i_d_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_3_i_wadr_d_iff : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_4_i_d_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_4_i_wadr_d_iff : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_5_i_d_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_5_i_wadr_d_iff : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_6_i_d_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_6_i_wadr_d_iff : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_7_i_d_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_8_i_d_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_9_i_d_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_10_i_d_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_10_i_wadr_d_iff : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_11_i_d_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_11_i_wadr_d_iff : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_12_i_d_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_13_i_d_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_14_i_d_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_15_i_d_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_16_i_we_d_iff : STD_LOGIC;
  SIGNAL yt_rsc_1_0_i_we_d_iff : STD_LOGIC;
  SIGNAL yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff : STD_LOGIC;
  SIGNAL yt_rsc_1_16_i_we_d_iff : STD_LOGIC;
  SIGNAL yt_rsc_2_0_i_we_d_iff : STD_LOGIC;
  SIGNAL yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff : STD_LOGIC;
  SIGNAL yt_rsc_2_16_i_we_d_iff : STD_LOGIC;
  SIGNAL yt_rsc_3_0_i_we_d_iff : STD_LOGIC;
  SIGNAL yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff : STD_LOGIC;
  SIGNAL yt_rsc_3_16_i_we_d_iff : STD_LOGIC;
  SIGNAL yt_rsc_4_0_i_d_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_0_i_wadr_d_iff : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_0_i_we_d_iff : STD_LOGIC;
  SIGNAL yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff : STD_LOGIC;
  SIGNAL yt_rsc_4_1_i_d_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_1_i_wadr_d_iff : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_2_i_d_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_2_i_wadr_d_iff : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_3_i_d_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_3_i_wadr_d_iff : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_4_i_d_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_4_i_wadr_d_iff : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_5_i_d_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_5_i_wadr_d_iff : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_6_i_d_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_6_i_wadr_d_iff : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_7_i_d_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_8_i_d_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_9_i_d_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_9_i_wadr_d_iff : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_10_i_d_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_10_i_wadr_d_iff : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_11_i_d_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_11_i_wadr_d_iff : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_12_i_d_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_13_i_d_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_14_i_d_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_15_i_d_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_16_i_we_d_iff : STD_LOGIC;
  SIGNAL yt_rsc_5_0_i_we_d_iff : STD_LOGIC;
  SIGNAL yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff : STD_LOGIC;
  SIGNAL yt_rsc_5_16_i_we_d_iff : STD_LOGIC;
  SIGNAL yt_rsc_6_0_i_we_d_iff : STD_LOGIC;
  SIGNAL yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff : STD_LOGIC;
  SIGNAL yt_rsc_6_16_i_we_d_iff : STD_LOGIC;
  SIGNAL yt_rsc_7_0_i_we_d_iff : STD_LOGIC;
  SIGNAL yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff : STD_LOGIC;
  SIGNAL yt_rsc_7_16_i_we_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_0_0_i_adra_d_iff : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_0_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_0_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_0_1_i_adra_d_iff : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_1_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_2_i_adra_d_iff : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_2_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_3_i_adra_d_iff : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_3_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_4_i_adra_d_iff : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_4_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_5_i_adra_d_iff : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_5_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_6_i_adra_d_iff : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_6_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_7_i_adra_d_iff : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_7_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_8_i_adra_d_iff : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_8_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_9_i_adra_d_iff : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_9_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_10_i_adra_d_iff : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_10_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_11_i_adra_d_iff : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_11_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_12_i_adra_d_iff : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_12_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_13_i_adra_d_iff : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_13_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_14_i_adra_d_iff : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_14_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_15_i_adra_d_iff : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_15_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_16_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_1_0_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_1_16_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_2_0_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_2_16_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_3_0_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_3_16_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_4_0_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_4_1_i_adra_d_iff : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_1_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_2_i_adra_d_iff : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_2_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_3_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_4_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_5_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_6_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_7_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_8_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_9_i_adra_d_iff : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_9_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_10_i_adra_d_iff : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_10_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_11_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_12_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_13_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_14_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_15_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff : STD_LOGIC;

  SIGNAL yt_rsc_0_0_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_0_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_0_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_0_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_0_1_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_1_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_1_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_1_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_0_2_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_2_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_2_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_2_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_0_3_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_3_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_3_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_3_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_0_4_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_4_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_4_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_4_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_0_5_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_5_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_5_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_5_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_0_6_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_6_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_6_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_6_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_0_7_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_7_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_7_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_7_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_0_8_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_8_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_8_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_8_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_0_9_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_9_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_9_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_9_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_0_10_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_10_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_10_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_10_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_0_11_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_11_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_11_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_11_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_0_12_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_12_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_12_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_12_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_0_13_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_13_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_13_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_13_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_0_14_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_14_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_14_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_14_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_0_15_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_15_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_15_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_15_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_0_16_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_16_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_16_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_16_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_0_17_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_17_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_17_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_17_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_0_18_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_18_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_18_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_18_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_0_19_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_19_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_19_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_19_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_0_20_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_20_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_20_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_20_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_0_21_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_21_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_21_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_21_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_0_22_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_22_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_22_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_22_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_0_23_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_23_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_23_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_23_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_0_24_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_24_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_24_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_24_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_0_25_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_25_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_25_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_25_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_0_26_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_26_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_26_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_26_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_0_27_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_27_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_27_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_27_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_0_28_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_28_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_28_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_28_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_0_29_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_29_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_29_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_29_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_0_30_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_30_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_30_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_30_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_0_31_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_31_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_31_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_31_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_1_0_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_0_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_0_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_0_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_1_1_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_1_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_1_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_1_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_1_2_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_2_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_2_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_2_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_1_3_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_3_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_3_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_3_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_1_4_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_4_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_4_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_4_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_1_5_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_5_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_5_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_5_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_1_6_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_6_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_6_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_6_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_1_7_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_7_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_7_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_7_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_1_8_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_8_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_8_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_8_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_1_9_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_9_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_9_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_9_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_1_10_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_10_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_10_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_10_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_1_11_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_11_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_11_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_11_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_1_12_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_12_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_12_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_12_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_1_13_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_13_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_13_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_13_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_1_14_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_14_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_14_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_14_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_1_15_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_15_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_15_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_15_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_1_16_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_16_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_16_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_16_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_1_17_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_17_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_17_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_17_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_1_18_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_18_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_18_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_18_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_1_19_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_19_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_19_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_19_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_1_20_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_20_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_20_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_20_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_1_21_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_21_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_21_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_21_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_1_22_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_22_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_22_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_22_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_1_23_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_23_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_23_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_23_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_1_24_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_24_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_24_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_24_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_1_25_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_25_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_25_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_25_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_1_26_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_26_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_26_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_26_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_1_27_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_27_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_27_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_27_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_1_28_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_28_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_28_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_28_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_1_29_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_29_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_29_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_29_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_1_30_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_30_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_30_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_30_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_1_31_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_31_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_31_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_31_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_2_0_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_0_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_0_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_0_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_2_1_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_1_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_1_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_1_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_2_2_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_2_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_2_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_2_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_2_3_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_3_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_3_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_3_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_2_4_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_4_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_4_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_4_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_2_5_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_5_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_5_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_5_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_2_6_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_6_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_6_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_6_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_2_7_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_7_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_7_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_7_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_2_8_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_8_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_8_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_8_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_2_9_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_9_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_9_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_9_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_2_10_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_10_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_10_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_10_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_2_11_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_11_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_11_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_11_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_2_12_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_12_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_12_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_12_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_2_13_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_13_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_13_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_13_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_2_14_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_14_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_14_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_14_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_2_15_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_15_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_15_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_15_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_2_16_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_16_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_16_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_16_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_2_17_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_17_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_17_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_17_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_2_18_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_18_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_18_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_18_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_2_19_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_19_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_19_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_19_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_2_20_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_20_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_20_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_20_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_2_21_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_21_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_21_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_21_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_2_22_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_22_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_22_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_22_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_2_23_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_23_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_23_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_23_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_2_24_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_24_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_24_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_24_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_2_25_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_25_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_25_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_25_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_2_26_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_26_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_26_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_26_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_2_27_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_27_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_27_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_27_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_2_28_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_28_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_28_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_28_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_2_29_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_29_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_29_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_29_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_2_30_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_30_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_30_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_30_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_2_31_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_31_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_31_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_31_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_3_0_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_0_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_0_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_0_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_3_1_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_1_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_1_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_1_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_3_2_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_2_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_2_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_2_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_3_3_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_3_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_3_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_3_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_3_4_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_4_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_4_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_4_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_3_5_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_5_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_5_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_5_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_3_6_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_6_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_6_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_6_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_3_7_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_7_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_7_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_7_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_3_8_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_8_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_8_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_8_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_3_9_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_9_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_9_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_9_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_3_10_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_10_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_10_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_10_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_3_11_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_11_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_11_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_11_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_3_12_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_12_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_12_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_12_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_3_13_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_13_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_13_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_13_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_3_14_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_14_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_14_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_14_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_3_15_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_15_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_15_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_15_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_3_16_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_16_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_16_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_16_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_3_17_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_17_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_17_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_17_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_3_18_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_18_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_18_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_18_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_3_19_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_19_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_19_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_19_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_3_20_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_20_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_20_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_20_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_3_21_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_21_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_21_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_21_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_3_22_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_22_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_22_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_22_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_3_23_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_23_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_23_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_23_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_3_24_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_24_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_24_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_24_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_3_25_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_25_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_25_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_25_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_3_26_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_26_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_26_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_26_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_3_27_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_27_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_27_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_27_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_3_28_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_28_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_28_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_28_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_3_29_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_29_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_29_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_29_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_3_30_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_30_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_30_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_30_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_3_31_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_31_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_31_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_31_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_4_0_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_0_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_0_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_0_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_4_1_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_1_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_1_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_1_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_4_2_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_2_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_2_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_2_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_4_3_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_3_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_3_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_3_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_4_4_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_4_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_4_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_4_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_4_5_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_5_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_5_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_5_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_4_6_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_6_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_6_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_6_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_4_7_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_7_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_7_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_7_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_4_8_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_8_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_8_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_8_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_4_9_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_9_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_9_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_9_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_4_10_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_10_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_10_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_10_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_4_11_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_11_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_11_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_11_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_4_12_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_12_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_12_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_12_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_4_13_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_13_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_13_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_13_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_4_14_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_14_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_14_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_14_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_4_15_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_15_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_15_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_15_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_4_16_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_16_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_16_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_16_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_4_17_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_17_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_17_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_17_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_4_18_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_18_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_18_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_18_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_4_19_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_19_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_19_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_19_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_4_20_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_20_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_20_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_20_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_4_21_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_21_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_21_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_21_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_4_22_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_22_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_22_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_22_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_4_23_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_23_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_23_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_23_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_4_24_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_24_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_24_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_24_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_4_25_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_25_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_25_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_25_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_4_26_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_26_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_26_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_26_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_4_27_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_27_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_27_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_27_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_4_28_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_28_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_28_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_28_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_4_29_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_29_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_29_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_29_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_4_30_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_30_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_30_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_30_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_4_31_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_31_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_31_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_31_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_5_0_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_0_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_0_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_0_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_5_1_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_1_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_1_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_1_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_5_2_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_2_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_2_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_2_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_5_3_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_3_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_3_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_3_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_5_4_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_4_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_4_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_4_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_5_5_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_5_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_5_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_5_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_5_6_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_6_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_6_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_6_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_5_7_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_7_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_7_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_7_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_5_8_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_8_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_8_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_8_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_5_9_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_9_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_9_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_9_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_5_10_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_10_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_10_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_10_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_5_11_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_11_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_11_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_11_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_5_12_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_12_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_12_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_12_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_5_13_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_13_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_13_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_13_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_5_14_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_14_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_14_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_14_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_5_15_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_15_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_15_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_15_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_5_16_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_16_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_16_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_16_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_5_17_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_17_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_17_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_17_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_5_18_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_18_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_18_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_18_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_5_19_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_19_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_19_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_19_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_5_20_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_20_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_20_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_20_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_5_21_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_21_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_21_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_21_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_5_22_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_22_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_22_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_22_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_5_23_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_23_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_23_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_23_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_5_24_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_24_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_24_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_24_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_5_25_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_25_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_25_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_25_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_5_26_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_26_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_26_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_26_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_5_27_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_27_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_27_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_27_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_5_28_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_28_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_28_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_28_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_5_29_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_29_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_29_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_29_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_5_30_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_30_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_30_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_30_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_5_31_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_31_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_31_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_31_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_6_0_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_0_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_0_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_0_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_6_1_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_1_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_1_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_1_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_6_2_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_2_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_2_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_2_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_6_3_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_3_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_3_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_3_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_6_4_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_4_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_4_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_4_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_6_5_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_5_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_5_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_5_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_6_6_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_6_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_6_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_6_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_6_7_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_7_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_7_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_7_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_6_8_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_8_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_8_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_8_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_6_9_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_9_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_9_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_9_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_6_10_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_10_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_10_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_10_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_6_11_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_11_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_11_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_11_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_6_12_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_12_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_12_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_12_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_6_13_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_13_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_13_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_13_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_6_14_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_14_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_14_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_14_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_6_15_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_15_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_15_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_15_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_6_16_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_16_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_16_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_16_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_6_17_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_17_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_17_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_17_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_6_18_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_18_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_18_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_18_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_6_19_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_19_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_19_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_19_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_6_20_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_20_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_20_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_20_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_6_21_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_21_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_21_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_21_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_6_22_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_22_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_22_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_22_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_6_23_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_23_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_23_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_23_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_6_24_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_24_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_24_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_24_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_6_25_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_25_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_25_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_25_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_6_26_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_26_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_26_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_26_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_6_27_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_27_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_27_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_27_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_6_28_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_28_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_28_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_28_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_6_29_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_29_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_29_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_29_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_6_30_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_30_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_30_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_30_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_6_31_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_31_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_31_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_31_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_7_0_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_0_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_0_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_0_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_7_1_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_1_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_1_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_1_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_7_2_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_2_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_2_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_2_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_7_3_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_3_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_3_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_3_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_7_4_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_4_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_4_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_4_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_7_5_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_5_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_5_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_5_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_7_6_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_6_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_6_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_6_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_7_7_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_7_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_7_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_7_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_7_8_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_8_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_8_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_8_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_7_9_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_9_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_9_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_9_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_7_10_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_10_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_10_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_10_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_7_11_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_11_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_11_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_11_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_7_12_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_12_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_12_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_12_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_7_13_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_13_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_13_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_13_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_7_14_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_14_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_14_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_14_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_7_15_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_15_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_15_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_15_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_7_16_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_16_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_16_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_16_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_7_17_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_17_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_17_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_17_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_7_18_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_18_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_18_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_18_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_7_19_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_19_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_19_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_19_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_7_20_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_20_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_20_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_20_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_7_21_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_21_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_21_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_21_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_7_22_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_22_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_22_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_22_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_7_23_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_23_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_23_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_23_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_7_24_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_24_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_24_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_24_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_7_25_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_25_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_25_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_25_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_7_26_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_26_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_26_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_26_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_7_27_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_27_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_27_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_27_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_7_28_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_28_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_28_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_28_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_7_29_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_29_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_29_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_29_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_7_30_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_30_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_30_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_30_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  SIGNAL yt_rsc_7_31_comp_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_31_comp_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_31_comp_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_31_comp_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_7_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_0_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_0_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_0_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_0_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_0_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_0_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_0_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_0_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_8_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_1_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_1_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_1_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_1_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_1_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_1_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_1_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_1_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_9_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_2_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_2_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_2_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_2_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_2_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_2_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_2_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_2_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_10_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_3_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_3_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_3_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_3_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_3_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_3_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_3_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_3_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_11_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_4_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_4_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_4_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_4_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_4_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_4_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_4_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_4_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_12_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_5_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_5_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_5_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_5_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_5_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_5_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_5_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_5_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_13_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_6_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_6_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_6_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_6_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_6_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_6_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_6_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_6_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_14_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_7_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_7_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_7_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_7_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_7_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_7_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_7_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_7_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_15_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_8_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_8_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_8_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_8_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_8_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_8_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_8_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_8_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_16_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_9_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_9_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_9_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_9_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_9_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_9_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_9_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_9_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_17_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_10_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_10_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_10_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_10_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_10_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_10_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_10_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_10_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_18_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_11_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_11_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_11_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_11_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_11_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_11_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_11_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_11_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_19_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_12_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_12_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_12_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_12_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_12_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_12_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_12_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_12_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_20_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_13_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_13_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_13_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_13_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_13_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_13_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_13_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_13_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_21_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_14_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_14_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_14_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_14_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_14_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_14_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_14_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_14_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_22_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_15_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_15_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_15_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_15_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_15_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_15_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_15_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_15_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_23_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_16_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_16_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_16_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_16_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_16_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_16_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_16_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_16_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_24_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_17_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_17_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_17_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_17_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_17_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_17_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_17_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_17_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_25_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_18_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_18_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_18_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_18_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_18_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_18_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_18_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_18_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_26_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_19_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_19_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_19_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_19_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_19_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_19_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_19_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_19_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_27_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_20_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_20_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_20_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_20_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_20_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_20_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_20_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_20_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_28_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_21_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_21_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_21_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_21_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_21_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_21_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_21_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_21_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_29_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_22_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_22_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_22_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_22_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_22_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_22_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_22_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_22_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_30_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_23_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_23_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_23_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_23_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_23_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_23_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_23_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_23_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_31_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_24_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_24_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_24_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_24_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_24_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_24_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_24_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_24_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_32_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_25_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_25_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_25_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_25_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_25_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_25_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_25_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_25_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_33_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_26_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_26_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_26_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_26_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_26_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_26_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_26_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_26_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_34_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_27_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_27_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_27_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_27_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_27_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_27_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_27_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_27_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_35_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_28_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_28_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_28_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_28_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_28_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_28_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_28_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_28_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_36_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_29_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_29_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_29_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_29_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_29_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_29_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_29_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_29_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_37_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_30_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_30_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_30_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_30_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_30_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_30_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_30_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_30_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_38_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_31_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_31_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_31_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_31_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_31_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_31_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_31_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_31_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_39_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_1_0_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_0_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_0_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_0_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_0_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_0_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_0_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_0_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_40_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_1_1_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_1_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_1_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_1_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_1_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_1_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_1_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_1_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_41_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_1_2_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_2_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_2_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_2_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_2_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_2_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_2_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_2_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_42_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_1_3_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_3_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_3_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_3_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_3_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_3_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_3_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_3_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_43_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_1_4_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_4_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_4_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_4_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_4_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_4_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_4_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_4_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_44_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_1_5_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_5_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_5_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_5_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_5_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_5_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_5_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_5_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_45_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_1_6_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_6_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_6_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_6_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_6_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_6_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_6_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_6_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_46_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_1_7_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_7_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_7_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_7_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_7_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_7_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_7_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_7_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_47_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_1_8_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_8_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_8_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_8_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_8_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_8_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_8_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_8_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_48_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_1_9_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_9_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_9_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_9_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_9_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_9_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_9_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_9_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_49_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_1_10_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_10_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_10_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_10_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_10_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_10_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_10_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_10_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_50_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_1_11_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_11_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_11_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_11_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_11_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_11_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_11_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_11_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_51_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_1_12_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_12_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_12_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_12_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_12_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_12_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_12_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_12_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_52_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_1_13_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_13_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_13_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_13_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_13_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_13_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_13_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_13_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_53_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_1_14_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_14_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_14_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_14_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_14_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_14_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_14_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_14_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_54_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_1_15_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_15_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_15_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_15_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_15_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_15_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_15_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_15_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_55_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_1_16_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_16_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_16_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_16_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_16_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_16_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_16_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_16_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_56_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_1_17_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_17_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_17_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_17_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_17_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_17_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_17_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_17_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_57_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_1_18_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_18_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_18_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_18_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_18_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_18_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_18_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_18_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_58_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_1_19_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_19_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_19_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_19_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_19_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_19_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_19_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_19_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_59_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_1_20_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_20_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_20_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_20_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_20_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_20_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_20_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_20_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_60_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_1_21_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_21_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_21_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_21_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_21_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_21_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_21_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_21_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_61_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_1_22_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_22_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_22_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_22_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_22_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_22_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_22_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_22_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_62_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_1_23_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_23_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_23_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_23_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_23_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_23_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_23_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_23_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_63_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_1_24_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_24_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_24_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_24_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_24_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_24_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_24_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_24_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_64_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_1_25_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_25_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_25_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_25_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_25_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_25_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_25_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_25_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_65_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_1_26_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_26_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_26_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_26_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_26_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_26_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_26_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_26_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_66_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_1_27_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_27_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_27_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_27_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_27_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_27_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_27_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_27_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_67_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_1_28_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_28_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_28_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_28_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_28_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_28_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_28_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_28_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_68_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_1_29_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_29_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_29_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_29_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_29_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_29_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_29_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_29_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_69_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_1_30_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_30_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_30_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_30_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_30_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_30_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_30_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_30_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_70_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_1_31_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_31_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_31_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_31_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_31_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_31_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_31_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_31_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_71_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_2_0_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_0_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_0_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_0_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_0_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_0_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_0_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_0_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_72_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_2_1_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_1_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_1_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_1_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_1_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_1_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_1_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_1_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_73_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_2_2_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_2_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_2_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_2_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_2_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_2_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_2_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_2_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_74_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_2_3_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_3_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_3_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_3_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_3_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_3_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_3_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_3_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_75_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_2_4_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_4_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_4_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_4_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_4_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_4_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_4_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_4_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_76_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_2_5_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_5_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_5_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_5_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_5_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_5_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_5_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_5_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_77_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_2_6_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_6_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_6_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_6_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_6_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_6_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_6_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_6_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_78_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_2_7_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_7_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_7_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_7_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_7_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_7_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_7_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_7_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_79_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_2_8_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_8_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_8_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_8_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_8_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_8_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_8_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_8_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_80_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_2_9_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_9_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_9_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_9_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_9_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_9_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_9_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_9_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_81_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_2_10_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_10_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_10_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_10_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_10_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_10_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_10_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_10_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_82_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_2_11_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_11_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_11_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_11_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_11_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_11_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_11_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_11_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_83_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_2_12_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_12_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_12_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_12_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_12_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_12_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_12_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_12_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_84_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_2_13_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_13_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_13_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_13_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_13_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_13_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_13_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_13_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_85_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_2_14_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_14_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_14_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_14_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_14_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_14_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_14_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_14_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_86_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_2_15_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_15_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_15_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_15_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_15_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_15_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_15_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_15_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_87_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_2_16_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_16_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_16_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_16_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_16_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_16_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_16_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_16_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_88_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_2_17_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_17_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_17_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_17_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_17_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_17_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_17_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_17_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_89_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_2_18_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_18_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_18_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_18_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_18_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_18_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_18_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_18_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_90_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_2_19_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_19_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_19_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_19_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_19_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_19_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_19_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_19_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_91_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_2_20_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_20_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_20_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_20_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_20_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_20_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_20_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_20_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_92_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_2_21_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_21_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_21_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_21_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_21_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_21_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_21_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_21_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_93_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_2_22_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_22_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_22_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_22_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_22_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_22_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_22_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_22_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_94_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_2_23_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_23_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_23_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_23_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_23_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_23_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_23_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_23_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_95_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_2_24_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_24_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_24_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_24_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_24_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_24_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_24_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_24_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_96_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_2_25_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_25_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_25_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_25_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_25_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_25_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_25_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_25_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_97_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_2_26_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_26_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_26_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_26_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_26_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_26_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_26_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_26_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_98_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_2_27_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_27_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_27_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_27_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_27_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_27_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_27_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_27_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_99_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_2_28_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_28_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_28_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_28_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_28_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_28_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_28_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_28_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_100_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_2_29_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_29_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_29_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_29_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_29_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_29_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_29_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_29_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_101_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_2_30_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_30_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_30_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_30_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_30_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_30_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_30_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_30_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_102_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_2_31_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_31_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_31_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_31_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_31_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_31_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_2_31_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_2_31_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_103_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_3_0_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_0_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_0_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_0_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_0_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_0_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_0_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_0_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_104_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_3_1_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_1_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_1_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_1_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_1_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_1_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_1_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_1_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_105_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_3_2_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_2_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_2_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_2_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_2_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_2_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_2_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_2_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_106_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_3_3_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_3_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_3_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_3_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_3_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_3_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_3_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_3_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_107_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_3_4_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_4_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_4_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_4_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_4_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_4_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_4_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_4_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_108_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_3_5_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_5_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_5_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_5_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_5_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_5_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_5_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_5_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_109_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_3_6_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_6_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_6_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_6_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_6_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_6_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_6_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_6_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_110_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_3_7_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_7_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_7_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_7_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_7_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_7_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_7_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_7_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_111_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_3_8_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_8_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_8_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_8_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_8_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_8_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_8_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_8_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_112_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_3_9_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_9_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_9_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_9_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_9_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_9_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_9_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_9_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_113_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_3_10_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_10_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_10_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_10_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_10_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_10_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_10_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_10_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_114_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_3_11_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_11_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_11_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_11_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_11_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_11_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_11_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_11_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_115_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_3_12_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_12_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_12_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_12_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_12_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_12_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_12_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_12_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_116_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_3_13_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_13_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_13_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_13_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_13_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_13_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_13_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_13_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_117_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_3_14_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_14_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_14_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_14_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_14_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_14_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_14_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_14_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_118_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_3_15_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_15_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_15_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_15_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_15_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_15_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_15_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_15_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_119_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_3_16_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_16_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_16_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_16_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_16_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_16_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_16_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_16_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_120_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_3_17_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_17_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_17_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_17_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_17_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_17_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_17_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_17_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_121_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_3_18_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_18_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_18_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_18_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_18_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_18_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_18_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_18_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_122_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_3_19_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_19_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_19_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_19_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_19_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_19_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_19_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_19_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_123_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_3_20_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_20_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_20_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_20_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_20_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_20_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_20_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_20_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_124_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_3_21_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_21_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_21_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_21_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_21_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_21_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_21_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_21_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_125_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_3_22_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_22_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_22_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_22_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_22_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_22_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_22_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_22_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_126_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_3_23_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_23_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_23_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_23_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_23_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_23_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_23_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_23_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_127_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_3_24_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_24_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_24_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_24_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_24_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_24_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_24_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_24_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_128_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_3_25_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_25_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_25_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_25_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_25_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_25_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_25_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_25_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_129_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_3_26_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_26_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_26_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_26_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_26_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_26_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_26_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_26_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_130_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_3_27_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_27_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_27_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_27_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_27_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_27_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_27_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_27_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_131_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_3_28_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_28_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_28_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_28_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_28_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_28_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_28_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_28_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_132_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_3_29_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_29_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_29_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_29_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_29_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_29_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_29_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_29_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_133_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_3_30_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_30_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_30_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_30_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_30_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_30_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_30_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_30_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_134_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_3_31_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_31_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_31_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_31_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_31_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_31_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_3_31_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_3_31_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_135_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_4_0_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_0_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_0_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_0_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_0_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_0_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_0_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_0_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_136_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_4_1_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_1_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_1_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_1_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_1_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_1_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_1_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_1_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_137_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_4_2_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_2_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_2_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_2_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_2_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_2_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_2_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_2_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_138_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_4_3_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_3_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_3_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_3_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_3_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_3_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_3_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_3_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_139_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_4_4_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_4_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_4_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_4_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_4_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_4_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_4_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_4_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_140_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_4_5_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_5_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_5_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_5_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_5_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_5_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_5_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_5_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_141_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_4_6_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_6_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_6_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_6_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_6_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_6_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_6_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_6_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_142_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_4_7_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_7_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_7_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_7_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_7_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_7_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_7_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_7_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_143_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_4_8_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_8_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_8_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_8_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_8_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_8_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_8_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_8_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_144_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_4_9_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_9_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_9_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_9_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_9_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_9_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_9_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_9_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_145_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_4_10_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_10_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_10_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_10_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_10_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_10_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_10_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_10_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_146_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_4_11_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_11_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_11_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_11_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_11_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_11_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_11_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_11_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_147_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_4_12_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_12_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_12_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_12_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_12_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_12_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_12_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_12_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_148_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_4_13_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_13_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_13_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_13_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_13_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_13_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_13_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_13_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_149_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_4_14_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_14_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_14_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_14_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_14_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_14_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_14_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_14_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_150_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_4_15_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_15_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_15_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_15_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_15_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_15_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_15_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_15_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_151_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_4_16_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_16_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_16_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_16_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_16_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_16_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_16_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_16_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_152_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_4_17_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_17_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_17_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_17_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_17_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_17_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_17_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_17_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_153_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_4_18_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_18_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_18_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_18_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_18_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_18_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_18_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_18_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_154_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_4_19_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_19_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_19_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_19_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_19_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_19_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_19_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_19_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_155_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_4_20_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_20_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_20_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_20_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_20_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_20_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_20_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_20_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_156_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_4_21_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_21_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_21_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_21_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_21_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_21_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_21_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_21_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_157_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_4_22_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_22_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_22_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_22_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_22_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_22_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_22_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_22_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_158_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_4_23_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_23_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_23_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_23_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_23_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_23_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_23_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_23_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_159_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_4_24_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_24_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_24_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_24_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_24_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_24_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_24_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_24_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_160_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_4_25_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_25_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_25_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_25_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_25_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_25_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_25_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_25_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_161_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_4_26_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_26_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_26_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_26_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_26_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_26_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_26_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_26_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_162_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_4_27_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_27_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_27_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_27_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_27_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_27_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_27_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_27_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_163_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_4_28_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_28_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_28_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_28_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_28_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_28_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_28_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_28_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_164_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_4_29_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_29_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_29_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_29_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_29_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_29_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_29_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_29_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_165_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_4_30_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_30_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_30_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_30_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_30_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_30_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_30_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_30_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_166_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_4_31_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_31_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_31_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_31_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_31_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_31_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_4_31_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_4_31_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_167_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_5_0_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_0_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_0_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_0_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_0_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_0_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_0_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_0_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_168_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_5_1_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_1_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_1_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_1_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_1_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_1_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_1_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_1_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_169_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_5_2_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_2_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_2_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_2_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_2_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_2_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_2_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_2_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_170_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_5_3_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_3_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_3_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_3_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_3_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_3_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_3_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_3_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_171_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_5_4_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_4_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_4_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_4_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_4_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_4_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_4_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_4_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_172_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_5_5_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_5_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_5_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_5_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_5_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_5_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_5_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_5_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_173_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_5_6_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_6_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_6_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_6_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_6_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_6_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_6_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_6_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_174_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_5_7_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_7_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_7_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_7_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_7_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_7_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_7_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_7_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_175_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_5_8_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_8_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_8_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_8_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_8_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_8_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_8_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_8_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_176_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_5_9_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_9_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_9_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_9_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_9_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_9_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_9_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_9_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_177_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_5_10_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_10_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_10_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_10_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_10_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_10_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_10_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_10_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_178_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_5_11_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_11_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_11_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_11_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_11_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_11_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_11_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_11_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_179_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_5_12_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_12_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_12_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_12_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_12_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_12_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_12_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_12_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_180_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_5_13_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_13_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_13_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_13_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_13_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_13_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_13_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_13_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_181_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_5_14_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_14_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_14_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_14_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_14_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_14_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_14_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_14_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_182_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_5_15_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_15_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_15_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_15_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_15_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_15_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_15_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_15_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_183_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_5_16_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_16_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_16_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_16_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_16_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_16_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_16_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_16_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_184_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_5_17_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_17_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_17_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_17_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_17_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_17_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_17_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_17_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_185_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_5_18_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_18_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_18_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_18_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_18_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_18_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_18_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_18_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_186_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_5_19_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_19_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_19_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_19_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_19_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_19_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_19_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_19_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_187_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_5_20_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_20_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_20_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_20_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_20_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_20_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_20_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_20_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_188_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_5_21_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_21_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_21_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_21_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_21_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_21_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_21_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_21_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_189_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_5_22_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_22_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_22_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_22_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_22_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_22_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_22_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_22_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_190_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_5_23_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_23_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_23_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_23_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_23_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_23_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_23_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_23_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_191_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_5_24_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_24_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_24_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_24_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_24_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_24_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_24_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_24_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_192_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_5_25_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_25_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_25_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_25_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_25_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_25_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_25_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_25_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_193_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_5_26_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_26_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_26_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_26_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_26_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_26_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_26_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_26_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_194_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_5_27_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_27_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_27_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_27_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_27_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_27_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_27_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_27_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_195_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_5_28_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_28_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_28_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_28_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_28_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_28_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_28_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_28_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_196_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_5_29_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_29_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_29_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_29_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_29_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_29_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_29_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_29_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_197_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_5_30_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_30_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_30_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_30_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_30_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_30_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_30_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_30_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_198_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_5_31_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_31_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_31_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_31_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_31_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_31_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_5_31_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_5_31_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_199_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_6_0_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_0_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_0_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_0_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_0_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_0_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_0_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_0_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_200_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_6_1_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_1_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_1_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_1_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_1_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_1_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_1_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_1_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_201_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_6_2_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_2_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_2_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_2_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_2_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_2_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_2_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_2_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_202_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_6_3_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_3_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_3_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_3_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_3_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_3_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_3_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_3_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_203_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_6_4_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_4_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_4_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_4_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_4_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_4_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_4_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_4_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_204_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_6_5_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_5_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_5_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_5_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_5_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_5_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_5_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_5_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_205_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_6_6_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_6_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_6_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_6_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_6_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_6_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_6_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_6_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_206_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_6_7_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_7_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_7_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_7_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_7_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_7_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_7_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_7_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_207_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_6_8_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_8_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_8_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_8_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_8_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_8_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_8_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_8_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_208_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_6_9_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_9_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_9_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_9_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_9_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_9_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_9_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_9_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_209_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_6_10_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_10_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_10_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_10_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_10_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_10_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_10_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_10_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_210_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_6_11_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_11_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_11_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_11_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_11_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_11_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_11_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_11_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_211_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_6_12_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_12_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_12_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_12_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_12_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_12_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_12_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_12_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_212_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_6_13_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_13_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_13_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_13_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_13_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_13_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_13_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_13_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_213_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_6_14_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_14_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_14_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_14_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_14_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_14_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_14_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_14_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_214_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_6_15_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_15_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_15_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_15_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_15_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_15_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_15_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_15_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_215_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_6_16_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_16_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_16_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_16_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_16_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_16_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_16_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_16_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_216_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_6_17_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_17_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_17_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_17_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_17_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_17_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_17_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_17_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_217_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_6_18_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_18_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_18_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_18_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_18_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_18_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_18_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_18_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_218_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_6_19_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_19_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_19_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_19_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_19_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_19_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_19_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_19_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_219_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_6_20_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_20_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_20_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_20_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_20_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_20_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_20_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_20_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_220_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_6_21_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_21_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_21_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_21_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_21_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_21_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_21_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_21_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_221_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_6_22_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_22_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_22_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_22_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_22_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_22_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_22_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_22_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_222_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_6_23_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_23_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_23_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_23_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_23_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_23_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_23_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_23_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_223_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_6_24_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_24_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_24_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_24_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_24_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_24_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_24_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_24_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_224_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_6_25_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_25_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_25_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_25_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_25_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_25_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_25_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_25_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_225_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_6_26_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_26_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_26_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_26_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_26_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_26_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_26_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_26_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_226_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_6_27_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_27_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_27_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_27_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_27_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_27_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_27_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_27_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_227_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_6_28_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_28_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_28_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_28_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_28_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_28_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_28_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_28_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_228_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_6_29_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_29_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_29_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_29_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_29_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_29_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_29_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_29_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_229_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_6_30_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_30_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_30_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_30_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_30_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_30_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_30_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_30_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_230_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_6_31_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_31_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_31_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_31_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_31_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_31_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_6_31_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_6_31_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_231_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_7_0_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_0_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_0_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_0_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_0_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_0_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_0_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_0_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_232_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_7_1_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_1_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_1_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_1_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_1_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_1_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_1_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_1_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_233_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_7_2_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_2_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_2_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_2_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_2_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_2_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_2_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_2_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_234_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_7_3_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_3_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_3_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_3_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_3_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_3_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_3_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_3_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_235_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_7_4_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_4_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_4_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_4_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_4_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_4_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_4_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_4_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_236_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_7_5_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_5_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_5_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_5_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_5_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_5_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_5_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_5_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_237_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_7_6_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_6_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_6_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_6_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_6_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_6_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_6_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_6_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_238_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_7_7_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_7_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_7_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_7_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_7_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_7_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_7_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_7_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_239_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_7_8_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_8_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_8_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_8_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_8_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_8_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_8_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_8_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_240_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_7_9_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_9_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_9_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_9_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_9_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_9_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_9_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_9_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_241_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_7_10_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_10_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_10_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_10_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_10_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_10_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_10_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_10_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_242_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_7_11_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_11_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_11_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_11_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_11_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_11_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_11_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_11_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_243_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_7_12_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_12_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_12_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_12_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_12_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_12_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_12_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_12_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_244_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_7_13_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_13_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_13_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_13_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_13_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_13_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_13_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_13_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_245_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_7_14_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_14_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_14_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_14_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_14_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_14_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_14_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_14_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_246_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_7_15_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_15_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_15_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_15_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_15_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_15_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_15_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_15_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_247_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_7_16_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_16_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_16_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_16_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_16_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_16_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_16_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_16_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_248_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_7_17_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_17_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_17_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_17_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_17_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_17_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_17_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_17_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_249_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_7_18_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_18_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_18_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_18_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_18_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_18_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_18_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_18_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_250_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_7_19_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_19_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_19_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_19_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_19_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_19_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_19_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_19_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_251_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_7_20_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_20_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_20_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_20_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_20_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_20_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_20_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_20_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_252_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_7_21_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_21_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_21_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_21_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_21_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_21_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_21_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_21_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_253_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_7_22_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_22_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_22_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_22_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_22_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_22_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_22_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_22_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_254_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_7_23_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_23_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_23_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_23_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_23_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_23_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_23_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_23_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_255_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_7_24_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_24_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_24_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_24_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_24_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_24_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_24_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_24_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_256_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_7_25_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_25_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_25_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_25_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_25_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_25_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_25_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_25_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_257_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_7_26_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_26_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_26_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_26_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_26_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_26_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_26_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_26_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_258_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_7_27_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_27_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_27_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_27_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_27_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_27_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_27_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_27_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_259_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_7_28_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_28_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_28_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_28_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_28_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_28_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_28_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_28_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_260_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_7_29_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_29_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_29_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_29_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_29_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_29_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_29_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_29_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_261_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_7_30_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_30_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_30_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_30_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_30_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_30_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_30_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_30_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_262_4_32_16_16_32_1_gen
    PORT(
      clkr_en : OUT STD_LOGIC;
      clkw_en : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      clkr : IN STD_LOGIC;
      clkr_en_d : IN STD_LOGIC;
      clkw_en_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_7_31_i_q : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_31_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_31_i_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_31_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_31_i_d_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_31_i_q_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_7_31_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_7_31_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_263_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_0_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_0_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_0_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_0_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_264_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_1_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_1_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_1_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_1_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_1_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_1_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_265_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_2_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_2_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_2_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_2_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_2_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_2_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_266_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_3_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_3_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_3_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_3_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_3_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_3_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_267_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_4_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_4_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_4_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_4_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_4_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_4_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_268_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_5_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_5_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_5_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_5_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_5_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_5_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_269_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_6_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_6_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_6_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_6_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_6_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_6_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_270_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_7_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_7_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_7_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_7_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_7_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_7_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_271_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_8_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_8_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_8_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_8_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_8_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_8_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_272_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_9_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_9_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_9_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_9_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_9_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_9_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_273_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_10_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_10_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_10_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_10_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_10_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_10_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_274_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_11_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_11_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_11_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_11_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_11_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_11_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_275_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_12_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_12_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_12_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_12_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_12_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_12_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_276_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_13_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_13_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_13_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_13_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_13_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_13_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_277_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_14_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_14_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_14_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_14_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_14_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_14_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_278_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_15_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_15_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_15_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_15_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_15_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_15_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_279_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_16_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_16_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_16_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_16_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_16_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_16_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_280_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_17_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_17_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_17_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_17_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_17_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_17_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_281_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_18_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_18_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_18_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_18_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_18_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_18_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_282_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_19_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_19_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_19_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_19_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_19_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_19_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_283_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_20_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_20_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_20_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_20_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_20_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_20_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_284_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_21_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_21_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_21_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_21_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_21_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_21_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_285_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_22_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_22_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_22_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_22_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_22_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_22_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_286_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_23_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_23_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_23_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_23_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_23_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_23_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_287_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_24_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_24_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_24_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_24_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_24_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_24_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_288_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_25_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_25_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_25_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_25_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_25_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_25_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_289_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_26_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_26_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_26_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_26_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_26_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_26_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_290_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_27_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_27_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_27_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_27_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_27_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_27_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_291_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_28_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_28_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_28_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_28_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_28_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_28_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_292_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_29_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_29_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_29_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_29_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_29_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_29_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_293_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_30_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_30_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_30_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_30_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_30_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_30_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_294_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_31_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_31_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_31_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_31_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_31_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_31_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_295_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_1_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_0_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_0_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_0_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_0_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_296_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_1_1_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_1_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_1_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_1_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_1_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_1_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_297_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_1_2_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_2_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_2_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_2_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_2_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_2_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_298_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_1_3_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_3_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_3_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_3_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_3_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_3_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_299_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_1_4_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_4_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_4_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_4_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_4_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_4_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_300_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_1_5_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_5_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_5_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_5_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_5_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_5_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_301_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_1_6_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_6_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_6_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_6_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_6_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_6_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_302_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_1_7_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_7_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_7_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_7_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_7_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_7_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_303_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_1_8_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_8_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_8_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_8_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_8_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_8_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_304_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_1_9_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_9_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_9_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_9_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_9_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_9_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_305_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_1_10_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_10_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_10_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_10_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_10_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_10_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_306_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_1_11_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_11_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_11_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_11_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_11_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_11_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_307_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_1_12_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_12_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_12_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_12_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_12_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_12_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_308_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_1_13_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_13_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_13_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_13_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_13_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_13_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_309_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_1_14_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_14_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_14_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_14_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_14_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_14_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_310_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_1_15_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_15_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_15_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_15_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_15_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_15_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_311_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_1_16_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_16_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_16_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_16_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_16_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_16_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_312_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_1_17_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_17_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_17_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_17_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_17_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_17_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_313_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_1_18_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_18_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_18_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_18_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_18_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_18_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_314_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_1_19_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_19_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_19_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_19_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_19_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_19_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_315_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_1_20_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_20_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_20_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_20_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_20_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_20_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_316_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_1_21_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_21_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_21_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_21_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_21_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_21_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_317_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_1_22_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_22_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_22_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_22_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_22_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_22_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_318_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_1_23_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_23_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_23_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_23_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_23_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_23_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_319_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_1_24_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_24_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_24_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_24_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_24_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_24_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_320_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_1_25_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_25_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_25_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_25_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_25_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_25_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_321_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_1_26_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_26_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_26_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_26_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_26_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_26_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_322_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_1_27_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_27_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_27_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_27_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_27_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_27_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_323_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_1_28_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_28_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_28_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_28_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_28_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_28_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_324_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_1_29_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_29_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_29_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_29_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_29_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_29_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_325_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_1_30_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_30_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_30_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_30_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_30_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_30_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_326_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_1_31_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_31_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_31_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_31_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_31_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_31_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_327_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_2_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_0_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_2_0_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_2_0_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_0_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_328_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_2_1_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_1_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_1_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_2_1_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_2_1_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_1_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_329_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_2_2_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_2_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_2_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_2_2_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_2_2_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_2_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_330_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_2_3_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_3_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_3_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_2_3_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_2_3_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_3_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_331_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_2_4_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_4_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_4_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_2_4_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_2_4_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_4_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_332_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_2_5_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_5_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_5_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_2_5_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_2_5_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_5_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_333_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_2_6_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_6_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_6_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_2_6_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_2_6_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_6_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_334_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_2_7_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_7_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_7_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_2_7_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_2_7_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_7_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_335_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_2_8_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_8_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_8_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_2_8_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_2_8_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_8_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_336_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_2_9_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_9_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_9_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_2_9_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_2_9_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_9_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_337_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_2_10_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_10_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_10_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_2_10_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_2_10_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_10_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_338_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_2_11_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_11_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_11_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_2_11_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_2_11_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_11_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_339_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_2_12_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_12_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_12_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_2_12_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_2_12_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_12_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_340_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_2_13_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_13_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_13_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_2_13_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_2_13_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_13_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_341_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_2_14_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_14_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_14_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_2_14_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_2_14_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_14_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_342_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_2_15_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_15_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_15_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_2_15_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_2_15_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_15_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_343_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_2_16_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_16_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_16_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_2_16_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_2_16_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_16_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_344_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_2_17_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_17_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_17_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_2_17_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_2_17_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_17_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_345_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_2_18_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_18_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_18_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_2_18_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_2_18_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_18_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_346_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_2_19_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_19_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_19_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_2_19_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_2_19_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_19_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_347_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_2_20_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_20_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_20_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_2_20_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_2_20_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_20_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_348_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_2_21_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_21_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_21_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_2_21_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_2_21_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_21_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_349_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_2_22_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_22_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_22_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_2_22_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_2_22_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_22_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_350_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_2_23_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_23_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_23_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_2_23_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_2_23_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_23_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_351_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_2_24_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_24_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_24_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_2_24_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_2_24_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_24_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_352_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_2_25_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_25_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_25_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_2_25_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_2_25_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_25_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_353_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_2_26_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_26_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_26_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_2_26_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_2_26_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_26_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_354_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_2_27_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_27_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_27_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_2_27_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_2_27_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_27_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_355_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_2_28_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_28_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_28_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_2_28_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_2_28_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_28_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_356_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_2_29_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_29_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_29_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_2_29_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_2_29_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_29_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_357_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_2_30_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_30_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_30_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_2_30_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_2_30_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_30_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_358_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_2_31_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_31_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_31_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_2_31_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_2_31_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_2_31_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_359_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_3_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_0_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_3_0_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_3_0_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_0_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_360_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_3_1_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_1_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_1_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_3_1_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_3_1_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_1_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_361_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_3_2_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_2_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_2_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_3_2_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_3_2_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_2_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_362_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_3_3_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_3_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_3_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_3_3_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_3_3_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_3_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_363_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_3_4_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_4_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_4_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_3_4_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_3_4_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_4_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_364_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_3_5_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_5_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_5_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_3_5_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_3_5_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_5_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_365_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_3_6_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_6_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_6_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_3_6_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_3_6_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_6_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_366_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_3_7_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_7_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_7_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_3_7_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_3_7_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_7_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_367_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_3_8_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_8_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_8_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_3_8_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_3_8_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_8_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_368_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_3_9_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_9_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_9_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_3_9_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_3_9_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_9_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_369_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_3_10_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_10_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_10_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_3_10_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_3_10_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_10_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_370_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_3_11_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_11_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_11_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_3_11_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_3_11_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_11_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_371_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_3_12_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_12_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_12_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_3_12_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_3_12_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_12_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_372_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_3_13_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_13_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_13_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_3_13_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_3_13_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_13_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_373_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_3_14_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_14_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_14_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_3_14_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_3_14_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_14_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_374_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_3_15_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_15_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_15_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_3_15_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_3_15_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_15_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_375_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_3_16_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_16_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_16_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_3_16_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_3_16_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_16_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_376_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_3_17_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_17_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_17_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_3_17_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_3_17_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_17_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_377_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_3_18_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_18_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_18_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_3_18_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_3_18_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_18_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_378_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_3_19_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_19_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_19_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_3_19_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_3_19_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_19_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_379_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_3_20_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_20_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_20_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_3_20_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_3_20_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_20_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_380_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_3_21_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_21_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_21_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_3_21_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_3_21_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_21_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_381_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_3_22_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_22_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_22_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_3_22_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_3_22_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_22_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_382_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_3_23_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_23_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_23_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_3_23_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_3_23_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_23_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_383_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_3_24_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_24_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_24_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_3_24_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_3_24_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_24_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_384_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_3_25_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_25_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_25_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_3_25_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_3_25_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_25_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_385_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_3_26_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_26_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_26_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_3_26_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_3_26_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_26_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_386_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_3_27_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_27_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_27_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_3_27_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_3_27_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_27_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_387_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_3_28_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_28_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_28_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_3_28_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_3_28_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_28_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_388_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_3_29_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_29_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_29_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_3_29_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_3_29_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_29_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_389_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_3_30_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_30_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_30_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_3_30_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_3_30_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_30_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_390_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_3_31_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_31_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_31_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_3_31_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_3_31_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_3_31_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_391_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_4_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_0_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_0_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_0_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_0_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_392_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_4_1_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_1_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_1_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_1_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_1_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_1_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_393_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_4_2_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_2_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_2_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_2_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_2_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_2_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_394_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_4_3_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_3_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_3_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_3_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_3_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_3_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_395_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_4_4_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_4_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_4_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_4_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_4_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_4_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_396_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_4_5_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_5_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_5_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_5_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_5_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_5_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_397_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_4_6_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_6_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_6_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_6_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_6_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_6_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_398_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_4_7_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_7_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_7_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_7_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_7_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_7_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_399_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_4_8_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_8_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_8_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_8_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_8_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_8_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_400_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_4_9_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_9_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_9_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_9_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_9_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_9_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_401_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_4_10_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_10_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_10_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_10_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_10_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_10_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_402_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_4_11_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_11_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_11_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_11_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_11_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_11_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_403_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_4_12_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_12_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_12_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_12_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_12_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_12_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_404_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_4_13_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_13_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_13_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_13_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_13_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_13_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_405_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_4_14_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_14_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_14_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_14_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_14_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_14_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_406_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_4_15_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_15_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_15_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_15_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_15_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_15_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_407_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_4_16_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_16_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_16_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_16_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_16_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_16_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_408_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_4_17_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_17_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_17_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_17_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_17_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_17_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_409_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_4_18_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_18_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_18_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_18_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_18_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_18_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_410_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_4_19_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_19_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_19_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_19_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_19_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_19_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_411_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_4_20_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_20_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_20_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_20_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_20_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_20_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_412_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_4_21_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_21_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_21_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_21_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_21_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_21_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_413_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_4_22_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_22_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_22_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_22_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_22_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_22_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_414_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_4_23_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_23_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_23_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_23_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_23_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_23_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_415_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_4_24_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_24_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_24_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_24_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_24_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_24_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_416_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_4_25_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_25_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_25_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_25_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_25_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_25_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_417_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_4_26_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_26_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_26_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_26_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_26_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_26_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_418_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_4_27_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_27_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_27_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_27_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_27_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_27_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_419_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_4_28_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_28_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_28_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_28_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_28_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_28_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_420_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_4_29_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_29_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_29_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_29_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_29_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_29_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_421_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_4_30_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_30_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_30_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_30_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_30_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_30_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_422_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_4_31_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_31_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_31_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_31_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_4_31_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_4_31_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_423_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_5_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_0_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_5_0_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_5_0_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_0_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_424_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_5_1_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_1_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_1_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_5_1_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_5_1_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_1_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_425_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_5_2_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_2_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_2_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_5_2_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_5_2_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_2_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_426_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_5_3_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_3_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_3_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_5_3_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_5_3_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_3_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_427_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_5_4_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_4_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_4_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_5_4_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_5_4_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_4_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_428_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_5_5_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_5_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_5_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_5_5_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_5_5_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_5_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_429_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_5_6_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_6_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_6_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_5_6_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_5_6_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_6_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_430_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_5_7_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_7_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_7_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_5_7_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_5_7_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_7_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_431_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_5_8_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_8_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_8_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_5_8_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_5_8_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_8_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_432_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_5_9_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_9_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_9_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_5_9_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_5_9_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_9_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_433_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_5_10_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_10_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_10_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_5_10_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_5_10_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_10_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_434_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_5_11_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_11_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_11_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_5_11_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_5_11_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_11_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_435_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_5_12_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_12_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_12_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_5_12_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_5_12_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_12_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_436_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_5_13_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_13_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_13_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_5_13_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_5_13_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_13_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_437_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_5_14_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_14_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_14_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_5_14_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_5_14_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_14_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_438_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_5_15_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_15_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_15_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_5_15_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_5_15_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_15_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_439_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_5_16_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_16_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_16_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_5_16_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_5_16_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_16_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_440_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_5_17_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_17_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_17_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_5_17_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_5_17_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_17_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_441_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_5_18_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_18_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_18_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_5_18_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_5_18_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_18_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_442_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_5_19_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_19_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_19_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_5_19_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_5_19_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_19_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_443_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_5_20_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_20_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_20_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_5_20_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_5_20_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_20_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_444_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_5_21_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_21_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_21_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_5_21_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_5_21_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_21_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_445_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_5_22_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_22_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_22_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_5_22_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_5_22_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_22_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_446_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_5_23_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_23_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_23_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_5_23_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_5_23_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_23_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_447_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_5_24_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_24_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_24_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_5_24_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_5_24_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_24_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_448_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_5_25_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_25_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_25_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_5_25_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_5_25_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_25_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_449_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_5_26_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_26_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_26_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_5_26_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_5_26_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_26_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_450_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_5_27_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_27_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_27_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_5_27_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_5_27_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_27_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_451_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_5_28_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_28_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_28_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_5_28_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_5_28_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_28_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_452_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_5_29_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_29_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_29_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_5_29_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_5_29_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_29_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_453_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_5_30_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_30_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_30_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_5_30_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_5_30_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_30_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_454_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_5_31_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_31_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_31_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_5_31_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_5_31_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_5_31_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_455_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_6_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_0_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_6_0_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_6_0_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_0_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_456_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_6_1_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_1_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_1_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_6_1_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_6_1_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_1_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_457_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_6_2_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_2_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_2_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_6_2_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_6_2_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_2_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_458_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_6_3_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_3_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_3_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_6_3_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_6_3_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_3_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_459_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_6_4_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_4_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_4_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_6_4_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_6_4_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_4_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_460_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_6_5_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_5_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_5_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_6_5_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_6_5_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_5_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_461_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_6_6_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_6_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_6_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_6_6_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_6_6_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_6_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_462_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_6_7_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_7_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_7_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_6_7_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_6_7_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_7_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_463_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_6_8_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_8_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_8_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_6_8_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_6_8_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_8_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_464_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_6_9_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_9_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_9_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_6_9_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_6_9_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_9_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_465_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_6_10_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_10_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_10_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_6_10_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_6_10_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_10_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_466_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_6_11_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_11_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_11_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_6_11_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_6_11_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_11_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_467_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_6_12_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_12_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_12_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_6_12_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_6_12_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_12_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_468_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_6_13_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_13_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_13_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_6_13_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_6_13_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_13_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_469_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_6_14_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_14_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_14_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_6_14_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_6_14_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_14_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_470_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_6_15_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_15_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_15_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_6_15_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_6_15_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_15_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_471_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_6_16_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_16_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_16_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_6_16_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_6_16_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_16_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_472_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_6_17_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_17_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_17_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_6_17_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_6_17_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_17_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_473_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_6_18_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_18_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_18_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_6_18_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_6_18_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_18_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_474_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_6_19_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_19_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_19_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_6_19_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_6_19_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_19_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_475_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_6_20_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_20_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_20_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_6_20_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_6_20_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_20_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_476_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_6_21_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_21_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_21_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_6_21_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_6_21_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_21_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_477_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_6_22_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_22_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_22_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_6_22_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_6_22_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_22_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_478_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_6_23_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_23_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_23_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_6_23_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_6_23_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_23_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_479_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_6_24_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_24_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_24_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_6_24_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_6_24_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_24_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_480_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_6_25_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_25_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_25_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_6_25_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_6_25_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_25_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_481_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_6_26_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_26_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_26_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_6_26_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_6_26_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_26_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_482_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_6_27_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_27_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_27_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_6_27_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_6_27_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_27_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_483_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_6_28_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_28_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_28_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_6_28_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_6_28_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_28_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_484_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_6_29_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_29_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_29_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_6_29_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_6_29_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_29_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_485_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_6_30_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_30_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_30_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_6_30_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_6_30_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_30_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_486_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_6_31_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_31_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_31_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_6_31_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_6_31_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_6_31_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_487_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_7_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_0_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_7_0_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_7_0_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_0_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_488_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_7_1_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_1_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_1_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_7_1_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_7_1_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_1_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_489_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_7_2_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_2_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_2_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_7_2_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_7_2_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_2_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_490_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_7_3_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_3_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_3_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_7_3_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_7_3_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_3_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_491_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_7_4_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_4_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_4_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_7_4_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_7_4_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_4_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_492_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_7_5_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_5_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_5_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_7_5_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_7_5_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_5_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_493_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_7_6_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_6_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_6_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_7_6_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_7_6_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_6_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_494_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_7_7_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_7_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_7_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_7_7_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_7_7_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_7_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_495_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_7_8_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_8_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_8_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_7_8_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_7_8_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_8_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_496_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_7_9_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_9_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_9_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_7_9_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_7_9_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_9_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_497_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_7_10_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_10_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_10_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_7_10_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_7_10_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_10_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_498_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_7_11_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_11_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_11_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_7_11_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_7_11_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_11_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_499_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_7_12_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_12_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_12_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_7_12_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_7_12_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_12_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_500_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_7_13_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_13_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_13_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_7_13_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_7_13_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_13_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_501_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_7_14_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_14_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_14_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_7_14_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_7_14_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_14_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_502_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_7_15_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_15_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_15_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_7_15_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_7_15_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_15_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_503_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_7_16_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_16_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_16_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_7_16_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_7_16_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_16_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_504_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_7_17_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_17_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_17_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_7_17_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_7_17_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_17_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_505_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_7_18_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_18_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_18_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_7_18_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_7_18_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_18_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_506_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_7_19_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_19_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_19_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_7_19_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_7_19_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_19_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_507_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_7_20_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_20_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_20_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_7_20_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_7_20_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_20_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_508_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_7_21_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_21_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_21_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_7_21_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_7_21_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_21_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_509_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_7_22_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_22_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_22_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_7_22_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_7_22_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_22_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_510_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_7_23_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_23_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_23_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_7_23_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_7_23_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_23_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_511_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_7_24_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_24_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_24_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_7_24_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_7_24_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_24_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_512_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_7_25_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_25_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_25_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_7_25_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_7_25_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_25_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_513_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_7_26_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_26_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_26_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_7_26_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_7_26_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_26_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_514_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_7_27_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_27_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_27_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_7_27_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_7_27_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_27_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_515_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_7_28_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_28_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_28_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_7_28_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_7_28_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_28_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_516_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_7_29_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_29_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_29_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_7_29_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_7_29_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_29_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_517_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_7_30_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_30_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_30_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_7_30_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_7_30_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_30_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_518_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_7_31_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_31_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_31_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_7_31_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_7_31_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_7_31_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_519_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1
      DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_520_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_1_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1
      DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_521_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_2_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1
      DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_522_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_3_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1
      DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_523_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_4_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1
      DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_524_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_5_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1
      DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_525_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_6_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1
      DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_526_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_7_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1
      DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_527_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_8_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1
      DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_528_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_9_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1
      DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_529_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_10_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1
      DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_530_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_11_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1
      DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_531_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_12_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1
      DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_532_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_13_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1
      DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_533_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_14_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1
      DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_534_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_15_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1
      DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_535_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL twiddle_h_rsc_0_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_536_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL twiddle_h_rsc_0_1_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_537_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL twiddle_h_rsc_0_2_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_538_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL twiddle_h_rsc_0_3_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_539_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL twiddle_h_rsc_0_4_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_540_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL twiddle_h_rsc_0_5_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_541_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL twiddle_h_rsc_0_6_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_542_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL twiddle_h_rsc_0_7_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_543_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL twiddle_h_rsc_0_8_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_8_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_8_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_8_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_8_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_8_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_8_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_8_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_8_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_8_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_8_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_544_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL twiddle_h_rsc_0_9_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_9_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_9_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_9_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_9_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_9_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_9_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_9_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_9_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_9_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_9_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_545_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL twiddle_h_rsc_0_10_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_10_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_10_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_10_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_10_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_10_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_10_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_10_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_10_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_10_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_10_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_546_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL twiddle_h_rsc_0_11_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_11_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_11_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_11_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_11_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_11_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_11_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_11_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_11_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_11_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_11_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_547_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL twiddle_h_rsc_0_12_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_12_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_12_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_12_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_12_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_12_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_12_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_12_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_12_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_12_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_12_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_548_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL twiddle_h_rsc_0_13_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_13_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_13_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_13_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_13_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_13_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_13_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_13_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_13_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_13_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_13_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_549_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL twiddle_h_rsc_0_14_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_14_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_14_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_14_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_14_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_14_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_14_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_14_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_14_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_14_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_14_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_550_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL twiddle_h_rsc_0_15_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_15_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_15_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_15_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_15_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_15_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_15_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_15_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_15_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_15_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_15_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);

  COMPONENT peaseNTT_core
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_triosy_0_0_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_1_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_2_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_3_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_4_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_5_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_6_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_7_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_8_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_9_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_10_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_11_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_12_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_13_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_14_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_15_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_16_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_17_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_18_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_19_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_20_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_21_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_22_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_23_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_24_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_25_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_26_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_27_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_28_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_29_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_30_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_31_lz : OUT STD_LOGIC;
      xt_rsc_triosy_1_0_lz : OUT STD_LOGIC;
      xt_rsc_triosy_1_1_lz : OUT STD_LOGIC;
      xt_rsc_triosy_1_2_lz : OUT STD_LOGIC;
      xt_rsc_triosy_1_3_lz : OUT STD_LOGIC;
      xt_rsc_triosy_1_4_lz : OUT STD_LOGIC;
      xt_rsc_triosy_1_5_lz : OUT STD_LOGIC;
      xt_rsc_triosy_1_6_lz : OUT STD_LOGIC;
      xt_rsc_triosy_1_7_lz : OUT STD_LOGIC;
      xt_rsc_triosy_1_8_lz : OUT STD_LOGIC;
      xt_rsc_triosy_1_9_lz : OUT STD_LOGIC;
      xt_rsc_triosy_1_10_lz : OUT STD_LOGIC;
      xt_rsc_triosy_1_11_lz : OUT STD_LOGIC;
      xt_rsc_triosy_1_12_lz : OUT STD_LOGIC;
      xt_rsc_triosy_1_13_lz : OUT STD_LOGIC;
      xt_rsc_triosy_1_14_lz : OUT STD_LOGIC;
      xt_rsc_triosy_1_15_lz : OUT STD_LOGIC;
      xt_rsc_triosy_1_16_lz : OUT STD_LOGIC;
      xt_rsc_triosy_1_17_lz : OUT STD_LOGIC;
      xt_rsc_triosy_1_18_lz : OUT STD_LOGIC;
      xt_rsc_triosy_1_19_lz : OUT STD_LOGIC;
      xt_rsc_triosy_1_20_lz : OUT STD_LOGIC;
      xt_rsc_triosy_1_21_lz : OUT STD_LOGIC;
      xt_rsc_triosy_1_22_lz : OUT STD_LOGIC;
      xt_rsc_triosy_1_23_lz : OUT STD_LOGIC;
      xt_rsc_triosy_1_24_lz : OUT STD_LOGIC;
      xt_rsc_triosy_1_25_lz : OUT STD_LOGIC;
      xt_rsc_triosy_1_26_lz : OUT STD_LOGIC;
      xt_rsc_triosy_1_27_lz : OUT STD_LOGIC;
      xt_rsc_triosy_1_28_lz : OUT STD_LOGIC;
      xt_rsc_triosy_1_29_lz : OUT STD_LOGIC;
      xt_rsc_triosy_1_30_lz : OUT STD_LOGIC;
      xt_rsc_triosy_1_31_lz : OUT STD_LOGIC;
      xt_rsc_triosy_2_0_lz : OUT STD_LOGIC;
      xt_rsc_triosy_2_1_lz : OUT STD_LOGIC;
      xt_rsc_triosy_2_2_lz : OUT STD_LOGIC;
      xt_rsc_triosy_2_3_lz : OUT STD_LOGIC;
      xt_rsc_triosy_2_4_lz : OUT STD_LOGIC;
      xt_rsc_triosy_2_5_lz : OUT STD_LOGIC;
      xt_rsc_triosy_2_6_lz : OUT STD_LOGIC;
      xt_rsc_triosy_2_7_lz : OUT STD_LOGIC;
      xt_rsc_triosy_2_8_lz : OUT STD_LOGIC;
      xt_rsc_triosy_2_9_lz : OUT STD_LOGIC;
      xt_rsc_triosy_2_10_lz : OUT STD_LOGIC;
      xt_rsc_triosy_2_11_lz : OUT STD_LOGIC;
      xt_rsc_triosy_2_12_lz : OUT STD_LOGIC;
      xt_rsc_triosy_2_13_lz : OUT STD_LOGIC;
      xt_rsc_triosy_2_14_lz : OUT STD_LOGIC;
      xt_rsc_triosy_2_15_lz : OUT STD_LOGIC;
      xt_rsc_triosy_2_16_lz : OUT STD_LOGIC;
      xt_rsc_triosy_2_17_lz : OUT STD_LOGIC;
      xt_rsc_triosy_2_18_lz : OUT STD_LOGIC;
      xt_rsc_triosy_2_19_lz : OUT STD_LOGIC;
      xt_rsc_triosy_2_20_lz : OUT STD_LOGIC;
      xt_rsc_triosy_2_21_lz : OUT STD_LOGIC;
      xt_rsc_triosy_2_22_lz : OUT STD_LOGIC;
      xt_rsc_triosy_2_23_lz : OUT STD_LOGIC;
      xt_rsc_triosy_2_24_lz : OUT STD_LOGIC;
      xt_rsc_triosy_2_25_lz : OUT STD_LOGIC;
      xt_rsc_triosy_2_26_lz : OUT STD_LOGIC;
      xt_rsc_triosy_2_27_lz : OUT STD_LOGIC;
      xt_rsc_triosy_2_28_lz : OUT STD_LOGIC;
      xt_rsc_triosy_2_29_lz : OUT STD_LOGIC;
      xt_rsc_triosy_2_30_lz : OUT STD_LOGIC;
      xt_rsc_triosy_2_31_lz : OUT STD_LOGIC;
      xt_rsc_triosy_3_0_lz : OUT STD_LOGIC;
      xt_rsc_triosy_3_1_lz : OUT STD_LOGIC;
      xt_rsc_triosy_3_2_lz : OUT STD_LOGIC;
      xt_rsc_triosy_3_3_lz : OUT STD_LOGIC;
      xt_rsc_triosy_3_4_lz : OUT STD_LOGIC;
      xt_rsc_triosy_3_5_lz : OUT STD_LOGIC;
      xt_rsc_triosy_3_6_lz : OUT STD_LOGIC;
      xt_rsc_triosy_3_7_lz : OUT STD_LOGIC;
      xt_rsc_triosy_3_8_lz : OUT STD_LOGIC;
      xt_rsc_triosy_3_9_lz : OUT STD_LOGIC;
      xt_rsc_triosy_3_10_lz : OUT STD_LOGIC;
      xt_rsc_triosy_3_11_lz : OUT STD_LOGIC;
      xt_rsc_triosy_3_12_lz : OUT STD_LOGIC;
      xt_rsc_triosy_3_13_lz : OUT STD_LOGIC;
      xt_rsc_triosy_3_14_lz : OUT STD_LOGIC;
      xt_rsc_triosy_3_15_lz : OUT STD_LOGIC;
      xt_rsc_triosy_3_16_lz : OUT STD_LOGIC;
      xt_rsc_triosy_3_17_lz : OUT STD_LOGIC;
      xt_rsc_triosy_3_18_lz : OUT STD_LOGIC;
      xt_rsc_triosy_3_19_lz : OUT STD_LOGIC;
      xt_rsc_triosy_3_20_lz : OUT STD_LOGIC;
      xt_rsc_triosy_3_21_lz : OUT STD_LOGIC;
      xt_rsc_triosy_3_22_lz : OUT STD_LOGIC;
      xt_rsc_triosy_3_23_lz : OUT STD_LOGIC;
      xt_rsc_triosy_3_24_lz : OUT STD_LOGIC;
      xt_rsc_triosy_3_25_lz : OUT STD_LOGIC;
      xt_rsc_triosy_3_26_lz : OUT STD_LOGIC;
      xt_rsc_triosy_3_27_lz : OUT STD_LOGIC;
      xt_rsc_triosy_3_28_lz : OUT STD_LOGIC;
      xt_rsc_triosy_3_29_lz : OUT STD_LOGIC;
      xt_rsc_triosy_3_30_lz : OUT STD_LOGIC;
      xt_rsc_triosy_3_31_lz : OUT STD_LOGIC;
      xt_rsc_triosy_4_0_lz : OUT STD_LOGIC;
      xt_rsc_triosy_4_1_lz : OUT STD_LOGIC;
      xt_rsc_triosy_4_2_lz : OUT STD_LOGIC;
      xt_rsc_triosy_4_3_lz : OUT STD_LOGIC;
      xt_rsc_triosy_4_4_lz : OUT STD_LOGIC;
      xt_rsc_triosy_4_5_lz : OUT STD_LOGIC;
      xt_rsc_triosy_4_6_lz : OUT STD_LOGIC;
      xt_rsc_triosy_4_7_lz : OUT STD_LOGIC;
      xt_rsc_triosy_4_8_lz : OUT STD_LOGIC;
      xt_rsc_triosy_4_9_lz : OUT STD_LOGIC;
      xt_rsc_triosy_4_10_lz : OUT STD_LOGIC;
      xt_rsc_triosy_4_11_lz : OUT STD_LOGIC;
      xt_rsc_triosy_4_12_lz : OUT STD_LOGIC;
      xt_rsc_triosy_4_13_lz : OUT STD_LOGIC;
      xt_rsc_triosy_4_14_lz : OUT STD_LOGIC;
      xt_rsc_triosy_4_15_lz : OUT STD_LOGIC;
      xt_rsc_triosy_4_16_lz : OUT STD_LOGIC;
      xt_rsc_triosy_4_17_lz : OUT STD_LOGIC;
      xt_rsc_triosy_4_18_lz : OUT STD_LOGIC;
      xt_rsc_triosy_4_19_lz : OUT STD_LOGIC;
      xt_rsc_triosy_4_20_lz : OUT STD_LOGIC;
      xt_rsc_triosy_4_21_lz : OUT STD_LOGIC;
      xt_rsc_triosy_4_22_lz : OUT STD_LOGIC;
      xt_rsc_triosy_4_23_lz : OUT STD_LOGIC;
      xt_rsc_triosy_4_24_lz : OUT STD_LOGIC;
      xt_rsc_triosy_4_25_lz : OUT STD_LOGIC;
      xt_rsc_triosy_4_26_lz : OUT STD_LOGIC;
      xt_rsc_triosy_4_27_lz : OUT STD_LOGIC;
      xt_rsc_triosy_4_28_lz : OUT STD_LOGIC;
      xt_rsc_triosy_4_29_lz : OUT STD_LOGIC;
      xt_rsc_triosy_4_30_lz : OUT STD_LOGIC;
      xt_rsc_triosy_4_31_lz : OUT STD_LOGIC;
      xt_rsc_triosy_5_0_lz : OUT STD_LOGIC;
      xt_rsc_triosy_5_1_lz : OUT STD_LOGIC;
      xt_rsc_triosy_5_2_lz : OUT STD_LOGIC;
      xt_rsc_triosy_5_3_lz : OUT STD_LOGIC;
      xt_rsc_triosy_5_4_lz : OUT STD_LOGIC;
      xt_rsc_triosy_5_5_lz : OUT STD_LOGIC;
      xt_rsc_triosy_5_6_lz : OUT STD_LOGIC;
      xt_rsc_triosy_5_7_lz : OUT STD_LOGIC;
      xt_rsc_triosy_5_8_lz : OUT STD_LOGIC;
      xt_rsc_triosy_5_9_lz : OUT STD_LOGIC;
      xt_rsc_triosy_5_10_lz : OUT STD_LOGIC;
      xt_rsc_triosy_5_11_lz : OUT STD_LOGIC;
      xt_rsc_triosy_5_12_lz : OUT STD_LOGIC;
      xt_rsc_triosy_5_13_lz : OUT STD_LOGIC;
      xt_rsc_triosy_5_14_lz : OUT STD_LOGIC;
      xt_rsc_triosy_5_15_lz : OUT STD_LOGIC;
      xt_rsc_triosy_5_16_lz : OUT STD_LOGIC;
      xt_rsc_triosy_5_17_lz : OUT STD_LOGIC;
      xt_rsc_triosy_5_18_lz : OUT STD_LOGIC;
      xt_rsc_triosy_5_19_lz : OUT STD_LOGIC;
      xt_rsc_triosy_5_20_lz : OUT STD_LOGIC;
      xt_rsc_triosy_5_21_lz : OUT STD_LOGIC;
      xt_rsc_triosy_5_22_lz : OUT STD_LOGIC;
      xt_rsc_triosy_5_23_lz : OUT STD_LOGIC;
      xt_rsc_triosy_5_24_lz : OUT STD_LOGIC;
      xt_rsc_triosy_5_25_lz : OUT STD_LOGIC;
      xt_rsc_triosy_5_26_lz : OUT STD_LOGIC;
      xt_rsc_triosy_5_27_lz : OUT STD_LOGIC;
      xt_rsc_triosy_5_28_lz : OUT STD_LOGIC;
      xt_rsc_triosy_5_29_lz : OUT STD_LOGIC;
      xt_rsc_triosy_5_30_lz : OUT STD_LOGIC;
      xt_rsc_triosy_5_31_lz : OUT STD_LOGIC;
      xt_rsc_triosy_6_0_lz : OUT STD_LOGIC;
      xt_rsc_triosy_6_1_lz : OUT STD_LOGIC;
      xt_rsc_triosy_6_2_lz : OUT STD_LOGIC;
      xt_rsc_triosy_6_3_lz : OUT STD_LOGIC;
      xt_rsc_triosy_6_4_lz : OUT STD_LOGIC;
      xt_rsc_triosy_6_5_lz : OUT STD_LOGIC;
      xt_rsc_triosy_6_6_lz : OUT STD_LOGIC;
      xt_rsc_triosy_6_7_lz : OUT STD_LOGIC;
      xt_rsc_triosy_6_8_lz : OUT STD_LOGIC;
      xt_rsc_triosy_6_9_lz : OUT STD_LOGIC;
      xt_rsc_triosy_6_10_lz : OUT STD_LOGIC;
      xt_rsc_triosy_6_11_lz : OUT STD_LOGIC;
      xt_rsc_triosy_6_12_lz : OUT STD_LOGIC;
      xt_rsc_triosy_6_13_lz : OUT STD_LOGIC;
      xt_rsc_triosy_6_14_lz : OUT STD_LOGIC;
      xt_rsc_triosy_6_15_lz : OUT STD_LOGIC;
      xt_rsc_triosy_6_16_lz : OUT STD_LOGIC;
      xt_rsc_triosy_6_17_lz : OUT STD_LOGIC;
      xt_rsc_triosy_6_18_lz : OUT STD_LOGIC;
      xt_rsc_triosy_6_19_lz : OUT STD_LOGIC;
      xt_rsc_triosy_6_20_lz : OUT STD_LOGIC;
      xt_rsc_triosy_6_21_lz : OUT STD_LOGIC;
      xt_rsc_triosy_6_22_lz : OUT STD_LOGIC;
      xt_rsc_triosy_6_23_lz : OUT STD_LOGIC;
      xt_rsc_triosy_6_24_lz : OUT STD_LOGIC;
      xt_rsc_triosy_6_25_lz : OUT STD_LOGIC;
      xt_rsc_triosy_6_26_lz : OUT STD_LOGIC;
      xt_rsc_triosy_6_27_lz : OUT STD_LOGIC;
      xt_rsc_triosy_6_28_lz : OUT STD_LOGIC;
      xt_rsc_triosy_6_29_lz : OUT STD_LOGIC;
      xt_rsc_triosy_6_30_lz : OUT STD_LOGIC;
      xt_rsc_triosy_6_31_lz : OUT STD_LOGIC;
      xt_rsc_triosy_7_0_lz : OUT STD_LOGIC;
      xt_rsc_triosy_7_1_lz : OUT STD_LOGIC;
      xt_rsc_triosy_7_2_lz : OUT STD_LOGIC;
      xt_rsc_triosy_7_3_lz : OUT STD_LOGIC;
      xt_rsc_triosy_7_4_lz : OUT STD_LOGIC;
      xt_rsc_triosy_7_5_lz : OUT STD_LOGIC;
      xt_rsc_triosy_7_6_lz : OUT STD_LOGIC;
      xt_rsc_triosy_7_7_lz : OUT STD_LOGIC;
      xt_rsc_triosy_7_8_lz : OUT STD_LOGIC;
      xt_rsc_triosy_7_9_lz : OUT STD_LOGIC;
      xt_rsc_triosy_7_10_lz : OUT STD_LOGIC;
      xt_rsc_triosy_7_11_lz : OUT STD_LOGIC;
      xt_rsc_triosy_7_12_lz : OUT STD_LOGIC;
      xt_rsc_triosy_7_13_lz : OUT STD_LOGIC;
      xt_rsc_triosy_7_14_lz : OUT STD_LOGIC;
      xt_rsc_triosy_7_15_lz : OUT STD_LOGIC;
      xt_rsc_triosy_7_16_lz : OUT STD_LOGIC;
      xt_rsc_triosy_7_17_lz : OUT STD_LOGIC;
      xt_rsc_triosy_7_18_lz : OUT STD_LOGIC;
      xt_rsc_triosy_7_19_lz : OUT STD_LOGIC;
      xt_rsc_triosy_7_20_lz : OUT STD_LOGIC;
      xt_rsc_triosy_7_21_lz : OUT STD_LOGIC;
      xt_rsc_triosy_7_22_lz : OUT STD_LOGIC;
      xt_rsc_triosy_7_23_lz : OUT STD_LOGIC;
      xt_rsc_triosy_7_24_lz : OUT STD_LOGIC;
      xt_rsc_triosy_7_25_lz : OUT STD_LOGIC;
      xt_rsc_triosy_7_26_lz : OUT STD_LOGIC;
      xt_rsc_triosy_7_27_lz : OUT STD_LOGIC;
      xt_rsc_triosy_7_28_lz : OUT STD_LOGIC;
      xt_rsc_triosy_7_29_lz : OUT STD_LOGIC;
      xt_rsc_triosy_7_30_lz : OUT STD_LOGIC;
      xt_rsc_triosy_7_31_lz : OUT STD_LOGIC;
      p_rsc_dat : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      p_rsc_triosy_lz : OUT STD_LOGIC;
      r_rsc_triosy_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_0_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_1_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_2_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_3_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_4_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_5_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_6_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_7_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_8_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_9_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_10_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_11_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_12_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_13_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_14_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_15_lz : OUT STD_LOGIC;
      twiddle_h_rsc_triosy_0_0_lz : OUT STD_LOGIC;
      twiddle_h_rsc_triosy_0_1_lz : OUT STD_LOGIC;
      twiddle_h_rsc_triosy_0_2_lz : OUT STD_LOGIC;
      twiddle_h_rsc_triosy_0_3_lz : OUT STD_LOGIC;
      twiddle_h_rsc_triosy_0_4_lz : OUT STD_LOGIC;
      twiddle_h_rsc_triosy_0_5_lz : OUT STD_LOGIC;
      twiddle_h_rsc_triosy_0_6_lz : OUT STD_LOGIC;
      twiddle_h_rsc_triosy_0_7_lz : OUT STD_LOGIC;
      twiddle_h_rsc_triosy_0_8_lz : OUT STD_LOGIC;
      twiddle_h_rsc_triosy_0_9_lz : OUT STD_LOGIC;
      twiddle_h_rsc_triosy_0_10_lz : OUT STD_LOGIC;
      twiddle_h_rsc_triosy_0_11_lz : OUT STD_LOGIC;
      twiddle_h_rsc_triosy_0_12_lz : OUT STD_LOGIC;
      twiddle_h_rsc_triosy_0_13_lz : OUT STD_LOGIC;
      twiddle_h_rsc_triosy_0_14_lz : OUT STD_LOGIC;
      twiddle_h_rsc_triosy_0_15_lz : OUT STD_LOGIC;
      yt_rsc_0_0_i_clkr_en_d : OUT STD_LOGIC;
      yt_rsc_0_0_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_1_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_2_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_3_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_4_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_5_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_6_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_7_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_8_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_9_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_10_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_11_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_12_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_13_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_14_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_15_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_16_i_clkr_en_d : OUT STD_LOGIC;
      yt_rsc_0_16_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_17_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_18_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_19_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_20_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_21_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_22_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_23_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_24_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_25_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_26_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_27_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_28_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_29_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_30_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_31_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_0_i_clkr_en_d : OUT STD_LOGIC;
      yt_rsc_1_0_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_1_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_2_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_3_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_4_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_5_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_6_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_7_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_8_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_9_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_10_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_11_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_12_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_13_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_14_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_15_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_16_i_clkr_en_d : OUT STD_LOGIC;
      yt_rsc_1_16_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_17_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_18_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_19_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_20_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_21_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_22_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_23_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_24_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_25_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_26_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_27_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_28_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_29_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_30_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_31_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_2_0_i_clkr_en_d : OUT STD_LOGIC;
      yt_rsc_2_0_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_2_1_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_2_2_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_2_3_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_2_4_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_2_5_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_2_6_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_2_7_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_2_8_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_2_9_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_2_10_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_2_11_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_2_12_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_2_13_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_2_14_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_2_15_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_2_16_i_clkr_en_d : OUT STD_LOGIC;
      yt_rsc_2_16_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_2_17_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_2_18_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_2_19_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_2_20_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_2_21_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_2_22_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_2_23_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_2_24_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_2_25_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_2_26_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_2_27_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_2_28_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_2_29_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_2_30_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_2_31_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_3_0_i_clkr_en_d : OUT STD_LOGIC;
      yt_rsc_3_0_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_3_1_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_3_2_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_3_3_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_3_4_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_3_5_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_3_6_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_3_7_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_3_8_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_3_9_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_3_10_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_3_11_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_3_12_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_3_13_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_3_14_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_3_15_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_3_16_i_clkr_en_d : OUT STD_LOGIC;
      yt_rsc_3_16_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_3_17_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_3_18_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_3_19_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_3_20_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_3_21_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_3_22_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_3_23_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_3_24_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_3_25_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_3_26_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_3_27_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_3_28_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_3_29_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_3_30_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_3_31_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_4_0_i_clkr_en_d : OUT STD_LOGIC;
      yt_rsc_4_0_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_4_1_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_4_2_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_4_3_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_4_4_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_4_5_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_4_6_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_4_7_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_4_8_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_4_9_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_4_10_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_4_11_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_4_12_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_4_13_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_4_14_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_4_15_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_4_16_i_clkr_en_d : OUT STD_LOGIC;
      yt_rsc_4_16_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_4_17_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_4_18_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_4_19_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_4_20_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_4_21_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_4_22_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_4_23_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_4_24_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_4_25_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_4_26_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_4_27_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_4_28_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_4_29_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_4_30_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_4_31_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_5_0_i_clkr_en_d : OUT STD_LOGIC;
      yt_rsc_5_0_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_5_1_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_5_2_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_5_3_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_5_4_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_5_5_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_5_6_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_5_7_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_5_8_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_5_9_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_5_10_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_5_11_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_5_12_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_5_13_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_5_14_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_5_15_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_5_16_i_clkr_en_d : OUT STD_LOGIC;
      yt_rsc_5_16_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_5_17_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_5_18_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_5_19_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_5_20_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_5_21_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_5_22_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_5_23_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_5_24_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_5_25_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_5_26_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_5_27_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_5_28_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_5_29_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_5_30_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_5_31_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_6_0_i_clkr_en_d : OUT STD_LOGIC;
      yt_rsc_6_0_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_6_1_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_6_2_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_6_3_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_6_4_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_6_5_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_6_6_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_6_7_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_6_8_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_6_9_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_6_10_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_6_11_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_6_12_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_6_13_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_6_14_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_6_15_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_6_16_i_clkr_en_d : OUT STD_LOGIC;
      yt_rsc_6_16_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_6_17_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_6_18_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_6_19_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_6_20_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_6_21_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_6_22_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_6_23_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_6_24_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_6_25_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_6_26_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_6_27_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_6_28_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_6_29_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_6_30_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_6_31_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_7_0_i_clkr_en_d : OUT STD_LOGIC;
      yt_rsc_7_0_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_7_1_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_7_2_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_7_3_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_7_4_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_7_5_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_7_6_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_7_7_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_7_8_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_7_9_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_7_10_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_7_11_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_7_12_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_7_13_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_7_14_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_7_15_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_7_16_i_clkr_en_d : OUT STD_LOGIC;
      yt_rsc_7_16_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_7_17_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_7_18_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_7_19_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_7_20_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_7_21_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_7_22_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_7_23_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_7_24_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_7_25_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_7_26_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_7_27_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_7_28_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_7_29_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_7_30_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_7_31_i_q_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_0_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_1_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_2_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_3_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_4_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_5_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_6_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_7_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_8_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_9_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_10_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_11_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_12_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_13_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_14_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_15_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_16_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_17_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_18_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_19_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_20_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_21_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_22_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_23_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_24_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_25_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_26_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_27_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_28_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_29_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_30_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_31_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_0_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_1_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_2_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_3_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_4_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_5_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_6_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_7_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_8_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_9_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_10_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_11_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_12_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_13_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_14_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_15_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_16_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_17_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_18_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_19_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_20_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_21_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_22_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_23_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_24_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_25_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_26_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_27_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_28_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_29_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_30_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_31_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_2_0_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_2_1_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_2_2_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_2_3_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_2_4_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_2_5_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_2_6_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_2_7_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_2_8_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_2_9_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_2_10_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_2_11_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_2_12_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_2_13_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_2_14_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_2_15_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_2_16_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_2_17_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_2_18_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_2_19_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_2_20_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_2_21_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_2_22_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_2_23_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_2_24_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_2_25_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_2_26_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_2_27_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_2_28_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_2_29_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_2_30_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_2_31_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_3_0_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_3_1_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_3_2_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_3_3_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_3_4_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_3_5_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_3_6_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_3_7_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_3_8_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_3_9_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_3_10_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_3_11_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_3_12_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_3_13_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_3_14_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_3_15_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_3_16_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_3_17_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_3_18_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_3_19_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_3_20_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_3_21_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_3_22_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_3_23_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_3_24_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_3_25_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_3_26_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_3_27_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_3_28_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_3_29_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_3_30_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_3_31_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_4_0_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_4_1_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_4_2_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_4_3_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_4_4_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_4_5_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_4_6_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_4_7_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_4_8_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_4_9_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_4_10_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_4_11_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_4_12_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_4_13_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_4_14_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_4_15_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_4_16_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_4_17_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_4_18_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_4_19_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_4_20_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_4_21_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_4_22_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_4_23_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_4_24_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_4_25_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_4_26_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_4_27_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_4_28_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_4_29_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_4_30_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_4_31_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_5_0_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_5_1_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_5_2_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_5_3_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_5_4_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_5_5_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_5_6_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_5_7_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_5_8_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_5_9_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_5_10_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_5_11_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_5_12_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_5_13_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_5_14_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_5_15_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_5_16_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_5_17_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_5_18_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_5_19_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_5_20_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_5_21_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_5_22_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_5_23_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_5_24_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_5_25_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_5_26_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_5_27_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_5_28_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_5_29_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_5_30_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_5_31_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_6_0_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_6_1_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_6_2_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_6_3_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_6_4_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_6_5_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_6_6_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_6_7_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_6_8_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_6_9_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_6_10_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_6_11_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_6_12_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_6_13_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_6_14_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_6_15_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_6_16_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_6_17_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_6_18_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_6_19_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_6_20_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_6_21_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_6_22_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_6_23_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_6_24_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_6_25_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_6_26_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_6_27_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_6_28_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_6_29_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_6_30_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_6_31_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_7_0_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_7_1_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_7_2_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_7_3_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_7_4_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_7_5_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_7_6_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_7_7_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_7_8_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_7_9_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_7_10_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_7_11_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_7_12_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_7_13_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_7_14_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_7_15_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_7_16_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_7_17_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_7_18_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_7_19_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_7_20_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_7_21_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_7_22_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_7_23_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_7_24_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_7_25_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_7_26_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_7_27_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_7_28_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_7_29_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_7_30_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_7_31_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_0_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
          DOWNTO 0);
      twiddle_rsc_0_1_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_1_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
          DOWNTO 0);
      twiddle_rsc_0_2_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_2_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
          DOWNTO 0);
      twiddle_rsc_0_3_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_3_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
          DOWNTO 0);
      twiddle_rsc_0_4_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_4_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
          DOWNTO 0);
      twiddle_rsc_0_5_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_5_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
          DOWNTO 0);
      twiddle_rsc_0_6_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_6_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
          DOWNTO 0);
      twiddle_rsc_0_7_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_7_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
          DOWNTO 0);
      twiddle_rsc_0_8_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_8_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
          DOWNTO 0);
      twiddle_rsc_0_9_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_9_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
          DOWNTO 0);
      twiddle_rsc_0_10_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_10_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      twiddle_rsc_0_11_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_11_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      twiddle_rsc_0_12_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_12_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      twiddle_rsc_0_13_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_13_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      twiddle_rsc_0_14_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_14_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      twiddle_rsc_0_15_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_15_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      twiddle_h_rsc_0_0_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_h_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      twiddle_h_rsc_0_1_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_1_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_h_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      twiddle_h_rsc_0_2_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_2_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_h_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      twiddle_h_rsc_0_3_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_3_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_h_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      twiddle_h_rsc_0_4_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_4_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_h_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      twiddle_h_rsc_0_5_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_5_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_h_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      twiddle_h_rsc_0_6_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_6_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_h_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      twiddle_h_rsc_0_7_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_7_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_h_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      twiddle_h_rsc_0_8_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_8_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_h_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      twiddle_h_rsc_0_9_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_9_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_h_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      twiddle_h_rsc_0_10_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_10_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_h_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      twiddle_h_rsc_0_11_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_11_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_h_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      twiddle_h_rsc_0_12_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_12_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_h_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      twiddle_h_rsc_0_13_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_13_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_h_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      twiddle_h_rsc_0_14_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_14_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_h_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      twiddle_h_rsc_0_15_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_15_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_h_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      yt_rsc_0_0_i_d_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_0_i_radr_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      yt_rsc_0_0_i_wadr_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      yt_rsc_0_0_i_we_d_pff : OUT STD_LOGIC;
      yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_pff : OUT STD_LOGIC;
      yt_rsc_0_1_i_d_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_1_i_wadr_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      yt_rsc_0_2_i_d_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_2_i_wadr_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      yt_rsc_0_3_i_d_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_3_i_wadr_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      yt_rsc_0_4_i_d_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_4_i_wadr_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      yt_rsc_0_5_i_d_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_5_i_wadr_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      yt_rsc_0_6_i_d_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_6_i_wadr_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      yt_rsc_0_7_i_d_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_8_i_d_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_9_i_d_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_10_i_d_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_10_i_wadr_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      yt_rsc_0_11_i_d_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_11_i_wadr_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      yt_rsc_0_12_i_d_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_13_i_d_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_14_i_d_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_15_i_d_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_16_i_we_d_pff : OUT STD_LOGIC;
      yt_rsc_1_0_i_we_d_pff : OUT STD_LOGIC;
      yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_pff : OUT STD_LOGIC;
      yt_rsc_1_16_i_we_d_pff : OUT STD_LOGIC;
      yt_rsc_2_0_i_we_d_pff : OUT STD_LOGIC;
      yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_pff : OUT STD_LOGIC;
      yt_rsc_2_16_i_we_d_pff : OUT STD_LOGIC;
      yt_rsc_3_0_i_we_d_pff : OUT STD_LOGIC;
      yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_pff : OUT STD_LOGIC;
      yt_rsc_3_16_i_we_d_pff : OUT STD_LOGIC;
      yt_rsc_4_0_i_d_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_4_0_i_wadr_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      yt_rsc_4_0_i_we_d_pff : OUT STD_LOGIC;
      yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_pff : OUT STD_LOGIC;
      yt_rsc_4_1_i_d_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_4_1_i_wadr_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      yt_rsc_4_2_i_d_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_4_2_i_wadr_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      yt_rsc_4_3_i_d_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_4_3_i_wadr_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      yt_rsc_4_4_i_d_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_4_4_i_wadr_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      yt_rsc_4_5_i_d_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_4_5_i_wadr_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      yt_rsc_4_6_i_d_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_4_6_i_wadr_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      yt_rsc_4_7_i_d_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_4_8_i_d_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_4_9_i_d_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_4_9_i_wadr_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      yt_rsc_4_10_i_d_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_4_10_i_wadr_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      yt_rsc_4_11_i_d_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_4_11_i_wadr_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      yt_rsc_4_12_i_d_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_4_13_i_d_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_4_14_i_d_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_4_15_i_d_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_4_16_i_we_d_pff : OUT STD_LOGIC;
      yt_rsc_5_0_i_we_d_pff : OUT STD_LOGIC;
      yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_pff : OUT STD_LOGIC;
      yt_rsc_5_16_i_we_d_pff : OUT STD_LOGIC;
      yt_rsc_6_0_i_we_d_pff : OUT STD_LOGIC;
      yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_pff : OUT STD_LOGIC;
      yt_rsc_6_16_i_we_d_pff : OUT STD_LOGIC;
      yt_rsc_7_0_i_we_d_pff : OUT STD_LOGIC;
      yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_pff : OUT STD_LOGIC;
      yt_rsc_7_16_i_we_d_pff : OUT STD_LOGIC;
      xt_rsc_0_0_i_adra_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      xt_rsc_0_0_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_0_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff : OUT STD_LOGIC;
      xt_rsc_0_1_i_adra_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      xt_rsc_0_1_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_2_i_adra_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      xt_rsc_0_2_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_3_i_adra_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      xt_rsc_0_3_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_4_i_adra_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      xt_rsc_0_4_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_5_i_adra_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      xt_rsc_0_5_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_6_i_adra_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      xt_rsc_0_6_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_7_i_adra_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      xt_rsc_0_7_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_8_i_adra_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      xt_rsc_0_8_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_9_i_adra_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      xt_rsc_0_9_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_10_i_adra_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      xt_rsc_0_10_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_11_i_adra_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      xt_rsc_0_11_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_12_i_adra_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      xt_rsc_0_12_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_13_i_adra_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      xt_rsc_0_13_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_14_i_adra_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      xt_rsc_0_14_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_15_i_adra_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      xt_rsc_0_15_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_16_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_1_0_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff : OUT STD_LOGIC;
      xt_rsc_1_16_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_2_0_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff : OUT STD_LOGIC;
      xt_rsc_2_16_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_3_0_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff : OUT STD_LOGIC;
      xt_rsc_3_16_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_4_0_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff : OUT STD_LOGIC;
      xt_rsc_4_1_i_adra_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      xt_rsc_4_1_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_4_2_i_adra_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      xt_rsc_4_2_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_4_3_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_4_4_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_4_5_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_4_6_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_4_7_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_4_8_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_4_9_i_adra_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      xt_rsc_4_9_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_4_10_i_adra_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      xt_rsc_4_10_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_4_11_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_4_12_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_4_13_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_4_14_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_4_15_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff : OUT STD_LOGIC;
      xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff : OUT STD_LOGIC;
      xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff : OUT STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_inst_p_rsc_dat : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_0_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_1_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_2_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_3_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_4_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_5_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_6_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_7_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_8_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_9_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_10_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_11_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_12_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_13_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_14_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_15_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_16_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_17_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_18_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_19_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_20_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_21_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_22_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_23_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_24_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_25_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_26_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_27_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_28_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_29_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_30_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_31_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_0_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_1_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_2_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_3_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_4_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_5_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_6_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_7_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_8_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_9_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_10_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_11_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_12_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_13_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_14_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_15_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_16_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_17_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_18_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_19_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_20_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_21_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_22_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_23_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_24_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_25_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_26_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_27_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_28_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_29_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_30_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_31_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_2_0_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_2_1_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_2_2_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_2_3_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_2_4_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_2_5_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_2_6_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_2_7_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_2_8_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_2_9_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_2_10_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_2_11_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_2_12_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_2_13_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_2_14_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_2_15_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_2_16_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_2_17_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_2_18_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_2_19_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_2_20_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_2_21_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_2_22_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_2_23_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_2_24_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_2_25_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_2_26_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_2_27_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_2_28_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_2_29_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_2_30_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_2_31_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_3_0_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_3_1_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_3_2_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_3_3_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_3_4_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_3_5_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_3_6_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_3_7_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_3_8_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_3_9_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_3_10_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_3_11_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_3_12_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_3_13_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_3_14_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_3_15_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_3_16_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_3_17_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_3_18_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_3_19_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_3_20_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_3_21_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_3_22_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_3_23_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_3_24_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_3_25_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_3_26_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_3_27_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_3_28_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_3_29_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_3_30_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_3_31_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_4_0_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_4_1_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_4_2_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_4_3_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_4_4_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_4_5_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_4_6_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_4_7_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_4_8_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_4_9_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_4_10_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_4_11_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_4_12_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_4_13_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_4_14_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_4_15_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_4_16_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_4_17_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_4_18_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_4_19_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_4_20_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_4_21_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_4_22_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_4_23_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_4_24_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_4_25_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_4_26_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_4_27_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_4_28_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_4_29_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_4_30_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_4_31_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_5_0_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_5_1_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_5_2_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_5_3_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_5_4_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_5_5_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_5_6_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_5_7_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_5_8_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_5_9_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_5_10_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_5_11_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_5_12_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_5_13_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_5_14_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_5_15_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_5_16_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_5_17_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_5_18_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_5_19_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_5_20_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_5_21_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_5_22_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_5_23_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_5_24_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_5_25_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_5_26_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_5_27_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_5_28_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_5_29_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_5_30_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_5_31_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_6_0_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_6_1_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_6_2_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_6_3_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_6_4_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_6_5_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_6_6_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_6_7_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_6_8_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_6_9_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_6_10_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_6_11_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_6_12_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_6_13_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_6_14_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_6_15_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_6_16_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_6_17_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_6_18_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_6_19_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_6_20_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_6_21_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_6_22_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_6_23_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_6_24_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_6_25_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_6_26_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_6_27_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_6_28_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_6_29_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_6_30_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_6_31_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_7_0_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_7_1_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_7_2_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_7_3_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_7_4_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_7_5_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_7_6_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_7_7_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_7_8_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_7_9_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_7_10_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_7_11_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_7_12_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_7_13_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_7_14_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_7_15_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_7_16_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_7_17_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_7_18_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_7_19_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_7_20_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_7_21_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_7_22_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_7_23_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_7_24_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_7_25_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_7_26_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_7_27_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_7_28_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_7_29_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_7_30_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_7_31_i_q_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_0_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_1_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_2_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_3_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_4_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_5_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_6_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_7_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_8_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_9_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_10_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_11_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_12_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_13_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_14_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_15_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_16_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_17_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_18_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_19_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_20_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_21_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_22_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_23_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_24_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_25_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_26_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_27_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_28_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_29_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_30_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_31_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_0_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_1_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_2_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_3_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_4_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_5_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_6_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_7_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_8_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_9_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_10_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_11_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_12_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_13_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_14_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_15_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_16_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_17_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_18_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_19_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_20_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_21_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_22_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_23_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_24_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_25_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_26_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_27_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_28_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_29_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_30_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_31_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_2_0_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_2_1_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_2_2_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_2_3_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_2_4_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_2_5_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_2_6_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_2_7_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_2_8_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_2_9_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_2_10_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_2_11_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_2_12_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_2_13_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_2_14_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_2_15_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_2_16_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_2_17_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_2_18_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_2_19_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_2_20_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_2_21_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_2_22_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_2_23_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_2_24_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_2_25_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_2_26_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_2_27_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_2_28_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_2_29_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_2_30_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_2_31_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_3_0_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_3_1_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_3_2_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_3_3_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_3_4_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_3_5_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_3_6_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_3_7_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_3_8_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_3_9_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_3_10_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_3_11_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_3_12_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_3_13_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_3_14_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_3_15_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_3_16_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_3_17_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_3_18_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_3_19_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_3_20_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_3_21_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_3_22_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_3_23_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_3_24_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_3_25_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_3_26_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_3_27_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_3_28_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_3_29_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_3_30_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_3_31_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_4_0_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_4_1_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_4_2_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_4_3_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_4_4_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_4_5_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_4_6_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_4_7_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_4_8_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_4_9_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_4_10_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_4_11_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_4_12_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_4_13_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_4_14_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_4_15_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_4_16_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_4_17_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_4_18_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_4_19_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_4_20_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_4_21_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_4_22_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_4_23_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_4_24_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_4_25_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_4_26_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_4_27_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_4_28_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_4_29_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_4_30_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_4_31_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_5_0_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_5_1_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_5_2_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_5_3_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_5_4_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_5_5_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_5_6_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_5_7_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_5_8_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_5_9_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_5_10_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_5_11_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_5_12_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_5_13_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_5_14_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_5_15_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_5_16_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_5_17_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_5_18_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_5_19_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_5_20_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_5_21_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_5_22_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_5_23_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_5_24_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_5_25_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_5_26_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_5_27_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_5_28_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_5_29_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_5_30_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_5_31_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_6_0_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_6_1_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_6_2_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_6_3_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_6_4_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_6_5_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_6_6_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_6_7_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_6_8_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_6_9_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_6_10_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_6_11_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_6_12_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_6_13_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_6_14_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_6_15_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_6_16_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_6_17_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_6_18_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_6_19_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_6_20_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_6_21_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_6_22_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_6_23_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_6_24_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_6_25_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_6_26_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_6_27_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_6_28_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_6_29_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_6_30_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_6_31_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_7_0_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_7_1_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_7_2_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_7_3_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_7_4_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_7_5_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_7_6_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_7_7_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_7_8_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_7_9_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_7_10_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_7_11_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_7_12_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_7_13_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_7_14_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_7_15_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_7_16_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_7_17_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_7_18_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_7_19_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_7_20_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_7_21_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_7_22_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_7_23_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_7_24_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_7_25_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_7_26_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_7_27_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_7_28_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_7_29_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_7_30_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_7_31_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_0_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d :
      STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_1_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_1_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d :
      STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_2_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_2_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d :
      STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_3_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_3_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d :
      STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_4_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_4_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d :
      STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_5_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_5_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d :
      STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_6_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_6_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d :
      STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_7_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_7_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d :
      STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_8_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_8_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d :
      STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_9_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_9_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d :
      STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_10_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_10_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d :
      STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_11_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_11_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d :
      STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_12_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_12_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d :
      STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_13_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_13_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d :
      STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_14_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_14_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d :
      STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_15_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_15_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d :
      STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_0_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_1_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_1_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_2_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_2_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_3_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_3_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_4_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_4_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_5_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_5_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_6_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_6_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_7_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_7_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_8_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_8_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_9_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_9_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_10_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_10_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_11_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_11_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_12_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_12_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_13_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_13_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_14_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_14_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_15_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_15_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_0_i_d_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_0_i_radr_d_pff : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_0_i_wadr_d_pff : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_1_i_d_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_1_i_wadr_d_pff : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_2_i_d_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_2_i_wadr_d_pff : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_3_i_d_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_3_i_wadr_d_pff : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_4_i_d_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_4_i_wadr_d_pff : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_5_i_d_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_5_i_wadr_d_pff : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_6_i_d_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_6_i_wadr_d_pff : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_7_i_d_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_8_i_d_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_9_i_d_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_10_i_d_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_10_i_wadr_d_pff : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_11_i_d_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_11_i_wadr_d_pff : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_12_i_d_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_13_i_d_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_14_i_d_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_15_i_d_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_4_0_i_d_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_4_0_i_wadr_d_pff : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_yt_rsc_4_1_i_d_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_4_1_i_wadr_d_pff : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_yt_rsc_4_2_i_d_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_4_2_i_wadr_d_pff : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_yt_rsc_4_3_i_d_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_4_3_i_wadr_d_pff : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_yt_rsc_4_4_i_d_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_4_4_i_wadr_d_pff : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_yt_rsc_4_5_i_d_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_4_5_i_wadr_d_pff : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_yt_rsc_4_6_i_d_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_4_6_i_wadr_d_pff : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_yt_rsc_4_7_i_d_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_4_8_i_d_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_4_9_i_d_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_4_9_i_wadr_d_pff : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_yt_rsc_4_10_i_d_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_4_10_i_wadr_d_pff : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_yt_rsc_4_11_i_d_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_4_11_i_wadr_d_pff : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_yt_rsc_4_12_i_d_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_4_13_i_d_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_4_14_i_d_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_4_15_i_d_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_0_i_adra_d_pff : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_0_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_1_i_adra_d_pff : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_1_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_2_i_adra_d_pff : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_2_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_3_i_adra_d_pff : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_3_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_4_i_adra_d_pff : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_4_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_5_i_adra_d_pff : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_5_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_6_i_adra_d_pff : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_6_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_7_i_adra_d_pff : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_7_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_8_i_adra_d_pff : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_8_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_9_i_adra_d_pff : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_9_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_10_i_adra_d_pff : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_10_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_11_i_adra_d_pff : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_11_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_12_i_adra_d_pff : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_12_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_13_i_adra_d_pff : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_13_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_14_i_adra_d_pff : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_14_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_15_i_adra_d_pff : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_15_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_xt_rsc_4_0_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_4_1_i_adra_d_pff : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_xt_rsc_4_1_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_4_2_i_adra_d_pff : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_xt_rsc_4_2_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_4_3_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_4_4_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_4_5_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_4_6_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_4_7_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_4_8_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_4_9_i_adra_d_pff : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_xt_rsc_4_9_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_4_10_i_adra_d_pff : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_xt_rsc_4_10_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_xt_rsc_4_11_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_xt_rsc_4_12_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_xt_rsc_4_13_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_xt_rsc_4_14_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_xt_rsc_4_15_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO
      0);

BEGIN
  yt_rsc_0_0_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_0_0_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_0_0_clkr_en,
      d => yt_rsc_0_0_comp_d,
      q => yt_rsc_0_0_comp_q,
      radr => yt_rsc_0_0_comp_radr,
      wadr => yt_rsc_0_0_comp_wadr,
      we => yt_rsc_0_0_we
    );
  yt_rsc_0_0_comp_d <= yt_rsc_0_0_d;
  yt_rsc_0_0_q <= yt_rsc_0_0_comp_q;
  yt_rsc_0_0_comp_radr <= yt_rsc_0_0_radr;
  yt_rsc_0_0_comp_wadr <= yt_rsc_0_0_wadr;

  yt_rsc_0_1_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_0_1_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_0_1_clkr_en,
      d => yt_rsc_0_1_comp_d,
      q => yt_rsc_0_1_comp_q,
      radr => yt_rsc_0_1_comp_radr,
      wadr => yt_rsc_0_1_comp_wadr,
      we => yt_rsc_0_1_we
    );
  yt_rsc_0_1_comp_d <= yt_rsc_0_1_d;
  yt_rsc_0_1_q <= yt_rsc_0_1_comp_q;
  yt_rsc_0_1_comp_radr <= yt_rsc_0_1_radr;
  yt_rsc_0_1_comp_wadr <= yt_rsc_0_1_wadr;

  yt_rsc_0_2_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_0_2_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_0_2_clkr_en,
      d => yt_rsc_0_2_comp_d,
      q => yt_rsc_0_2_comp_q,
      radr => yt_rsc_0_2_comp_radr,
      wadr => yt_rsc_0_2_comp_wadr,
      we => yt_rsc_0_2_we
    );
  yt_rsc_0_2_comp_d <= yt_rsc_0_2_d;
  yt_rsc_0_2_q <= yt_rsc_0_2_comp_q;
  yt_rsc_0_2_comp_radr <= yt_rsc_0_2_radr;
  yt_rsc_0_2_comp_wadr <= yt_rsc_0_2_wadr;

  yt_rsc_0_3_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_0_3_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_0_3_clkr_en,
      d => yt_rsc_0_3_comp_d,
      q => yt_rsc_0_3_comp_q,
      radr => yt_rsc_0_3_comp_radr,
      wadr => yt_rsc_0_3_comp_wadr,
      we => yt_rsc_0_3_we
    );
  yt_rsc_0_3_comp_d <= yt_rsc_0_3_d;
  yt_rsc_0_3_q <= yt_rsc_0_3_comp_q;
  yt_rsc_0_3_comp_radr <= yt_rsc_0_3_radr;
  yt_rsc_0_3_comp_wadr <= yt_rsc_0_3_wadr;

  yt_rsc_0_4_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_0_4_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_0_4_clkr_en,
      d => yt_rsc_0_4_comp_d,
      q => yt_rsc_0_4_comp_q,
      radr => yt_rsc_0_4_comp_radr,
      wadr => yt_rsc_0_4_comp_wadr,
      we => yt_rsc_0_4_we
    );
  yt_rsc_0_4_comp_d <= yt_rsc_0_4_d;
  yt_rsc_0_4_q <= yt_rsc_0_4_comp_q;
  yt_rsc_0_4_comp_radr <= yt_rsc_0_4_radr;
  yt_rsc_0_4_comp_wadr <= yt_rsc_0_4_wadr;

  yt_rsc_0_5_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_0_5_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_0_5_clkr_en,
      d => yt_rsc_0_5_comp_d,
      q => yt_rsc_0_5_comp_q,
      radr => yt_rsc_0_5_comp_radr,
      wadr => yt_rsc_0_5_comp_wadr,
      we => yt_rsc_0_5_we
    );
  yt_rsc_0_5_comp_d <= yt_rsc_0_5_d;
  yt_rsc_0_5_q <= yt_rsc_0_5_comp_q;
  yt_rsc_0_5_comp_radr <= yt_rsc_0_5_radr;
  yt_rsc_0_5_comp_wadr <= yt_rsc_0_5_wadr;

  yt_rsc_0_6_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_0_6_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_0_6_clkr_en,
      d => yt_rsc_0_6_comp_d,
      q => yt_rsc_0_6_comp_q,
      radr => yt_rsc_0_6_comp_radr,
      wadr => yt_rsc_0_6_comp_wadr,
      we => yt_rsc_0_6_we
    );
  yt_rsc_0_6_comp_d <= yt_rsc_0_6_d;
  yt_rsc_0_6_q <= yt_rsc_0_6_comp_q;
  yt_rsc_0_6_comp_radr <= yt_rsc_0_6_radr;
  yt_rsc_0_6_comp_wadr <= yt_rsc_0_6_wadr;

  yt_rsc_0_7_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_0_7_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_0_7_clkr_en,
      d => yt_rsc_0_7_comp_d,
      q => yt_rsc_0_7_comp_q,
      radr => yt_rsc_0_7_comp_radr,
      wadr => yt_rsc_0_7_comp_wadr,
      we => yt_rsc_0_7_we
    );
  yt_rsc_0_7_comp_d <= yt_rsc_0_7_d;
  yt_rsc_0_7_q <= yt_rsc_0_7_comp_q;
  yt_rsc_0_7_comp_radr <= yt_rsc_0_7_radr;
  yt_rsc_0_7_comp_wadr <= yt_rsc_0_7_wadr;

  yt_rsc_0_8_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_0_8_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_0_8_clkr_en,
      d => yt_rsc_0_8_comp_d,
      q => yt_rsc_0_8_comp_q,
      radr => yt_rsc_0_8_comp_radr,
      wadr => yt_rsc_0_8_comp_wadr,
      we => yt_rsc_0_8_we
    );
  yt_rsc_0_8_comp_d <= yt_rsc_0_8_d;
  yt_rsc_0_8_q <= yt_rsc_0_8_comp_q;
  yt_rsc_0_8_comp_radr <= yt_rsc_0_8_radr;
  yt_rsc_0_8_comp_wadr <= yt_rsc_0_8_wadr;

  yt_rsc_0_9_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_0_9_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_0_9_clkr_en,
      d => yt_rsc_0_9_comp_d,
      q => yt_rsc_0_9_comp_q,
      radr => yt_rsc_0_9_comp_radr,
      wadr => yt_rsc_0_9_comp_wadr,
      we => yt_rsc_0_9_we
    );
  yt_rsc_0_9_comp_d <= yt_rsc_0_9_d;
  yt_rsc_0_9_q <= yt_rsc_0_9_comp_q;
  yt_rsc_0_9_comp_radr <= yt_rsc_0_9_radr;
  yt_rsc_0_9_comp_wadr <= yt_rsc_0_9_wadr;

  yt_rsc_0_10_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_0_10_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_0_10_clkr_en,
      d => yt_rsc_0_10_comp_d,
      q => yt_rsc_0_10_comp_q,
      radr => yt_rsc_0_10_comp_radr,
      wadr => yt_rsc_0_10_comp_wadr,
      we => yt_rsc_0_10_we
    );
  yt_rsc_0_10_comp_d <= yt_rsc_0_10_d;
  yt_rsc_0_10_q <= yt_rsc_0_10_comp_q;
  yt_rsc_0_10_comp_radr <= yt_rsc_0_10_radr;
  yt_rsc_0_10_comp_wadr <= yt_rsc_0_10_wadr;

  yt_rsc_0_11_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_0_11_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_0_11_clkr_en,
      d => yt_rsc_0_11_comp_d,
      q => yt_rsc_0_11_comp_q,
      radr => yt_rsc_0_11_comp_radr,
      wadr => yt_rsc_0_11_comp_wadr,
      we => yt_rsc_0_11_we
    );
  yt_rsc_0_11_comp_d <= yt_rsc_0_11_d;
  yt_rsc_0_11_q <= yt_rsc_0_11_comp_q;
  yt_rsc_0_11_comp_radr <= yt_rsc_0_11_radr;
  yt_rsc_0_11_comp_wadr <= yt_rsc_0_11_wadr;

  yt_rsc_0_12_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_0_12_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_0_12_clkr_en,
      d => yt_rsc_0_12_comp_d,
      q => yt_rsc_0_12_comp_q,
      radr => yt_rsc_0_12_comp_radr,
      wadr => yt_rsc_0_12_comp_wadr,
      we => yt_rsc_0_12_we
    );
  yt_rsc_0_12_comp_d <= yt_rsc_0_12_d;
  yt_rsc_0_12_q <= yt_rsc_0_12_comp_q;
  yt_rsc_0_12_comp_radr <= yt_rsc_0_12_radr;
  yt_rsc_0_12_comp_wadr <= yt_rsc_0_12_wadr;

  yt_rsc_0_13_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_0_13_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_0_13_clkr_en,
      d => yt_rsc_0_13_comp_d,
      q => yt_rsc_0_13_comp_q,
      radr => yt_rsc_0_13_comp_radr,
      wadr => yt_rsc_0_13_comp_wadr,
      we => yt_rsc_0_13_we
    );
  yt_rsc_0_13_comp_d <= yt_rsc_0_13_d;
  yt_rsc_0_13_q <= yt_rsc_0_13_comp_q;
  yt_rsc_0_13_comp_radr <= yt_rsc_0_13_radr;
  yt_rsc_0_13_comp_wadr <= yt_rsc_0_13_wadr;

  yt_rsc_0_14_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_0_14_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_0_14_clkr_en,
      d => yt_rsc_0_14_comp_d,
      q => yt_rsc_0_14_comp_q,
      radr => yt_rsc_0_14_comp_radr,
      wadr => yt_rsc_0_14_comp_wadr,
      we => yt_rsc_0_14_we
    );
  yt_rsc_0_14_comp_d <= yt_rsc_0_14_d;
  yt_rsc_0_14_q <= yt_rsc_0_14_comp_q;
  yt_rsc_0_14_comp_radr <= yt_rsc_0_14_radr;
  yt_rsc_0_14_comp_wadr <= yt_rsc_0_14_wadr;

  yt_rsc_0_15_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_0_15_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_0_15_clkr_en,
      d => yt_rsc_0_15_comp_d,
      q => yt_rsc_0_15_comp_q,
      radr => yt_rsc_0_15_comp_radr,
      wadr => yt_rsc_0_15_comp_wadr,
      we => yt_rsc_0_15_we
    );
  yt_rsc_0_15_comp_d <= yt_rsc_0_15_d;
  yt_rsc_0_15_q <= yt_rsc_0_15_comp_q;
  yt_rsc_0_15_comp_radr <= yt_rsc_0_15_radr;
  yt_rsc_0_15_comp_wadr <= yt_rsc_0_15_wadr;

  yt_rsc_0_16_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_0_16_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_0_16_clkr_en,
      d => yt_rsc_0_16_comp_d,
      q => yt_rsc_0_16_comp_q,
      radr => yt_rsc_0_16_comp_radr,
      wadr => yt_rsc_0_16_comp_wadr,
      we => yt_rsc_0_16_we
    );
  yt_rsc_0_16_comp_d <= yt_rsc_0_16_d;
  yt_rsc_0_16_q <= yt_rsc_0_16_comp_q;
  yt_rsc_0_16_comp_radr <= yt_rsc_0_16_radr;
  yt_rsc_0_16_comp_wadr <= yt_rsc_0_16_wadr;

  yt_rsc_0_17_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_0_17_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_0_17_clkr_en,
      d => yt_rsc_0_17_comp_d,
      q => yt_rsc_0_17_comp_q,
      radr => yt_rsc_0_17_comp_radr,
      wadr => yt_rsc_0_17_comp_wadr,
      we => yt_rsc_0_17_we
    );
  yt_rsc_0_17_comp_d <= yt_rsc_0_17_d;
  yt_rsc_0_17_q <= yt_rsc_0_17_comp_q;
  yt_rsc_0_17_comp_radr <= yt_rsc_0_17_radr;
  yt_rsc_0_17_comp_wadr <= yt_rsc_0_17_wadr;

  yt_rsc_0_18_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_0_18_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_0_18_clkr_en,
      d => yt_rsc_0_18_comp_d,
      q => yt_rsc_0_18_comp_q,
      radr => yt_rsc_0_18_comp_radr,
      wadr => yt_rsc_0_18_comp_wadr,
      we => yt_rsc_0_18_we
    );
  yt_rsc_0_18_comp_d <= yt_rsc_0_18_d;
  yt_rsc_0_18_q <= yt_rsc_0_18_comp_q;
  yt_rsc_0_18_comp_radr <= yt_rsc_0_18_radr;
  yt_rsc_0_18_comp_wadr <= yt_rsc_0_18_wadr;

  yt_rsc_0_19_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_0_19_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_0_19_clkr_en,
      d => yt_rsc_0_19_comp_d,
      q => yt_rsc_0_19_comp_q,
      radr => yt_rsc_0_19_comp_radr,
      wadr => yt_rsc_0_19_comp_wadr,
      we => yt_rsc_0_19_we
    );
  yt_rsc_0_19_comp_d <= yt_rsc_0_19_d;
  yt_rsc_0_19_q <= yt_rsc_0_19_comp_q;
  yt_rsc_0_19_comp_radr <= yt_rsc_0_19_radr;
  yt_rsc_0_19_comp_wadr <= yt_rsc_0_19_wadr;

  yt_rsc_0_20_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_0_20_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_0_20_clkr_en,
      d => yt_rsc_0_20_comp_d,
      q => yt_rsc_0_20_comp_q,
      radr => yt_rsc_0_20_comp_radr,
      wadr => yt_rsc_0_20_comp_wadr,
      we => yt_rsc_0_20_we
    );
  yt_rsc_0_20_comp_d <= yt_rsc_0_20_d;
  yt_rsc_0_20_q <= yt_rsc_0_20_comp_q;
  yt_rsc_0_20_comp_radr <= yt_rsc_0_20_radr;
  yt_rsc_0_20_comp_wadr <= yt_rsc_0_20_wadr;

  yt_rsc_0_21_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_0_21_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_0_21_clkr_en,
      d => yt_rsc_0_21_comp_d,
      q => yt_rsc_0_21_comp_q,
      radr => yt_rsc_0_21_comp_radr,
      wadr => yt_rsc_0_21_comp_wadr,
      we => yt_rsc_0_21_we
    );
  yt_rsc_0_21_comp_d <= yt_rsc_0_21_d;
  yt_rsc_0_21_q <= yt_rsc_0_21_comp_q;
  yt_rsc_0_21_comp_radr <= yt_rsc_0_21_radr;
  yt_rsc_0_21_comp_wadr <= yt_rsc_0_21_wadr;

  yt_rsc_0_22_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_0_22_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_0_22_clkr_en,
      d => yt_rsc_0_22_comp_d,
      q => yt_rsc_0_22_comp_q,
      radr => yt_rsc_0_22_comp_radr,
      wadr => yt_rsc_0_22_comp_wadr,
      we => yt_rsc_0_22_we
    );
  yt_rsc_0_22_comp_d <= yt_rsc_0_22_d;
  yt_rsc_0_22_q <= yt_rsc_0_22_comp_q;
  yt_rsc_0_22_comp_radr <= yt_rsc_0_22_radr;
  yt_rsc_0_22_comp_wadr <= yt_rsc_0_22_wadr;

  yt_rsc_0_23_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_0_23_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_0_23_clkr_en,
      d => yt_rsc_0_23_comp_d,
      q => yt_rsc_0_23_comp_q,
      radr => yt_rsc_0_23_comp_radr,
      wadr => yt_rsc_0_23_comp_wadr,
      we => yt_rsc_0_23_we
    );
  yt_rsc_0_23_comp_d <= yt_rsc_0_23_d;
  yt_rsc_0_23_q <= yt_rsc_0_23_comp_q;
  yt_rsc_0_23_comp_radr <= yt_rsc_0_23_radr;
  yt_rsc_0_23_comp_wadr <= yt_rsc_0_23_wadr;

  yt_rsc_0_24_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_0_24_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_0_24_clkr_en,
      d => yt_rsc_0_24_comp_d,
      q => yt_rsc_0_24_comp_q,
      radr => yt_rsc_0_24_comp_radr,
      wadr => yt_rsc_0_24_comp_wadr,
      we => yt_rsc_0_24_we
    );
  yt_rsc_0_24_comp_d <= yt_rsc_0_24_d;
  yt_rsc_0_24_q <= yt_rsc_0_24_comp_q;
  yt_rsc_0_24_comp_radr <= yt_rsc_0_24_radr;
  yt_rsc_0_24_comp_wadr <= yt_rsc_0_24_wadr;

  yt_rsc_0_25_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_0_25_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_0_25_clkr_en,
      d => yt_rsc_0_25_comp_d,
      q => yt_rsc_0_25_comp_q,
      radr => yt_rsc_0_25_comp_radr,
      wadr => yt_rsc_0_25_comp_wadr,
      we => yt_rsc_0_25_we
    );
  yt_rsc_0_25_comp_d <= yt_rsc_0_25_d;
  yt_rsc_0_25_q <= yt_rsc_0_25_comp_q;
  yt_rsc_0_25_comp_radr <= yt_rsc_0_25_radr;
  yt_rsc_0_25_comp_wadr <= yt_rsc_0_25_wadr;

  yt_rsc_0_26_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_0_26_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_0_26_clkr_en,
      d => yt_rsc_0_26_comp_d,
      q => yt_rsc_0_26_comp_q,
      radr => yt_rsc_0_26_comp_radr,
      wadr => yt_rsc_0_26_comp_wadr,
      we => yt_rsc_0_26_we
    );
  yt_rsc_0_26_comp_d <= yt_rsc_0_26_d;
  yt_rsc_0_26_q <= yt_rsc_0_26_comp_q;
  yt_rsc_0_26_comp_radr <= yt_rsc_0_26_radr;
  yt_rsc_0_26_comp_wadr <= yt_rsc_0_26_wadr;

  yt_rsc_0_27_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_0_27_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_0_27_clkr_en,
      d => yt_rsc_0_27_comp_d,
      q => yt_rsc_0_27_comp_q,
      radr => yt_rsc_0_27_comp_radr,
      wadr => yt_rsc_0_27_comp_wadr,
      we => yt_rsc_0_27_we
    );
  yt_rsc_0_27_comp_d <= yt_rsc_0_27_d;
  yt_rsc_0_27_q <= yt_rsc_0_27_comp_q;
  yt_rsc_0_27_comp_radr <= yt_rsc_0_27_radr;
  yt_rsc_0_27_comp_wadr <= yt_rsc_0_27_wadr;

  yt_rsc_0_28_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_0_28_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_0_28_clkr_en,
      d => yt_rsc_0_28_comp_d,
      q => yt_rsc_0_28_comp_q,
      radr => yt_rsc_0_28_comp_radr,
      wadr => yt_rsc_0_28_comp_wadr,
      we => yt_rsc_0_28_we
    );
  yt_rsc_0_28_comp_d <= yt_rsc_0_28_d;
  yt_rsc_0_28_q <= yt_rsc_0_28_comp_q;
  yt_rsc_0_28_comp_radr <= yt_rsc_0_28_radr;
  yt_rsc_0_28_comp_wadr <= yt_rsc_0_28_wadr;

  yt_rsc_0_29_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_0_29_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_0_29_clkr_en,
      d => yt_rsc_0_29_comp_d,
      q => yt_rsc_0_29_comp_q,
      radr => yt_rsc_0_29_comp_radr,
      wadr => yt_rsc_0_29_comp_wadr,
      we => yt_rsc_0_29_we
    );
  yt_rsc_0_29_comp_d <= yt_rsc_0_29_d;
  yt_rsc_0_29_q <= yt_rsc_0_29_comp_q;
  yt_rsc_0_29_comp_radr <= yt_rsc_0_29_radr;
  yt_rsc_0_29_comp_wadr <= yt_rsc_0_29_wadr;

  yt_rsc_0_30_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_0_30_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_0_30_clkr_en,
      d => yt_rsc_0_30_comp_d,
      q => yt_rsc_0_30_comp_q,
      radr => yt_rsc_0_30_comp_radr,
      wadr => yt_rsc_0_30_comp_wadr,
      we => yt_rsc_0_30_we
    );
  yt_rsc_0_30_comp_d <= yt_rsc_0_30_d;
  yt_rsc_0_30_q <= yt_rsc_0_30_comp_q;
  yt_rsc_0_30_comp_radr <= yt_rsc_0_30_radr;
  yt_rsc_0_30_comp_wadr <= yt_rsc_0_30_wadr;

  yt_rsc_0_31_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_0_31_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_0_31_clkr_en,
      d => yt_rsc_0_31_comp_d,
      q => yt_rsc_0_31_comp_q,
      radr => yt_rsc_0_31_comp_radr,
      wadr => yt_rsc_0_31_comp_wadr,
      we => yt_rsc_0_31_we
    );
  yt_rsc_0_31_comp_d <= yt_rsc_0_31_d;
  yt_rsc_0_31_q <= yt_rsc_0_31_comp_q;
  yt_rsc_0_31_comp_radr <= yt_rsc_0_31_radr;
  yt_rsc_0_31_comp_wadr <= yt_rsc_0_31_wadr;

  yt_rsc_1_0_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_1_0_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_1_0_clkr_en,
      d => yt_rsc_1_0_comp_d,
      q => yt_rsc_1_0_comp_q,
      radr => yt_rsc_1_0_comp_radr,
      wadr => yt_rsc_1_0_comp_wadr,
      we => yt_rsc_1_0_we
    );
  yt_rsc_1_0_comp_d <= yt_rsc_1_0_d;
  yt_rsc_1_0_q <= yt_rsc_1_0_comp_q;
  yt_rsc_1_0_comp_radr <= yt_rsc_1_0_radr;
  yt_rsc_1_0_comp_wadr <= yt_rsc_1_0_wadr;

  yt_rsc_1_1_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_1_1_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_1_1_clkr_en,
      d => yt_rsc_1_1_comp_d,
      q => yt_rsc_1_1_comp_q,
      radr => yt_rsc_1_1_comp_radr,
      wadr => yt_rsc_1_1_comp_wadr,
      we => yt_rsc_1_1_we
    );
  yt_rsc_1_1_comp_d <= yt_rsc_1_1_d;
  yt_rsc_1_1_q <= yt_rsc_1_1_comp_q;
  yt_rsc_1_1_comp_radr <= yt_rsc_1_1_radr;
  yt_rsc_1_1_comp_wadr <= yt_rsc_1_1_wadr;

  yt_rsc_1_2_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_1_2_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_1_2_clkr_en,
      d => yt_rsc_1_2_comp_d,
      q => yt_rsc_1_2_comp_q,
      radr => yt_rsc_1_2_comp_radr,
      wadr => yt_rsc_1_2_comp_wadr,
      we => yt_rsc_1_2_we
    );
  yt_rsc_1_2_comp_d <= yt_rsc_1_2_d;
  yt_rsc_1_2_q <= yt_rsc_1_2_comp_q;
  yt_rsc_1_2_comp_radr <= yt_rsc_1_2_radr;
  yt_rsc_1_2_comp_wadr <= yt_rsc_1_2_wadr;

  yt_rsc_1_3_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_1_3_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_1_3_clkr_en,
      d => yt_rsc_1_3_comp_d,
      q => yt_rsc_1_3_comp_q,
      radr => yt_rsc_1_3_comp_radr,
      wadr => yt_rsc_1_3_comp_wadr,
      we => yt_rsc_1_3_we
    );
  yt_rsc_1_3_comp_d <= yt_rsc_1_3_d;
  yt_rsc_1_3_q <= yt_rsc_1_3_comp_q;
  yt_rsc_1_3_comp_radr <= yt_rsc_1_3_radr;
  yt_rsc_1_3_comp_wadr <= yt_rsc_1_3_wadr;

  yt_rsc_1_4_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_1_4_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_1_4_clkr_en,
      d => yt_rsc_1_4_comp_d,
      q => yt_rsc_1_4_comp_q,
      radr => yt_rsc_1_4_comp_radr,
      wadr => yt_rsc_1_4_comp_wadr,
      we => yt_rsc_1_4_we
    );
  yt_rsc_1_4_comp_d <= yt_rsc_1_4_d;
  yt_rsc_1_4_q <= yt_rsc_1_4_comp_q;
  yt_rsc_1_4_comp_radr <= yt_rsc_1_4_radr;
  yt_rsc_1_4_comp_wadr <= yt_rsc_1_4_wadr;

  yt_rsc_1_5_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_1_5_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_1_5_clkr_en,
      d => yt_rsc_1_5_comp_d,
      q => yt_rsc_1_5_comp_q,
      radr => yt_rsc_1_5_comp_radr,
      wadr => yt_rsc_1_5_comp_wadr,
      we => yt_rsc_1_5_we
    );
  yt_rsc_1_5_comp_d <= yt_rsc_1_5_d;
  yt_rsc_1_5_q <= yt_rsc_1_5_comp_q;
  yt_rsc_1_5_comp_radr <= yt_rsc_1_5_radr;
  yt_rsc_1_5_comp_wadr <= yt_rsc_1_5_wadr;

  yt_rsc_1_6_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_1_6_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_1_6_clkr_en,
      d => yt_rsc_1_6_comp_d,
      q => yt_rsc_1_6_comp_q,
      radr => yt_rsc_1_6_comp_radr,
      wadr => yt_rsc_1_6_comp_wadr,
      we => yt_rsc_1_6_we
    );
  yt_rsc_1_6_comp_d <= yt_rsc_1_6_d;
  yt_rsc_1_6_q <= yt_rsc_1_6_comp_q;
  yt_rsc_1_6_comp_radr <= yt_rsc_1_6_radr;
  yt_rsc_1_6_comp_wadr <= yt_rsc_1_6_wadr;

  yt_rsc_1_7_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_1_7_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_1_7_clkr_en,
      d => yt_rsc_1_7_comp_d,
      q => yt_rsc_1_7_comp_q,
      radr => yt_rsc_1_7_comp_radr,
      wadr => yt_rsc_1_7_comp_wadr,
      we => yt_rsc_1_7_we
    );
  yt_rsc_1_7_comp_d <= yt_rsc_1_7_d;
  yt_rsc_1_7_q <= yt_rsc_1_7_comp_q;
  yt_rsc_1_7_comp_radr <= yt_rsc_1_7_radr;
  yt_rsc_1_7_comp_wadr <= yt_rsc_1_7_wadr;

  yt_rsc_1_8_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_1_8_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_1_8_clkr_en,
      d => yt_rsc_1_8_comp_d,
      q => yt_rsc_1_8_comp_q,
      radr => yt_rsc_1_8_comp_radr,
      wadr => yt_rsc_1_8_comp_wadr,
      we => yt_rsc_1_8_we
    );
  yt_rsc_1_8_comp_d <= yt_rsc_1_8_d;
  yt_rsc_1_8_q <= yt_rsc_1_8_comp_q;
  yt_rsc_1_8_comp_radr <= yt_rsc_1_8_radr;
  yt_rsc_1_8_comp_wadr <= yt_rsc_1_8_wadr;

  yt_rsc_1_9_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_1_9_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_1_9_clkr_en,
      d => yt_rsc_1_9_comp_d,
      q => yt_rsc_1_9_comp_q,
      radr => yt_rsc_1_9_comp_radr,
      wadr => yt_rsc_1_9_comp_wadr,
      we => yt_rsc_1_9_we
    );
  yt_rsc_1_9_comp_d <= yt_rsc_1_9_d;
  yt_rsc_1_9_q <= yt_rsc_1_9_comp_q;
  yt_rsc_1_9_comp_radr <= yt_rsc_1_9_radr;
  yt_rsc_1_9_comp_wadr <= yt_rsc_1_9_wadr;

  yt_rsc_1_10_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_1_10_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_1_10_clkr_en,
      d => yt_rsc_1_10_comp_d,
      q => yt_rsc_1_10_comp_q,
      radr => yt_rsc_1_10_comp_radr,
      wadr => yt_rsc_1_10_comp_wadr,
      we => yt_rsc_1_10_we
    );
  yt_rsc_1_10_comp_d <= yt_rsc_1_10_d;
  yt_rsc_1_10_q <= yt_rsc_1_10_comp_q;
  yt_rsc_1_10_comp_radr <= yt_rsc_1_10_radr;
  yt_rsc_1_10_comp_wadr <= yt_rsc_1_10_wadr;

  yt_rsc_1_11_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_1_11_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_1_11_clkr_en,
      d => yt_rsc_1_11_comp_d,
      q => yt_rsc_1_11_comp_q,
      radr => yt_rsc_1_11_comp_radr,
      wadr => yt_rsc_1_11_comp_wadr,
      we => yt_rsc_1_11_we
    );
  yt_rsc_1_11_comp_d <= yt_rsc_1_11_d;
  yt_rsc_1_11_q <= yt_rsc_1_11_comp_q;
  yt_rsc_1_11_comp_radr <= yt_rsc_1_11_radr;
  yt_rsc_1_11_comp_wadr <= yt_rsc_1_11_wadr;

  yt_rsc_1_12_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_1_12_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_1_12_clkr_en,
      d => yt_rsc_1_12_comp_d,
      q => yt_rsc_1_12_comp_q,
      radr => yt_rsc_1_12_comp_radr,
      wadr => yt_rsc_1_12_comp_wadr,
      we => yt_rsc_1_12_we
    );
  yt_rsc_1_12_comp_d <= yt_rsc_1_12_d;
  yt_rsc_1_12_q <= yt_rsc_1_12_comp_q;
  yt_rsc_1_12_comp_radr <= yt_rsc_1_12_radr;
  yt_rsc_1_12_comp_wadr <= yt_rsc_1_12_wadr;

  yt_rsc_1_13_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_1_13_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_1_13_clkr_en,
      d => yt_rsc_1_13_comp_d,
      q => yt_rsc_1_13_comp_q,
      radr => yt_rsc_1_13_comp_radr,
      wadr => yt_rsc_1_13_comp_wadr,
      we => yt_rsc_1_13_we
    );
  yt_rsc_1_13_comp_d <= yt_rsc_1_13_d;
  yt_rsc_1_13_q <= yt_rsc_1_13_comp_q;
  yt_rsc_1_13_comp_radr <= yt_rsc_1_13_radr;
  yt_rsc_1_13_comp_wadr <= yt_rsc_1_13_wadr;

  yt_rsc_1_14_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_1_14_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_1_14_clkr_en,
      d => yt_rsc_1_14_comp_d,
      q => yt_rsc_1_14_comp_q,
      radr => yt_rsc_1_14_comp_radr,
      wadr => yt_rsc_1_14_comp_wadr,
      we => yt_rsc_1_14_we
    );
  yt_rsc_1_14_comp_d <= yt_rsc_1_14_d;
  yt_rsc_1_14_q <= yt_rsc_1_14_comp_q;
  yt_rsc_1_14_comp_radr <= yt_rsc_1_14_radr;
  yt_rsc_1_14_comp_wadr <= yt_rsc_1_14_wadr;

  yt_rsc_1_15_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_1_15_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_1_15_clkr_en,
      d => yt_rsc_1_15_comp_d,
      q => yt_rsc_1_15_comp_q,
      radr => yt_rsc_1_15_comp_radr,
      wadr => yt_rsc_1_15_comp_wadr,
      we => yt_rsc_1_15_we
    );
  yt_rsc_1_15_comp_d <= yt_rsc_1_15_d;
  yt_rsc_1_15_q <= yt_rsc_1_15_comp_q;
  yt_rsc_1_15_comp_radr <= yt_rsc_1_15_radr;
  yt_rsc_1_15_comp_wadr <= yt_rsc_1_15_wadr;

  yt_rsc_1_16_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_1_16_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_1_16_clkr_en,
      d => yt_rsc_1_16_comp_d,
      q => yt_rsc_1_16_comp_q,
      radr => yt_rsc_1_16_comp_radr,
      wadr => yt_rsc_1_16_comp_wadr,
      we => yt_rsc_1_16_we
    );
  yt_rsc_1_16_comp_d <= yt_rsc_1_16_d;
  yt_rsc_1_16_q <= yt_rsc_1_16_comp_q;
  yt_rsc_1_16_comp_radr <= yt_rsc_1_16_radr;
  yt_rsc_1_16_comp_wadr <= yt_rsc_1_16_wadr;

  yt_rsc_1_17_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_1_17_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_1_17_clkr_en,
      d => yt_rsc_1_17_comp_d,
      q => yt_rsc_1_17_comp_q,
      radr => yt_rsc_1_17_comp_radr,
      wadr => yt_rsc_1_17_comp_wadr,
      we => yt_rsc_1_17_we
    );
  yt_rsc_1_17_comp_d <= yt_rsc_1_17_d;
  yt_rsc_1_17_q <= yt_rsc_1_17_comp_q;
  yt_rsc_1_17_comp_radr <= yt_rsc_1_17_radr;
  yt_rsc_1_17_comp_wadr <= yt_rsc_1_17_wadr;

  yt_rsc_1_18_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_1_18_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_1_18_clkr_en,
      d => yt_rsc_1_18_comp_d,
      q => yt_rsc_1_18_comp_q,
      radr => yt_rsc_1_18_comp_radr,
      wadr => yt_rsc_1_18_comp_wadr,
      we => yt_rsc_1_18_we
    );
  yt_rsc_1_18_comp_d <= yt_rsc_1_18_d;
  yt_rsc_1_18_q <= yt_rsc_1_18_comp_q;
  yt_rsc_1_18_comp_radr <= yt_rsc_1_18_radr;
  yt_rsc_1_18_comp_wadr <= yt_rsc_1_18_wadr;

  yt_rsc_1_19_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_1_19_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_1_19_clkr_en,
      d => yt_rsc_1_19_comp_d,
      q => yt_rsc_1_19_comp_q,
      radr => yt_rsc_1_19_comp_radr,
      wadr => yt_rsc_1_19_comp_wadr,
      we => yt_rsc_1_19_we
    );
  yt_rsc_1_19_comp_d <= yt_rsc_1_19_d;
  yt_rsc_1_19_q <= yt_rsc_1_19_comp_q;
  yt_rsc_1_19_comp_radr <= yt_rsc_1_19_radr;
  yt_rsc_1_19_comp_wadr <= yt_rsc_1_19_wadr;

  yt_rsc_1_20_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_1_20_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_1_20_clkr_en,
      d => yt_rsc_1_20_comp_d,
      q => yt_rsc_1_20_comp_q,
      radr => yt_rsc_1_20_comp_radr,
      wadr => yt_rsc_1_20_comp_wadr,
      we => yt_rsc_1_20_we
    );
  yt_rsc_1_20_comp_d <= yt_rsc_1_20_d;
  yt_rsc_1_20_q <= yt_rsc_1_20_comp_q;
  yt_rsc_1_20_comp_radr <= yt_rsc_1_20_radr;
  yt_rsc_1_20_comp_wadr <= yt_rsc_1_20_wadr;

  yt_rsc_1_21_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_1_21_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_1_21_clkr_en,
      d => yt_rsc_1_21_comp_d,
      q => yt_rsc_1_21_comp_q,
      radr => yt_rsc_1_21_comp_radr,
      wadr => yt_rsc_1_21_comp_wadr,
      we => yt_rsc_1_21_we
    );
  yt_rsc_1_21_comp_d <= yt_rsc_1_21_d;
  yt_rsc_1_21_q <= yt_rsc_1_21_comp_q;
  yt_rsc_1_21_comp_radr <= yt_rsc_1_21_radr;
  yt_rsc_1_21_comp_wadr <= yt_rsc_1_21_wadr;

  yt_rsc_1_22_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_1_22_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_1_22_clkr_en,
      d => yt_rsc_1_22_comp_d,
      q => yt_rsc_1_22_comp_q,
      radr => yt_rsc_1_22_comp_radr,
      wadr => yt_rsc_1_22_comp_wadr,
      we => yt_rsc_1_22_we
    );
  yt_rsc_1_22_comp_d <= yt_rsc_1_22_d;
  yt_rsc_1_22_q <= yt_rsc_1_22_comp_q;
  yt_rsc_1_22_comp_radr <= yt_rsc_1_22_radr;
  yt_rsc_1_22_comp_wadr <= yt_rsc_1_22_wadr;

  yt_rsc_1_23_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_1_23_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_1_23_clkr_en,
      d => yt_rsc_1_23_comp_d,
      q => yt_rsc_1_23_comp_q,
      radr => yt_rsc_1_23_comp_radr,
      wadr => yt_rsc_1_23_comp_wadr,
      we => yt_rsc_1_23_we
    );
  yt_rsc_1_23_comp_d <= yt_rsc_1_23_d;
  yt_rsc_1_23_q <= yt_rsc_1_23_comp_q;
  yt_rsc_1_23_comp_radr <= yt_rsc_1_23_radr;
  yt_rsc_1_23_comp_wadr <= yt_rsc_1_23_wadr;

  yt_rsc_1_24_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_1_24_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_1_24_clkr_en,
      d => yt_rsc_1_24_comp_d,
      q => yt_rsc_1_24_comp_q,
      radr => yt_rsc_1_24_comp_radr,
      wadr => yt_rsc_1_24_comp_wadr,
      we => yt_rsc_1_24_we
    );
  yt_rsc_1_24_comp_d <= yt_rsc_1_24_d;
  yt_rsc_1_24_q <= yt_rsc_1_24_comp_q;
  yt_rsc_1_24_comp_radr <= yt_rsc_1_24_radr;
  yt_rsc_1_24_comp_wadr <= yt_rsc_1_24_wadr;

  yt_rsc_1_25_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_1_25_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_1_25_clkr_en,
      d => yt_rsc_1_25_comp_d,
      q => yt_rsc_1_25_comp_q,
      radr => yt_rsc_1_25_comp_radr,
      wadr => yt_rsc_1_25_comp_wadr,
      we => yt_rsc_1_25_we
    );
  yt_rsc_1_25_comp_d <= yt_rsc_1_25_d;
  yt_rsc_1_25_q <= yt_rsc_1_25_comp_q;
  yt_rsc_1_25_comp_radr <= yt_rsc_1_25_radr;
  yt_rsc_1_25_comp_wadr <= yt_rsc_1_25_wadr;

  yt_rsc_1_26_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_1_26_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_1_26_clkr_en,
      d => yt_rsc_1_26_comp_d,
      q => yt_rsc_1_26_comp_q,
      radr => yt_rsc_1_26_comp_radr,
      wadr => yt_rsc_1_26_comp_wadr,
      we => yt_rsc_1_26_we
    );
  yt_rsc_1_26_comp_d <= yt_rsc_1_26_d;
  yt_rsc_1_26_q <= yt_rsc_1_26_comp_q;
  yt_rsc_1_26_comp_radr <= yt_rsc_1_26_radr;
  yt_rsc_1_26_comp_wadr <= yt_rsc_1_26_wadr;

  yt_rsc_1_27_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_1_27_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_1_27_clkr_en,
      d => yt_rsc_1_27_comp_d,
      q => yt_rsc_1_27_comp_q,
      radr => yt_rsc_1_27_comp_radr,
      wadr => yt_rsc_1_27_comp_wadr,
      we => yt_rsc_1_27_we
    );
  yt_rsc_1_27_comp_d <= yt_rsc_1_27_d;
  yt_rsc_1_27_q <= yt_rsc_1_27_comp_q;
  yt_rsc_1_27_comp_radr <= yt_rsc_1_27_radr;
  yt_rsc_1_27_comp_wadr <= yt_rsc_1_27_wadr;

  yt_rsc_1_28_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_1_28_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_1_28_clkr_en,
      d => yt_rsc_1_28_comp_d,
      q => yt_rsc_1_28_comp_q,
      radr => yt_rsc_1_28_comp_radr,
      wadr => yt_rsc_1_28_comp_wadr,
      we => yt_rsc_1_28_we
    );
  yt_rsc_1_28_comp_d <= yt_rsc_1_28_d;
  yt_rsc_1_28_q <= yt_rsc_1_28_comp_q;
  yt_rsc_1_28_comp_radr <= yt_rsc_1_28_radr;
  yt_rsc_1_28_comp_wadr <= yt_rsc_1_28_wadr;

  yt_rsc_1_29_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_1_29_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_1_29_clkr_en,
      d => yt_rsc_1_29_comp_d,
      q => yt_rsc_1_29_comp_q,
      radr => yt_rsc_1_29_comp_radr,
      wadr => yt_rsc_1_29_comp_wadr,
      we => yt_rsc_1_29_we
    );
  yt_rsc_1_29_comp_d <= yt_rsc_1_29_d;
  yt_rsc_1_29_q <= yt_rsc_1_29_comp_q;
  yt_rsc_1_29_comp_radr <= yt_rsc_1_29_radr;
  yt_rsc_1_29_comp_wadr <= yt_rsc_1_29_wadr;

  yt_rsc_1_30_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_1_30_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_1_30_clkr_en,
      d => yt_rsc_1_30_comp_d,
      q => yt_rsc_1_30_comp_q,
      radr => yt_rsc_1_30_comp_radr,
      wadr => yt_rsc_1_30_comp_wadr,
      we => yt_rsc_1_30_we
    );
  yt_rsc_1_30_comp_d <= yt_rsc_1_30_d;
  yt_rsc_1_30_q <= yt_rsc_1_30_comp_q;
  yt_rsc_1_30_comp_radr <= yt_rsc_1_30_radr;
  yt_rsc_1_30_comp_wadr <= yt_rsc_1_30_wadr;

  yt_rsc_1_31_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_1_31_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_1_31_clkr_en,
      d => yt_rsc_1_31_comp_d,
      q => yt_rsc_1_31_comp_q,
      radr => yt_rsc_1_31_comp_radr,
      wadr => yt_rsc_1_31_comp_wadr,
      we => yt_rsc_1_31_we
    );
  yt_rsc_1_31_comp_d <= yt_rsc_1_31_d;
  yt_rsc_1_31_q <= yt_rsc_1_31_comp_q;
  yt_rsc_1_31_comp_radr <= yt_rsc_1_31_radr;
  yt_rsc_1_31_comp_wadr <= yt_rsc_1_31_wadr;

  yt_rsc_2_0_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_2_0_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_2_0_clkr_en,
      d => yt_rsc_2_0_comp_d,
      q => yt_rsc_2_0_comp_q,
      radr => yt_rsc_2_0_comp_radr,
      wadr => yt_rsc_2_0_comp_wadr,
      we => yt_rsc_2_0_we
    );
  yt_rsc_2_0_comp_d <= yt_rsc_2_0_d;
  yt_rsc_2_0_q <= yt_rsc_2_0_comp_q;
  yt_rsc_2_0_comp_radr <= yt_rsc_2_0_radr;
  yt_rsc_2_0_comp_wadr <= yt_rsc_2_0_wadr;

  yt_rsc_2_1_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_2_1_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_2_1_clkr_en,
      d => yt_rsc_2_1_comp_d,
      q => yt_rsc_2_1_comp_q,
      radr => yt_rsc_2_1_comp_radr,
      wadr => yt_rsc_2_1_comp_wadr,
      we => yt_rsc_2_1_we
    );
  yt_rsc_2_1_comp_d <= yt_rsc_2_1_d;
  yt_rsc_2_1_q <= yt_rsc_2_1_comp_q;
  yt_rsc_2_1_comp_radr <= yt_rsc_2_1_radr;
  yt_rsc_2_1_comp_wadr <= yt_rsc_2_1_wadr;

  yt_rsc_2_2_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_2_2_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_2_2_clkr_en,
      d => yt_rsc_2_2_comp_d,
      q => yt_rsc_2_2_comp_q,
      radr => yt_rsc_2_2_comp_radr,
      wadr => yt_rsc_2_2_comp_wadr,
      we => yt_rsc_2_2_we
    );
  yt_rsc_2_2_comp_d <= yt_rsc_2_2_d;
  yt_rsc_2_2_q <= yt_rsc_2_2_comp_q;
  yt_rsc_2_2_comp_radr <= yt_rsc_2_2_radr;
  yt_rsc_2_2_comp_wadr <= yt_rsc_2_2_wadr;

  yt_rsc_2_3_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_2_3_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_2_3_clkr_en,
      d => yt_rsc_2_3_comp_d,
      q => yt_rsc_2_3_comp_q,
      radr => yt_rsc_2_3_comp_radr,
      wadr => yt_rsc_2_3_comp_wadr,
      we => yt_rsc_2_3_we
    );
  yt_rsc_2_3_comp_d <= yt_rsc_2_3_d;
  yt_rsc_2_3_q <= yt_rsc_2_3_comp_q;
  yt_rsc_2_3_comp_radr <= yt_rsc_2_3_radr;
  yt_rsc_2_3_comp_wadr <= yt_rsc_2_3_wadr;

  yt_rsc_2_4_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_2_4_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_2_4_clkr_en,
      d => yt_rsc_2_4_comp_d,
      q => yt_rsc_2_4_comp_q,
      radr => yt_rsc_2_4_comp_radr,
      wadr => yt_rsc_2_4_comp_wadr,
      we => yt_rsc_2_4_we
    );
  yt_rsc_2_4_comp_d <= yt_rsc_2_4_d;
  yt_rsc_2_4_q <= yt_rsc_2_4_comp_q;
  yt_rsc_2_4_comp_radr <= yt_rsc_2_4_radr;
  yt_rsc_2_4_comp_wadr <= yt_rsc_2_4_wadr;

  yt_rsc_2_5_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_2_5_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_2_5_clkr_en,
      d => yt_rsc_2_5_comp_d,
      q => yt_rsc_2_5_comp_q,
      radr => yt_rsc_2_5_comp_radr,
      wadr => yt_rsc_2_5_comp_wadr,
      we => yt_rsc_2_5_we
    );
  yt_rsc_2_5_comp_d <= yt_rsc_2_5_d;
  yt_rsc_2_5_q <= yt_rsc_2_5_comp_q;
  yt_rsc_2_5_comp_radr <= yt_rsc_2_5_radr;
  yt_rsc_2_5_comp_wadr <= yt_rsc_2_5_wadr;

  yt_rsc_2_6_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_2_6_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_2_6_clkr_en,
      d => yt_rsc_2_6_comp_d,
      q => yt_rsc_2_6_comp_q,
      radr => yt_rsc_2_6_comp_radr,
      wadr => yt_rsc_2_6_comp_wadr,
      we => yt_rsc_2_6_we
    );
  yt_rsc_2_6_comp_d <= yt_rsc_2_6_d;
  yt_rsc_2_6_q <= yt_rsc_2_6_comp_q;
  yt_rsc_2_6_comp_radr <= yt_rsc_2_6_radr;
  yt_rsc_2_6_comp_wadr <= yt_rsc_2_6_wadr;

  yt_rsc_2_7_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_2_7_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_2_7_clkr_en,
      d => yt_rsc_2_7_comp_d,
      q => yt_rsc_2_7_comp_q,
      radr => yt_rsc_2_7_comp_radr,
      wadr => yt_rsc_2_7_comp_wadr,
      we => yt_rsc_2_7_we
    );
  yt_rsc_2_7_comp_d <= yt_rsc_2_7_d;
  yt_rsc_2_7_q <= yt_rsc_2_7_comp_q;
  yt_rsc_2_7_comp_radr <= yt_rsc_2_7_radr;
  yt_rsc_2_7_comp_wadr <= yt_rsc_2_7_wadr;

  yt_rsc_2_8_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_2_8_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_2_8_clkr_en,
      d => yt_rsc_2_8_comp_d,
      q => yt_rsc_2_8_comp_q,
      radr => yt_rsc_2_8_comp_radr,
      wadr => yt_rsc_2_8_comp_wadr,
      we => yt_rsc_2_8_we
    );
  yt_rsc_2_8_comp_d <= yt_rsc_2_8_d;
  yt_rsc_2_8_q <= yt_rsc_2_8_comp_q;
  yt_rsc_2_8_comp_radr <= yt_rsc_2_8_radr;
  yt_rsc_2_8_comp_wadr <= yt_rsc_2_8_wadr;

  yt_rsc_2_9_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_2_9_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_2_9_clkr_en,
      d => yt_rsc_2_9_comp_d,
      q => yt_rsc_2_9_comp_q,
      radr => yt_rsc_2_9_comp_radr,
      wadr => yt_rsc_2_9_comp_wadr,
      we => yt_rsc_2_9_we
    );
  yt_rsc_2_9_comp_d <= yt_rsc_2_9_d;
  yt_rsc_2_9_q <= yt_rsc_2_9_comp_q;
  yt_rsc_2_9_comp_radr <= yt_rsc_2_9_radr;
  yt_rsc_2_9_comp_wadr <= yt_rsc_2_9_wadr;

  yt_rsc_2_10_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_2_10_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_2_10_clkr_en,
      d => yt_rsc_2_10_comp_d,
      q => yt_rsc_2_10_comp_q,
      radr => yt_rsc_2_10_comp_radr,
      wadr => yt_rsc_2_10_comp_wadr,
      we => yt_rsc_2_10_we
    );
  yt_rsc_2_10_comp_d <= yt_rsc_2_10_d;
  yt_rsc_2_10_q <= yt_rsc_2_10_comp_q;
  yt_rsc_2_10_comp_radr <= yt_rsc_2_10_radr;
  yt_rsc_2_10_comp_wadr <= yt_rsc_2_10_wadr;

  yt_rsc_2_11_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_2_11_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_2_11_clkr_en,
      d => yt_rsc_2_11_comp_d,
      q => yt_rsc_2_11_comp_q,
      radr => yt_rsc_2_11_comp_radr,
      wadr => yt_rsc_2_11_comp_wadr,
      we => yt_rsc_2_11_we
    );
  yt_rsc_2_11_comp_d <= yt_rsc_2_11_d;
  yt_rsc_2_11_q <= yt_rsc_2_11_comp_q;
  yt_rsc_2_11_comp_radr <= yt_rsc_2_11_radr;
  yt_rsc_2_11_comp_wadr <= yt_rsc_2_11_wadr;

  yt_rsc_2_12_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_2_12_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_2_12_clkr_en,
      d => yt_rsc_2_12_comp_d,
      q => yt_rsc_2_12_comp_q,
      radr => yt_rsc_2_12_comp_radr,
      wadr => yt_rsc_2_12_comp_wadr,
      we => yt_rsc_2_12_we
    );
  yt_rsc_2_12_comp_d <= yt_rsc_2_12_d;
  yt_rsc_2_12_q <= yt_rsc_2_12_comp_q;
  yt_rsc_2_12_comp_radr <= yt_rsc_2_12_radr;
  yt_rsc_2_12_comp_wadr <= yt_rsc_2_12_wadr;

  yt_rsc_2_13_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_2_13_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_2_13_clkr_en,
      d => yt_rsc_2_13_comp_d,
      q => yt_rsc_2_13_comp_q,
      radr => yt_rsc_2_13_comp_radr,
      wadr => yt_rsc_2_13_comp_wadr,
      we => yt_rsc_2_13_we
    );
  yt_rsc_2_13_comp_d <= yt_rsc_2_13_d;
  yt_rsc_2_13_q <= yt_rsc_2_13_comp_q;
  yt_rsc_2_13_comp_radr <= yt_rsc_2_13_radr;
  yt_rsc_2_13_comp_wadr <= yt_rsc_2_13_wadr;

  yt_rsc_2_14_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_2_14_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_2_14_clkr_en,
      d => yt_rsc_2_14_comp_d,
      q => yt_rsc_2_14_comp_q,
      radr => yt_rsc_2_14_comp_radr,
      wadr => yt_rsc_2_14_comp_wadr,
      we => yt_rsc_2_14_we
    );
  yt_rsc_2_14_comp_d <= yt_rsc_2_14_d;
  yt_rsc_2_14_q <= yt_rsc_2_14_comp_q;
  yt_rsc_2_14_comp_radr <= yt_rsc_2_14_radr;
  yt_rsc_2_14_comp_wadr <= yt_rsc_2_14_wadr;

  yt_rsc_2_15_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_2_15_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_2_15_clkr_en,
      d => yt_rsc_2_15_comp_d,
      q => yt_rsc_2_15_comp_q,
      radr => yt_rsc_2_15_comp_radr,
      wadr => yt_rsc_2_15_comp_wadr,
      we => yt_rsc_2_15_we
    );
  yt_rsc_2_15_comp_d <= yt_rsc_2_15_d;
  yt_rsc_2_15_q <= yt_rsc_2_15_comp_q;
  yt_rsc_2_15_comp_radr <= yt_rsc_2_15_radr;
  yt_rsc_2_15_comp_wadr <= yt_rsc_2_15_wadr;

  yt_rsc_2_16_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_2_16_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_2_16_clkr_en,
      d => yt_rsc_2_16_comp_d,
      q => yt_rsc_2_16_comp_q,
      radr => yt_rsc_2_16_comp_radr,
      wadr => yt_rsc_2_16_comp_wadr,
      we => yt_rsc_2_16_we
    );
  yt_rsc_2_16_comp_d <= yt_rsc_2_16_d;
  yt_rsc_2_16_q <= yt_rsc_2_16_comp_q;
  yt_rsc_2_16_comp_radr <= yt_rsc_2_16_radr;
  yt_rsc_2_16_comp_wadr <= yt_rsc_2_16_wadr;

  yt_rsc_2_17_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_2_17_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_2_17_clkr_en,
      d => yt_rsc_2_17_comp_d,
      q => yt_rsc_2_17_comp_q,
      radr => yt_rsc_2_17_comp_radr,
      wadr => yt_rsc_2_17_comp_wadr,
      we => yt_rsc_2_17_we
    );
  yt_rsc_2_17_comp_d <= yt_rsc_2_17_d;
  yt_rsc_2_17_q <= yt_rsc_2_17_comp_q;
  yt_rsc_2_17_comp_radr <= yt_rsc_2_17_radr;
  yt_rsc_2_17_comp_wadr <= yt_rsc_2_17_wadr;

  yt_rsc_2_18_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_2_18_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_2_18_clkr_en,
      d => yt_rsc_2_18_comp_d,
      q => yt_rsc_2_18_comp_q,
      radr => yt_rsc_2_18_comp_radr,
      wadr => yt_rsc_2_18_comp_wadr,
      we => yt_rsc_2_18_we
    );
  yt_rsc_2_18_comp_d <= yt_rsc_2_18_d;
  yt_rsc_2_18_q <= yt_rsc_2_18_comp_q;
  yt_rsc_2_18_comp_radr <= yt_rsc_2_18_radr;
  yt_rsc_2_18_comp_wadr <= yt_rsc_2_18_wadr;

  yt_rsc_2_19_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_2_19_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_2_19_clkr_en,
      d => yt_rsc_2_19_comp_d,
      q => yt_rsc_2_19_comp_q,
      radr => yt_rsc_2_19_comp_radr,
      wadr => yt_rsc_2_19_comp_wadr,
      we => yt_rsc_2_19_we
    );
  yt_rsc_2_19_comp_d <= yt_rsc_2_19_d;
  yt_rsc_2_19_q <= yt_rsc_2_19_comp_q;
  yt_rsc_2_19_comp_radr <= yt_rsc_2_19_radr;
  yt_rsc_2_19_comp_wadr <= yt_rsc_2_19_wadr;

  yt_rsc_2_20_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_2_20_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_2_20_clkr_en,
      d => yt_rsc_2_20_comp_d,
      q => yt_rsc_2_20_comp_q,
      radr => yt_rsc_2_20_comp_radr,
      wadr => yt_rsc_2_20_comp_wadr,
      we => yt_rsc_2_20_we
    );
  yt_rsc_2_20_comp_d <= yt_rsc_2_20_d;
  yt_rsc_2_20_q <= yt_rsc_2_20_comp_q;
  yt_rsc_2_20_comp_radr <= yt_rsc_2_20_radr;
  yt_rsc_2_20_comp_wadr <= yt_rsc_2_20_wadr;

  yt_rsc_2_21_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_2_21_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_2_21_clkr_en,
      d => yt_rsc_2_21_comp_d,
      q => yt_rsc_2_21_comp_q,
      radr => yt_rsc_2_21_comp_radr,
      wadr => yt_rsc_2_21_comp_wadr,
      we => yt_rsc_2_21_we
    );
  yt_rsc_2_21_comp_d <= yt_rsc_2_21_d;
  yt_rsc_2_21_q <= yt_rsc_2_21_comp_q;
  yt_rsc_2_21_comp_radr <= yt_rsc_2_21_radr;
  yt_rsc_2_21_comp_wadr <= yt_rsc_2_21_wadr;

  yt_rsc_2_22_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_2_22_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_2_22_clkr_en,
      d => yt_rsc_2_22_comp_d,
      q => yt_rsc_2_22_comp_q,
      radr => yt_rsc_2_22_comp_radr,
      wadr => yt_rsc_2_22_comp_wadr,
      we => yt_rsc_2_22_we
    );
  yt_rsc_2_22_comp_d <= yt_rsc_2_22_d;
  yt_rsc_2_22_q <= yt_rsc_2_22_comp_q;
  yt_rsc_2_22_comp_radr <= yt_rsc_2_22_radr;
  yt_rsc_2_22_comp_wadr <= yt_rsc_2_22_wadr;

  yt_rsc_2_23_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_2_23_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_2_23_clkr_en,
      d => yt_rsc_2_23_comp_d,
      q => yt_rsc_2_23_comp_q,
      radr => yt_rsc_2_23_comp_radr,
      wadr => yt_rsc_2_23_comp_wadr,
      we => yt_rsc_2_23_we
    );
  yt_rsc_2_23_comp_d <= yt_rsc_2_23_d;
  yt_rsc_2_23_q <= yt_rsc_2_23_comp_q;
  yt_rsc_2_23_comp_radr <= yt_rsc_2_23_radr;
  yt_rsc_2_23_comp_wadr <= yt_rsc_2_23_wadr;

  yt_rsc_2_24_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_2_24_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_2_24_clkr_en,
      d => yt_rsc_2_24_comp_d,
      q => yt_rsc_2_24_comp_q,
      radr => yt_rsc_2_24_comp_radr,
      wadr => yt_rsc_2_24_comp_wadr,
      we => yt_rsc_2_24_we
    );
  yt_rsc_2_24_comp_d <= yt_rsc_2_24_d;
  yt_rsc_2_24_q <= yt_rsc_2_24_comp_q;
  yt_rsc_2_24_comp_radr <= yt_rsc_2_24_radr;
  yt_rsc_2_24_comp_wadr <= yt_rsc_2_24_wadr;

  yt_rsc_2_25_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_2_25_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_2_25_clkr_en,
      d => yt_rsc_2_25_comp_d,
      q => yt_rsc_2_25_comp_q,
      radr => yt_rsc_2_25_comp_radr,
      wadr => yt_rsc_2_25_comp_wadr,
      we => yt_rsc_2_25_we
    );
  yt_rsc_2_25_comp_d <= yt_rsc_2_25_d;
  yt_rsc_2_25_q <= yt_rsc_2_25_comp_q;
  yt_rsc_2_25_comp_radr <= yt_rsc_2_25_radr;
  yt_rsc_2_25_comp_wadr <= yt_rsc_2_25_wadr;

  yt_rsc_2_26_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_2_26_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_2_26_clkr_en,
      d => yt_rsc_2_26_comp_d,
      q => yt_rsc_2_26_comp_q,
      radr => yt_rsc_2_26_comp_radr,
      wadr => yt_rsc_2_26_comp_wadr,
      we => yt_rsc_2_26_we
    );
  yt_rsc_2_26_comp_d <= yt_rsc_2_26_d;
  yt_rsc_2_26_q <= yt_rsc_2_26_comp_q;
  yt_rsc_2_26_comp_radr <= yt_rsc_2_26_radr;
  yt_rsc_2_26_comp_wadr <= yt_rsc_2_26_wadr;

  yt_rsc_2_27_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_2_27_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_2_27_clkr_en,
      d => yt_rsc_2_27_comp_d,
      q => yt_rsc_2_27_comp_q,
      radr => yt_rsc_2_27_comp_radr,
      wadr => yt_rsc_2_27_comp_wadr,
      we => yt_rsc_2_27_we
    );
  yt_rsc_2_27_comp_d <= yt_rsc_2_27_d;
  yt_rsc_2_27_q <= yt_rsc_2_27_comp_q;
  yt_rsc_2_27_comp_radr <= yt_rsc_2_27_radr;
  yt_rsc_2_27_comp_wadr <= yt_rsc_2_27_wadr;

  yt_rsc_2_28_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_2_28_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_2_28_clkr_en,
      d => yt_rsc_2_28_comp_d,
      q => yt_rsc_2_28_comp_q,
      radr => yt_rsc_2_28_comp_radr,
      wadr => yt_rsc_2_28_comp_wadr,
      we => yt_rsc_2_28_we
    );
  yt_rsc_2_28_comp_d <= yt_rsc_2_28_d;
  yt_rsc_2_28_q <= yt_rsc_2_28_comp_q;
  yt_rsc_2_28_comp_radr <= yt_rsc_2_28_radr;
  yt_rsc_2_28_comp_wadr <= yt_rsc_2_28_wadr;

  yt_rsc_2_29_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_2_29_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_2_29_clkr_en,
      d => yt_rsc_2_29_comp_d,
      q => yt_rsc_2_29_comp_q,
      radr => yt_rsc_2_29_comp_radr,
      wadr => yt_rsc_2_29_comp_wadr,
      we => yt_rsc_2_29_we
    );
  yt_rsc_2_29_comp_d <= yt_rsc_2_29_d;
  yt_rsc_2_29_q <= yt_rsc_2_29_comp_q;
  yt_rsc_2_29_comp_radr <= yt_rsc_2_29_radr;
  yt_rsc_2_29_comp_wadr <= yt_rsc_2_29_wadr;

  yt_rsc_2_30_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_2_30_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_2_30_clkr_en,
      d => yt_rsc_2_30_comp_d,
      q => yt_rsc_2_30_comp_q,
      radr => yt_rsc_2_30_comp_radr,
      wadr => yt_rsc_2_30_comp_wadr,
      we => yt_rsc_2_30_we
    );
  yt_rsc_2_30_comp_d <= yt_rsc_2_30_d;
  yt_rsc_2_30_q <= yt_rsc_2_30_comp_q;
  yt_rsc_2_30_comp_radr <= yt_rsc_2_30_radr;
  yt_rsc_2_30_comp_wadr <= yt_rsc_2_30_wadr;

  yt_rsc_2_31_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_2_31_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_2_31_clkr_en,
      d => yt_rsc_2_31_comp_d,
      q => yt_rsc_2_31_comp_q,
      radr => yt_rsc_2_31_comp_radr,
      wadr => yt_rsc_2_31_comp_wadr,
      we => yt_rsc_2_31_we
    );
  yt_rsc_2_31_comp_d <= yt_rsc_2_31_d;
  yt_rsc_2_31_q <= yt_rsc_2_31_comp_q;
  yt_rsc_2_31_comp_radr <= yt_rsc_2_31_radr;
  yt_rsc_2_31_comp_wadr <= yt_rsc_2_31_wadr;

  yt_rsc_3_0_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_3_0_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_3_0_clkr_en,
      d => yt_rsc_3_0_comp_d,
      q => yt_rsc_3_0_comp_q,
      radr => yt_rsc_3_0_comp_radr,
      wadr => yt_rsc_3_0_comp_wadr,
      we => yt_rsc_3_0_we
    );
  yt_rsc_3_0_comp_d <= yt_rsc_3_0_d;
  yt_rsc_3_0_q <= yt_rsc_3_0_comp_q;
  yt_rsc_3_0_comp_radr <= yt_rsc_3_0_radr;
  yt_rsc_3_0_comp_wadr <= yt_rsc_3_0_wadr;

  yt_rsc_3_1_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_3_1_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_3_1_clkr_en,
      d => yt_rsc_3_1_comp_d,
      q => yt_rsc_3_1_comp_q,
      radr => yt_rsc_3_1_comp_radr,
      wadr => yt_rsc_3_1_comp_wadr,
      we => yt_rsc_3_1_we
    );
  yt_rsc_3_1_comp_d <= yt_rsc_3_1_d;
  yt_rsc_3_1_q <= yt_rsc_3_1_comp_q;
  yt_rsc_3_1_comp_radr <= yt_rsc_3_1_radr;
  yt_rsc_3_1_comp_wadr <= yt_rsc_3_1_wadr;

  yt_rsc_3_2_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_3_2_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_3_2_clkr_en,
      d => yt_rsc_3_2_comp_d,
      q => yt_rsc_3_2_comp_q,
      radr => yt_rsc_3_2_comp_radr,
      wadr => yt_rsc_3_2_comp_wadr,
      we => yt_rsc_3_2_we
    );
  yt_rsc_3_2_comp_d <= yt_rsc_3_2_d;
  yt_rsc_3_2_q <= yt_rsc_3_2_comp_q;
  yt_rsc_3_2_comp_radr <= yt_rsc_3_2_radr;
  yt_rsc_3_2_comp_wadr <= yt_rsc_3_2_wadr;

  yt_rsc_3_3_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_3_3_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_3_3_clkr_en,
      d => yt_rsc_3_3_comp_d,
      q => yt_rsc_3_3_comp_q,
      radr => yt_rsc_3_3_comp_radr,
      wadr => yt_rsc_3_3_comp_wadr,
      we => yt_rsc_3_3_we
    );
  yt_rsc_3_3_comp_d <= yt_rsc_3_3_d;
  yt_rsc_3_3_q <= yt_rsc_3_3_comp_q;
  yt_rsc_3_3_comp_radr <= yt_rsc_3_3_radr;
  yt_rsc_3_3_comp_wadr <= yt_rsc_3_3_wadr;

  yt_rsc_3_4_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_3_4_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_3_4_clkr_en,
      d => yt_rsc_3_4_comp_d,
      q => yt_rsc_3_4_comp_q,
      radr => yt_rsc_3_4_comp_radr,
      wadr => yt_rsc_3_4_comp_wadr,
      we => yt_rsc_3_4_we
    );
  yt_rsc_3_4_comp_d <= yt_rsc_3_4_d;
  yt_rsc_3_4_q <= yt_rsc_3_4_comp_q;
  yt_rsc_3_4_comp_radr <= yt_rsc_3_4_radr;
  yt_rsc_3_4_comp_wadr <= yt_rsc_3_4_wadr;

  yt_rsc_3_5_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_3_5_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_3_5_clkr_en,
      d => yt_rsc_3_5_comp_d,
      q => yt_rsc_3_5_comp_q,
      radr => yt_rsc_3_5_comp_radr,
      wadr => yt_rsc_3_5_comp_wadr,
      we => yt_rsc_3_5_we
    );
  yt_rsc_3_5_comp_d <= yt_rsc_3_5_d;
  yt_rsc_3_5_q <= yt_rsc_3_5_comp_q;
  yt_rsc_3_5_comp_radr <= yt_rsc_3_5_radr;
  yt_rsc_3_5_comp_wadr <= yt_rsc_3_5_wadr;

  yt_rsc_3_6_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_3_6_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_3_6_clkr_en,
      d => yt_rsc_3_6_comp_d,
      q => yt_rsc_3_6_comp_q,
      radr => yt_rsc_3_6_comp_radr,
      wadr => yt_rsc_3_6_comp_wadr,
      we => yt_rsc_3_6_we
    );
  yt_rsc_3_6_comp_d <= yt_rsc_3_6_d;
  yt_rsc_3_6_q <= yt_rsc_3_6_comp_q;
  yt_rsc_3_6_comp_radr <= yt_rsc_3_6_radr;
  yt_rsc_3_6_comp_wadr <= yt_rsc_3_6_wadr;

  yt_rsc_3_7_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_3_7_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_3_7_clkr_en,
      d => yt_rsc_3_7_comp_d,
      q => yt_rsc_3_7_comp_q,
      radr => yt_rsc_3_7_comp_radr,
      wadr => yt_rsc_3_7_comp_wadr,
      we => yt_rsc_3_7_we
    );
  yt_rsc_3_7_comp_d <= yt_rsc_3_7_d;
  yt_rsc_3_7_q <= yt_rsc_3_7_comp_q;
  yt_rsc_3_7_comp_radr <= yt_rsc_3_7_radr;
  yt_rsc_3_7_comp_wadr <= yt_rsc_3_7_wadr;

  yt_rsc_3_8_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_3_8_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_3_8_clkr_en,
      d => yt_rsc_3_8_comp_d,
      q => yt_rsc_3_8_comp_q,
      radr => yt_rsc_3_8_comp_radr,
      wadr => yt_rsc_3_8_comp_wadr,
      we => yt_rsc_3_8_we
    );
  yt_rsc_3_8_comp_d <= yt_rsc_3_8_d;
  yt_rsc_3_8_q <= yt_rsc_3_8_comp_q;
  yt_rsc_3_8_comp_radr <= yt_rsc_3_8_radr;
  yt_rsc_3_8_comp_wadr <= yt_rsc_3_8_wadr;

  yt_rsc_3_9_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_3_9_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_3_9_clkr_en,
      d => yt_rsc_3_9_comp_d,
      q => yt_rsc_3_9_comp_q,
      radr => yt_rsc_3_9_comp_radr,
      wadr => yt_rsc_3_9_comp_wadr,
      we => yt_rsc_3_9_we
    );
  yt_rsc_3_9_comp_d <= yt_rsc_3_9_d;
  yt_rsc_3_9_q <= yt_rsc_3_9_comp_q;
  yt_rsc_3_9_comp_radr <= yt_rsc_3_9_radr;
  yt_rsc_3_9_comp_wadr <= yt_rsc_3_9_wadr;

  yt_rsc_3_10_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_3_10_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_3_10_clkr_en,
      d => yt_rsc_3_10_comp_d,
      q => yt_rsc_3_10_comp_q,
      radr => yt_rsc_3_10_comp_radr,
      wadr => yt_rsc_3_10_comp_wadr,
      we => yt_rsc_3_10_we
    );
  yt_rsc_3_10_comp_d <= yt_rsc_3_10_d;
  yt_rsc_3_10_q <= yt_rsc_3_10_comp_q;
  yt_rsc_3_10_comp_radr <= yt_rsc_3_10_radr;
  yt_rsc_3_10_comp_wadr <= yt_rsc_3_10_wadr;

  yt_rsc_3_11_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_3_11_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_3_11_clkr_en,
      d => yt_rsc_3_11_comp_d,
      q => yt_rsc_3_11_comp_q,
      radr => yt_rsc_3_11_comp_radr,
      wadr => yt_rsc_3_11_comp_wadr,
      we => yt_rsc_3_11_we
    );
  yt_rsc_3_11_comp_d <= yt_rsc_3_11_d;
  yt_rsc_3_11_q <= yt_rsc_3_11_comp_q;
  yt_rsc_3_11_comp_radr <= yt_rsc_3_11_radr;
  yt_rsc_3_11_comp_wadr <= yt_rsc_3_11_wadr;

  yt_rsc_3_12_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_3_12_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_3_12_clkr_en,
      d => yt_rsc_3_12_comp_d,
      q => yt_rsc_3_12_comp_q,
      radr => yt_rsc_3_12_comp_radr,
      wadr => yt_rsc_3_12_comp_wadr,
      we => yt_rsc_3_12_we
    );
  yt_rsc_3_12_comp_d <= yt_rsc_3_12_d;
  yt_rsc_3_12_q <= yt_rsc_3_12_comp_q;
  yt_rsc_3_12_comp_radr <= yt_rsc_3_12_radr;
  yt_rsc_3_12_comp_wadr <= yt_rsc_3_12_wadr;

  yt_rsc_3_13_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_3_13_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_3_13_clkr_en,
      d => yt_rsc_3_13_comp_d,
      q => yt_rsc_3_13_comp_q,
      radr => yt_rsc_3_13_comp_radr,
      wadr => yt_rsc_3_13_comp_wadr,
      we => yt_rsc_3_13_we
    );
  yt_rsc_3_13_comp_d <= yt_rsc_3_13_d;
  yt_rsc_3_13_q <= yt_rsc_3_13_comp_q;
  yt_rsc_3_13_comp_radr <= yt_rsc_3_13_radr;
  yt_rsc_3_13_comp_wadr <= yt_rsc_3_13_wadr;

  yt_rsc_3_14_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_3_14_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_3_14_clkr_en,
      d => yt_rsc_3_14_comp_d,
      q => yt_rsc_3_14_comp_q,
      radr => yt_rsc_3_14_comp_radr,
      wadr => yt_rsc_3_14_comp_wadr,
      we => yt_rsc_3_14_we
    );
  yt_rsc_3_14_comp_d <= yt_rsc_3_14_d;
  yt_rsc_3_14_q <= yt_rsc_3_14_comp_q;
  yt_rsc_3_14_comp_radr <= yt_rsc_3_14_radr;
  yt_rsc_3_14_comp_wadr <= yt_rsc_3_14_wadr;

  yt_rsc_3_15_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_3_15_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_3_15_clkr_en,
      d => yt_rsc_3_15_comp_d,
      q => yt_rsc_3_15_comp_q,
      radr => yt_rsc_3_15_comp_radr,
      wadr => yt_rsc_3_15_comp_wadr,
      we => yt_rsc_3_15_we
    );
  yt_rsc_3_15_comp_d <= yt_rsc_3_15_d;
  yt_rsc_3_15_q <= yt_rsc_3_15_comp_q;
  yt_rsc_3_15_comp_radr <= yt_rsc_3_15_radr;
  yt_rsc_3_15_comp_wadr <= yt_rsc_3_15_wadr;

  yt_rsc_3_16_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_3_16_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_3_16_clkr_en,
      d => yt_rsc_3_16_comp_d,
      q => yt_rsc_3_16_comp_q,
      radr => yt_rsc_3_16_comp_radr,
      wadr => yt_rsc_3_16_comp_wadr,
      we => yt_rsc_3_16_we
    );
  yt_rsc_3_16_comp_d <= yt_rsc_3_16_d;
  yt_rsc_3_16_q <= yt_rsc_3_16_comp_q;
  yt_rsc_3_16_comp_radr <= yt_rsc_3_16_radr;
  yt_rsc_3_16_comp_wadr <= yt_rsc_3_16_wadr;

  yt_rsc_3_17_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_3_17_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_3_17_clkr_en,
      d => yt_rsc_3_17_comp_d,
      q => yt_rsc_3_17_comp_q,
      radr => yt_rsc_3_17_comp_radr,
      wadr => yt_rsc_3_17_comp_wadr,
      we => yt_rsc_3_17_we
    );
  yt_rsc_3_17_comp_d <= yt_rsc_3_17_d;
  yt_rsc_3_17_q <= yt_rsc_3_17_comp_q;
  yt_rsc_3_17_comp_radr <= yt_rsc_3_17_radr;
  yt_rsc_3_17_comp_wadr <= yt_rsc_3_17_wadr;

  yt_rsc_3_18_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_3_18_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_3_18_clkr_en,
      d => yt_rsc_3_18_comp_d,
      q => yt_rsc_3_18_comp_q,
      radr => yt_rsc_3_18_comp_radr,
      wadr => yt_rsc_3_18_comp_wadr,
      we => yt_rsc_3_18_we
    );
  yt_rsc_3_18_comp_d <= yt_rsc_3_18_d;
  yt_rsc_3_18_q <= yt_rsc_3_18_comp_q;
  yt_rsc_3_18_comp_radr <= yt_rsc_3_18_radr;
  yt_rsc_3_18_comp_wadr <= yt_rsc_3_18_wadr;

  yt_rsc_3_19_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_3_19_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_3_19_clkr_en,
      d => yt_rsc_3_19_comp_d,
      q => yt_rsc_3_19_comp_q,
      radr => yt_rsc_3_19_comp_radr,
      wadr => yt_rsc_3_19_comp_wadr,
      we => yt_rsc_3_19_we
    );
  yt_rsc_3_19_comp_d <= yt_rsc_3_19_d;
  yt_rsc_3_19_q <= yt_rsc_3_19_comp_q;
  yt_rsc_3_19_comp_radr <= yt_rsc_3_19_radr;
  yt_rsc_3_19_comp_wadr <= yt_rsc_3_19_wadr;

  yt_rsc_3_20_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_3_20_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_3_20_clkr_en,
      d => yt_rsc_3_20_comp_d,
      q => yt_rsc_3_20_comp_q,
      radr => yt_rsc_3_20_comp_radr,
      wadr => yt_rsc_3_20_comp_wadr,
      we => yt_rsc_3_20_we
    );
  yt_rsc_3_20_comp_d <= yt_rsc_3_20_d;
  yt_rsc_3_20_q <= yt_rsc_3_20_comp_q;
  yt_rsc_3_20_comp_radr <= yt_rsc_3_20_radr;
  yt_rsc_3_20_comp_wadr <= yt_rsc_3_20_wadr;

  yt_rsc_3_21_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_3_21_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_3_21_clkr_en,
      d => yt_rsc_3_21_comp_d,
      q => yt_rsc_3_21_comp_q,
      radr => yt_rsc_3_21_comp_radr,
      wadr => yt_rsc_3_21_comp_wadr,
      we => yt_rsc_3_21_we
    );
  yt_rsc_3_21_comp_d <= yt_rsc_3_21_d;
  yt_rsc_3_21_q <= yt_rsc_3_21_comp_q;
  yt_rsc_3_21_comp_radr <= yt_rsc_3_21_radr;
  yt_rsc_3_21_comp_wadr <= yt_rsc_3_21_wadr;

  yt_rsc_3_22_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_3_22_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_3_22_clkr_en,
      d => yt_rsc_3_22_comp_d,
      q => yt_rsc_3_22_comp_q,
      radr => yt_rsc_3_22_comp_radr,
      wadr => yt_rsc_3_22_comp_wadr,
      we => yt_rsc_3_22_we
    );
  yt_rsc_3_22_comp_d <= yt_rsc_3_22_d;
  yt_rsc_3_22_q <= yt_rsc_3_22_comp_q;
  yt_rsc_3_22_comp_radr <= yt_rsc_3_22_radr;
  yt_rsc_3_22_comp_wadr <= yt_rsc_3_22_wadr;

  yt_rsc_3_23_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_3_23_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_3_23_clkr_en,
      d => yt_rsc_3_23_comp_d,
      q => yt_rsc_3_23_comp_q,
      radr => yt_rsc_3_23_comp_radr,
      wadr => yt_rsc_3_23_comp_wadr,
      we => yt_rsc_3_23_we
    );
  yt_rsc_3_23_comp_d <= yt_rsc_3_23_d;
  yt_rsc_3_23_q <= yt_rsc_3_23_comp_q;
  yt_rsc_3_23_comp_radr <= yt_rsc_3_23_radr;
  yt_rsc_3_23_comp_wadr <= yt_rsc_3_23_wadr;

  yt_rsc_3_24_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_3_24_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_3_24_clkr_en,
      d => yt_rsc_3_24_comp_d,
      q => yt_rsc_3_24_comp_q,
      radr => yt_rsc_3_24_comp_radr,
      wadr => yt_rsc_3_24_comp_wadr,
      we => yt_rsc_3_24_we
    );
  yt_rsc_3_24_comp_d <= yt_rsc_3_24_d;
  yt_rsc_3_24_q <= yt_rsc_3_24_comp_q;
  yt_rsc_3_24_comp_radr <= yt_rsc_3_24_radr;
  yt_rsc_3_24_comp_wadr <= yt_rsc_3_24_wadr;

  yt_rsc_3_25_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_3_25_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_3_25_clkr_en,
      d => yt_rsc_3_25_comp_d,
      q => yt_rsc_3_25_comp_q,
      radr => yt_rsc_3_25_comp_radr,
      wadr => yt_rsc_3_25_comp_wadr,
      we => yt_rsc_3_25_we
    );
  yt_rsc_3_25_comp_d <= yt_rsc_3_25_d;
  yt_rsc_3_25_q <= yt_rsc_3_25_comp_q;
  yt_rsc_3_25_comp_radr <= yt_rsc_3_25_radr;
  yt_rsc_3_25_comp_wadr <= yt_rsc_3_25_wadr;

  yt_rsc_3_26_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_3_26_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_3_26_clkr_en,
      d => yt_rsc_3_26_comp_d,
      q => yt_rsc_3_26_comp_q,
      radr => yt_rsc_3_26_comp_radr,
      wadr => yt_rsc_3_26_comp_wadr,
      we => yt_rsc_3_26_we
    );
  yt_rsc_3_26_comp_d <= yt_rsc_3_26_d;
  yt_rsc_3_26_q <= yt_rsc_3_26_comp_q;
  yt_rsc_3_26_comp_radr <= yt_rsc_3_26_radr;
  yt_rsc_3_26_comp_wadr <= yt_rsc_3_26_wadr;

  yt_rsc_3_27_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_3_27_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_3_27_clkr_en,
      d => yt_rsc_3_27_comp_d,
      q => yt_rsc_3_27_comp_q,
      radr => yt_rsc_3_27_comp_radr,
      wadr => yt_rsc_3_27_comp_wadr,
      we => yt_rsc_3_27_we
    );
  yt_rsc_3_27_comp_d <= yt_rsc_3_27_d;
  yt_rsc_3_27_q <= yt_rsc_3_27_comp_q;
  yt_rsc_3_27_comp_radr <= yt_rsc_3_27_radr;
  yt_rsc_3_27_comp_wadr <= yt_rsc_3_27_wadr;

  yt_rsc_3_28_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_3_28_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_3_28_clkr_en,
      d => yt_rsc_3_28_comp_d,
      q => yt_rsc_3_28_comp_q,
      radr => yt_rsc_3_28_comp_radr,
      wadr => yt_rsc_3_28_comp_wadr,
      we => yt_rsc_3_28_we
    );
  yt_rsc_3_28_comp_d <= yt_rsc_3_28_d;
  yt_rsc_3_28_q <= yt_rsc_3_28_comp_q;
  yt_rsc_3_28_comp_radr <= yt_rsc_3_28_radr;
  yt_rsc_3_28_comp_wadr <= yt_rsc_3_28_wadr;

  yt_rsc_3_29_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_3_29_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_3_29_clkr_en,
      d => yt_rsc_3_29_comp_d,
      q => yt_rsc_3_29_comp_q,
      radr => yt_rsc_3_29_comp_radr,
      wadr => yt_rsc_3_29_comp_wadr,
      we => yt_rsc_3_29_we
    );
  yt_rsc_3_29_comp_d <= yt_rsc_3_29_d;
  yt_rsc_3_29_q <= yt_rsc_3_29_comp_q;
  yt_rsc_3_29_comp_radr <= yt_rsc_3_29_radr;
  yt_rsc_3_29_comp_wadr <= yt_rsc_3_29_wadr;

  yt_rsc_3_30_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_3_30_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_3_30_clkr_en,
      d => yt_rsc_3_30_comp_d,
      q => yt_rsc_3_30_comp_q,
      radr => yt_rsc_3_30_comp_radr,
      wadr => yt_rsc_3_30_comp_wadr,
      we => yt_rsc_3_30_we
    );
  yt_rsc_3_30_comp_d <= yt_rsc_3_30_d;
  yt_rsc_3_30_q <= yt_rsc_3_30_comp_q;
  yt_rsc_3_30_comp_radr <= yt_rsc_3_30_radr;
  yt_rsc_3_30_comp_wadr <= yt_rsc_3_30_wadr;

  yt_rsc_3_31_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_3_31_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_3_31_clkr_en,
      d => yt_rsc_3_31_comp_d,
      q => yt_rsc_3_31_comp_q,
      radr => yt_rsc_3_31_comp_radr,
      wadr => yt_rsc_3_31_comp_wadr,
      we => yt_rsc_3_31_we
    );
  yt_rsc_3_31_comp_d <= yt_rsc_3_31_d;
  yt_rsc_3_31_q <= yt_rsc_3_31_comp_q;
  yt_rsc_3_31_comp_radr <= yt_rsc_3_31_radr;
  yt_rsc_3_31_comp_wadr <= yt_rsc_3_31_wadr;

  yt_rsc_4_0_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_4_0_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_4_0_clkr_en,
      d => yt_rsc_4_0_comp_d,
      q => yt_rsc_4_0_comp_q,
      radr => yt_rsc_4_0_comp_radr,
      wadr => yt_rsc_4_0_comp_wadr,
      we => yt_rsc_4_0_we
    );
  yt_rsc_4_0_comp_d <= yt_rsc_4_0_d;
  yt_rsc_4_0_q <= yt_rsc_4_0_comp_q;
  yt_rsc_4_0_comp_radr <= yt_rsc_4_0_radr;
  yt_rsc_4_0_comp_wadr <= yt_rsc_4_0_wadr;

  yt_rsc_4_1_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_4_1_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_4_1_clkr_en,
      d => yt_rsc_4_1_comp_d,
      q => yt_rsc_4_1_comp_q,
      radr => yt_rsc_4_1_comp_radr,
      wadr => yt_rsc_4_1_comp_wadr,
      we => yt_rsc_4_1_we
    );
  yt_rsc_4_1_comp_d <= yt_rsc_4_1_d;
  yt_rsc_4_1_q <= yt_rsc_4_1_comp_q;
  yt_rsc_4_1_comp_radr <= yt_rsc_4_1_radr;
  yt_rsc_4_1_comp_wadr <= yt_rsc_4_1_wadr;

  yt_rsc_4_2_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_4_2_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_4_2_clkr_en,
      d => yt_rsc_4_2_comp_d,
      q => yt_rsc_4_2_comp_q,
      radr => yt_rsc_4_2_comp_radr,
      wadr => yt_rsc_4_2_comp_wadr,
      we => yt_rsc_4_2_we
    );
  yt_rsc_4_2_comp_d <= yt_rsc_4_2_d;
  yt_rsc_4_2_q <= yt_rsc_4_2_comp_q;
  yt_rsc_4_2_comp_radr <= yt_rsc_4_2_radr;
  yt_rsc_4_2_comp_wadr <= yt_rsc_4_2_wadr;

  yt_rsc_4_3_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_4_3_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_4_3_clkr_en,
      d => yt_rsc_4_3_comp_d,
      q => yt_rsc_4_3_comp_q,
      radr => yt_rsc_4_3_comp_radr,
      wadr => yt_rsc_4_3_comp_wadr,
      we => yt_rsc_4_3_we
    );
  yt_rsc_4_3_comp_d <= yt_rsc_4_3_d;
  yt_rsc_4_3_q <= yt_rsc_4_3_comp_q;
  yt_rsc_4_3_comp_radr <= yt_rsc_4_3_radr;
  yt_rsc_4_3_comp_wadr <= yt_rsc_4_3_wadr;

  yt_rsc_4_4_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_4_4_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_4_4_clkr_en,
      d => yt_rsc_4_4_comp_d,
      q => yt_rsc_4_4_comp_q,
      radr => yt_rsc_4_4_comp_radr,
      wadr => yt_rsc_4_4_comp_wadr,
      we => yt_rsc_4_4_we
    );
  yt_rsc_4_4_comp_d <= yt_rsc_4_4_d;
  yt_rsc_4_4_q <= yt_rsc_4_4_comp_q;
  yt_rsc_4_4_comp_radr <= yt_rsc_4_4_radr;
  yt_rsc_4_4_comp_wadr <= yt_rsc_4_4_wadr;

  yt_rsc_4_5_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_4_5_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_4_5_clkr_en,
      d => yt_rsc_4_5_comp_d,
      q => yt_rsc_4_5_comp_q,
      radr => yt_rsc_4_5_comp_radr,
      wadr => yt_rsc_4_5_comp_wadr,
      we => yt_rsc_4_5_we
    );
  yt_rsc_4_5_comp_d <= yt_rsc_4_5_d;
  yt_rsc_4_5_q <= yt_rsc_4_5_comp_q;
  yt_rsc_4_5_comp_radr <= yt_rsc_4_5_radr;
  yt_rsc_4_5_comp_wadr <= yt_rsc_4_5_wadr;

  yt_rsc_4_6_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_4_6_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_4_6_clkr_en,
      d => yt_rsc_4_6_comp_d,
      q => yt_rsc_4_6_comp_q,
      radr => yt_rsc_4_6_comp_radr,
      wadr => yt_rsc_4_6_comp_wadr,
      we => yt_rsc_4_6_we
    );
  yt_rsc_4_6_comp_d <= yt_rsc_4_6_d;
  yt_rsc_4_6_q <= yt_rsc_4_6_comp_q;
  yt_rsc_4_6_comp_radr <= yt_rsc_4_6_radr;
  yt_rsc_4_6_comp_wadr <= yt_rsc_4_6_wadr;

  yt_rsc_4_7_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_4_7_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_4_7_clkr_en,
      d => yt_rsc_4_7_comp_d,
      q => yt_rsc_4_7_comp_q,
      radr => yt_rsc_4_7_comp_radr,
      wadr => yt_rsc_4_7_comp_wadr,
      we => yt_rsc_4_7_we
    );
  yt_rsc_4_7_comp_d <= yt_rsc_4_7_d;
  yt_rsc_4_7_q <= yt_rsc_4_7_comp_q;
  yt_rsc_4_7_comp_radr <= yt_rsc_4_7_radr;
  yt_rsc_4_7_comp_wadr <= yt_rsc_4_7_wadr;

  yt_rsc_4_8_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_4_8_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_4_8_clkr_en,
      d => yt_rsc_4_8_comp_d,
      q => yt_rsc_4_8_comp_q,
      radr => yt_rsc_4_8_comp_radr,
      wadr => yt_rsc_4_8_comp_wadr,
      we => yt_rsc_4_8_we
    );
  yt_rsc_4_8_comp_d <= yt_rsc_4_8_d;
  yt_rsc_4_8_q <= yt_rsc_4_8_comp_q;
  yt_rsc_4_8_comp_radr <= yt_rsc_4_8_radr;
  yt_rsc_4_8_comp_wadr <= yt_rsc_4_8_wadr;

  yt_rsc_4_9_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_4_9_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_4_9_clkr_en,
      d => yt_rsc_4_9_comp_d,
      q => yt_rsc_4_9_comp_q,
      radr => yt_rsc_4_9_comp_radr,
      wadr => yt_rsc_4_9_comp_wadr,
      we => yt_rsc_4_9_we
    );
  yt_rsc_4_9_comp_d <= yt_rsc_4_9_d;
  yt_rsc_4_9_q <= yt_rsc_4_9_comp_q;
  yt_rsc_4_9_comp_radr <= yt_rsc_4_9_radr;
  yt_rsc_4_9_comp_wadr <= yt_rsc_4_9_wadr;

  yt_rsc_4_10_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_4_10_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_4_10_clkr_en,
      d => yt_rsc_4_10_comp_d,
      q => yt_rsc_4_10_comp_q,
      radr => yt_rsc_4_10_comp_radr,
      wadr => yt_rsc_4_10_comp_wadr,
      we => yt_rsc_4_10_we
    );
  yt_rsc_4_10_comp_d <= yt_rsc_4_10_d;
  yt_rsc_4_10_q <= yt_rsc_4_10_comp_q;
  yt_rsc_4_10_comp_radr <= yt_rsc_4_10_radr;
  yt_rsc_4_10_comp_wadr <= yt_rsc_4_10_wadr;

  yt_rsc_4_11_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_4_11_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_4_11_clkr_en,
      d => yt_rsc_4_11_comp_d,
      q => yt_rsc_4_11_comp_q,
      radr => yt_rsc_4_11_comp_radr,
      wadr => yt_rsc_4_11_comp_wadr,
      we => yt_rsc_4_11_we
    );
  yt_rsc_4_11_comp_d <= yt_rsc_4_11_d;
  yt_rsc_4_11_q <= yt_rsc_4_11_comp_q;
  yt_rsc_4_11_comp_radr <= yt_rsc_4_11_radr;
  yt_rsc_4_11_comp_wadr <= yt_rsc_4_11_wadr;

  yt_rsc_4_12_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_4_12_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_4_12_clkr_en,
      d => yt_rsc_4_12_comp_d,
      q => yt_rsc_4_12_comp_q,
      radr => yt_rsc_4_12_comp_radr,
      wadr => yt_rsc_4_12_comp_wadr,
      we => yt_rsc_4_12_we
    );
  yt_rsc_4_12_comp_d <= yt_rsc_4_12_d;
  yt_rsc_4_12_q <= yt_rsc_4_12_comp_q;
  yt_rsc_4_12_comp_radr <= yt_rsc_4_12_radr;
  yt_rsc_4_12_comp_wadr <= yt_rsc_4_12_wadr;

  yt_rsc_4_13_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_4_13_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_4_13_clkr_en,
      d => yt_rsc_4_13_comp_d,
      q => yt_rsc_4_13_comp_q,
      radr => yt_rsc_4_13_comp_radr,
      wadr => yt_rsc_4_13_comp_wadr,
      we => yt_rsc_4_13_we
    );
  yt_rsc_4_13_comp_d <= yt_rsc_4_13_d;
  yt_rsc_4_13_q <= yt_rsc_4_13_comp_q;
  yt_rsc_4_13_comp_radr <= yt_rsc_4_13_radr;
  yt_rsc_4_13_comp_wadr <= yt_rsc_4_13_wadr;

  yt_rsc_4_14_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_4_14_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_4_14_clkr_en,
      d => yt_rsc_4_14_comp_d,
      q => yt_rsc_4_14_comp_q,
      radr => yt_rsc_4_14_comp_radr,
      wadr => yt_rsc_4_14_comp_wadr,
      we => yt_rsc_4_14_we
    );
  yt_rsc_4_14_comp_d <= yt_rsc_4_14_d;
  yt_rsc_4_14_q <= yt_rsc_4_14_comp_q;
  yt_rsc_4_14_comp_radr <= yt_rsc_4_14_radr;
  yt_rsc_4_14_comp_wadr <= yt_rsc_4_14_wadr;

  yt_rsc_4_15_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_4_15_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_4_15_clkr_en,
      d => yt_rsc_4_15_comp_d,
      q => yt_rsc_4_15_comp_q,
      radr => yt_rsc_4_15_comp_radr,
      wadr => yt_rsc_4_15_comp_wadr,
      we => yt_rsc_4_15_we
    );
  yt_rsc_4_15_comp_d <= yt_rsc_4_15_d;
  yt_rsc_4_15_q <= yt_rsc_4_15_comp_q;
  yt_rsc_4_15_comp_radr <= yt_rsc_4_15_radr;
  yt_rsc_4_15_comp_wadr <= yt_rsc_4_15_wadr;

  yt_rsc_4_16_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_4_16_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_4_16_clkr_en,
      d => yt_rsc_4_16_comp_d,
      q => yt_rsc_4_16_comp_q,
      radr => yt_rsc_4_16_comp_radr,
      wadr => yt_rsc_4_16_comp_wadr,
      we => yt_rsc_4_16_we
    );
  yt_rsc_4_16_comp_d <= yt_rsc_4_16_d;
  yt_rsc_4_16_q <= yt_rsc_4_16_comp_q;
  yt_rsc_4_16_comp_radr <= yt_rsc_4_16_radr;
  yt_rsc_4_16_comp_wadr <= yt_rsc_4_16_wadr;

  yt_rsc_4_17_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_4_17_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_4_17_clkr_en,
      d => yt_rsc_4_17_comp_d,
      q => yt_rsc_4_17_comp_q,
      radr => yt_rsc_4_17_comp_radr,
      wadr => yt_rsc_4_17_comp_wadr,
      we => yt_rsc_4_17_we
    );
  yt_rsc_4_17_comp_d <= yt_rsc_4_17_d;
  yt_rsc_4_17_q <= yt_rsc_4_17_comp_q;
  yt_rsc_4_17_comp_radr <= yt_rsc_4_17_radr;
  yt_rsc_4_17_comp_wadr <= yt_rsc_4_17_wadr;

  yt_rsc_4_18_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_4_18_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_4_18_clkr_en,
      d => yt_rsc_4_18_comp_d,
      q => yt_rsc_4_18_comp_q,
      radr => yt_rsc_4_18_comp_radr,
      wadr => yt_rsc_4_18_comp_wadr,
      we => yt_rsc_4_18_we
    );
  yt_rsc_4_18_comp_d <= yt_rsc_4_18_d;
  yt_rsc_4_18_q <= yt_rsc_4_18_comp_q;
  yt_rsc_4_18_comp_radr <= yt_rsc_4_18_radr;
  yt_rsc_4_18_comp_wadr <= yt_rsc_4_18_wadr;

  yt_rsc_4_19_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_4_19_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_4_19_clkr_en,
      d => yt_rsc_4_19_comp_d,
      q => yt_rsc_4_19_comp_q,
      radr => yt_rsc_4_19_comp_radr,
      wadr => yt_rsc_4_19_comp_wadr,
      we => yt_rsc_4_19_we
    );
  yt_rsc_4_19_comp_d <= yt_rsc_4_19_d;
  yt_rsc_4_19_q <= yt_rsc_4_19_comp_q;
  yt_rsc_4_19_comp_radr <= yt_rsc_4_19_radr;
  yt_rsc_4_19_comp_wadr <= yt_rsc_4_19_wadr;

  yt_rsc_4_20_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_4_20_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_4_20_clkr_en,
      d => yt_rsc_4_20_comp_d,
      q => yt_rsc_4_20_comp_q,
      radr => yt_rsc_4_20_comp_radr,
      wadr => yt_rsc_4_20_comp_wadr,
      we => yt_rsc_4_20_we
    );
  yt_rsc_4_20_comp_d <= yt_rsc_4_20_d;
  yt_rsc_4_20_q <= yt_rsc_4_20_comp_q;
  yt_rsc_4_20_comp_radr <= yt_rsc_4_20_radr;
  yt_rsc_4_20_comp_wadr <= yt_rsc_4_20_wadr;

  yt_rsc_4_21_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_4_21_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_4_21_clkr_en,
      d => yt_rsc_4_21_comp_d,
      q => yt_rsc_4_21_comp_q,
      radr => yt_rsc_4_21_comp_radr,
      wadr => yt_rsc_4_21_comp_wadr,
      we => yt_rsc_4_21_we
    );
  yt_rsc_4_21_comp_d <= yt_rsc_4_21_d;
  yt_rsc_4_21_q <= yt_rsc_4_21_comp_q;
  yt_rsc_4_21_comp_radr <= yt_rsc_4_21_radr;
  yt_rsc_4_21_comp_wadr <= yt_rsc_4_21_wadr;

  yt_rsc_4_22_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_4_22_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_4_22_clkr_en,
      d => yt_rsc_4_22_comp_d,
      q => yt_rsc_4_22_comp_q,
      radr => yt_rsc_4_22_comp_radr,
      wadr => yt_rsc_4_22_comp_wadr,
      we => yt_rsc_4_22_we
    );
  yt_rsc_4_22_comp_d <= yt_rsc_4_22_d;
  yt_rsc_4_22_q <= yt_rsc_4_22_comp_q;
  yt_rsc_4_22_comp_radr <= yt_rsc_4_22_radr;
  yt_rsc_4_22_comp_wadr <= yt_rsc_4_22_wadr;

  yt_rsc_4_23_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_4_23_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_4_23_clkr_en,
      d => yt_rsc_4_23_comp_d,
      q => yt_rsc_4_23_comp_q,
      radr => yt_rsc_4_23_comp_radr,
      wadr => yt_rsc_4_23_comp_wadr,
      we => yt_rsc_4_23_we
    );
  yt_rsc_4_23_comp_d <= yt_rsc_4_23_d;
  yt_rsc_4_23_q <= yt_rsc_4_23_comp_q;
  yt_rsc_4_23_comp_radr <= yt_rsc_4_23_radr;
  yt_rsc_4_23_comp_wadr <= yt_rsc_4_23_wadr;

  yt_rsc_4_24_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_4_24_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_4_24_clkr_en,
      d => yt_rsc_4_24_comp_d,
      q => yt_rsc_4_24_comp_q,
      radr => yt_rsc_4_24_comp_radr,
      wadr => yt_rsc_4_24_comp_wadr,
      we => yt_rsc_4_24_we
    );
  yt_rsc_4_24_comp_d <= yt_rsc_4_24_d;
  yt_rsc_4_24_q <= yt_rsc_4_24_comp_q;
  yt_rsc_4_24_comp_radr <= yt_rsc_4_24_radr;
  yt_rsc_4_24_comp_wadr <= yt_rsc_4_24_wadr;

  yt_rsc_4_25_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_4_25_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_4_25_clkr_en,
      d => yt_rsc_4_25_comp_d,
      q => yt_rsc_4_25_comp_q,
      radr => yt_rsc_4_25_comp_radr,
      wadr => yt_rsc_4_25_comp_wadr,
      we => yt_rsc_4_25_we
    );
  yt_rsc_4_25_comp_d <= yt_rsc_4_25_d;
  yt_rsc_4_25_q <= yt_rsc_4_25_comp_q;
  yt_rsc_4_25_comp_radr <= yt_rsc_4_25_radr;
  yt_rsc_4_25_comp_wadr <= yt_rsc_4_25_wadr;

  yt_rsc_4_26_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_4_26_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_4_26_clkr_en,
      d => yt_rsc_4_26_comp_d,
      q => yt_rsc_4_26_comp_q,
      radr => yt_rsc_4_26_comp_radr,
      wadr => yt_rsc_4_26_comp_wadr,
      we => yt_rsc_4_26_we
    );
  yt_rsc_4_26_comp_d <= yt_rsc_4_26_d;
  yt_rsc_4_26_q <= yt_rsc_4_26_comp_q;
  yt_rsc_4_26_comp_radr <= yt_rsc_4_26_radr;
  yt_rsc_4_26_comp_wadr <= yt_rsc_4_26_wadr;

  yt_rsc_4_27_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_4_27_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_4_27_clkr_en,
      d => yt_rsc_4_27_comp_d,
      q => yt_rsc_4_27_comp_q,
      radr => yt_rsc_4_27_comp_radr,
      wadr => yt_rsc_4_27_comp_wadr,
      we => yt_rsc_4_27_we
    );
  yt_rsc_4_27_comp_d <= yt_rsc_4_27_d;
  yt_rsc_4_27_q <= yt_rsc_4_27_comp_q;
  yt_rsc_4_27_comp_radr <= yt_rsc_4_27_radr;
  yt_rsc_4_27_comp_wadr <= yt_rsc_4_27_wadr;

  yt_rsc_4_28_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_4_28_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_4_28_clkr_en,
      d => yt_rsc_4_28_comp_d,
      q => yt_rsc_4_28_comp_q,
      radr => yt_rsc_4_28_comp_radr,
      wadr => yt_rsc_4_28_comp_wadr,
      we => yt_rsc_4_28_we
    );
  yt_rsc_4_28_comp_d <= yt_rsc_4_28_d;
  yt_rsc_4_28_q <= yt_rsc_4_28_comp_q;
  yt_rsc_4_28_comp_radr <= yt_rsc_4_28_radr;
  yt_rsc_4_28_comp_wadr <= yt_rsc_4_28_wadr;

  yt_rsc_4_29_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_4_29_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_4_29_clkr_en,
      d => yt_rsc_4_29_comp_d,
      q => yt_rsc_4_29_comp_q,
      radr => yt_rsc_4_29_comp_radr,
      wadr => yt_rsc_4_29_comp_wadr,
      we => yt_rsc_4_29_we
    );
  yt_rsc_4_29_comp_d <= yt_rsc_4_29_d;
  yt_rsc_4_29_q <= yt_rsc_4_29_comp_q;
  yt_rsc_4_29_comp_radr <= yt_rsc_4_29_radr;
  yt_rsc_4_29_comp_wadr <= yt_rsc_4_29_wadr;

  yt_rsc_4_30_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_4_30_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_4_30_clkr_en,
      d => yt_rsc_4_30_comp_d,
      q => yt_rsc_4_30_comp_q,
      radr => yt_rsc_4_30_comp_radr,
      wadr => yt_rsc_4_30_comp_wadr,
      we => yt_rsc_4_30_we
    );
  yt_rsc_4_30_comp_d <= yt_rsc_4_30_d;
  yt_rsc_4_30_q <= yt_rsc_4_30_comp_q;
  yt_rsc_4_30_comp_radr <= yt_rsc_4_30_radr;
  yt_rsc_4_30_comp_wadr <= yt_rsc_4_30_wadr;

  yt_rsc_4_31_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_4_31_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_4_31_clkr_en,
      d => yt_rsc_4_31_comp_d,
      q => yt_rsc_4_31_comp_q,
      radr => yt_rsc_4_31_comp_radr,
      wadr => yt_rsc_4_31_comp_wadr,
      we => yt_rsc_4_31_we
    );
  yt_rsc_4_31_comp_d <= yt_rsc_4_31_d;
  yt_rsc_4_31_q <= yt_rsc_4_31_comp_q;
  yt_rsc_4_31_comp_radr <= yt_rsc_4_31_radr;
  yt_rsc_4_31_comp_wadr <= yt_rsc_4_31_wadr;

  yt_rsc_5_0_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_5_0_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_5_0_clkr_en,
      d => yt_rsc_5_0_comp_d,
      q => yt_rsc_5_0_comp_q,
      radr => yt_rsc_5_0_comp_radr,
      wadr => yt_rsc_5_0_comp_wadr,
      we => yt_rsc_5_0_we
    );
  yt_rsc_5_0_comp_d <= yt_rsc_5_0_d;
  yt_rsc_5_0_q <= yt_rsc_5_0_comp_q;
  yt_rsc_5_0_comp_radr <= yt_rsc_5_0_radr;
  yt_rsc_5_0_comp_wadr <= yt_rsc_5_0_wadr;

  yt_rsc_5_1_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_5_1_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_5_1_clkr_en,
      d => yt_rsc_5_1_comp_d,
      q => yt_rsc_5_1_comp_q,
      radr => yt_rsc_5_1_comp_radr,
      wadr => yt_rsc_5_1_comp_wadr,
      we => yt_rsc_5_1_we
    );
  yt_rsc_5_1_comp_d <= yt_rsc_5_1_d;
  yt_rsc_5_1_q <= yt_rsc_5_1_comp_q;
  yt_rsc_5_1_comp_radr <= yt_rsc_5_1_radr;
  yt_rsc_5_1_comp_wadr <= yt_rsc_5_1_wadr;

  yt_rsc_5_2_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_5_2_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_5_2_clkr_en,
      d => yt_rsc_5_2_comp_d,
      q => yt_rsc_5_2_comp_q,
      radr => yt_rsc_5_2_comp_radr,
      wadr => yt_rsc_5_2_comp_wadr,
      we => yt_rsc_5_2_we
    );
  yt_rsc_5_2_comp_d <= yt_rsc_5_2_d;
  yt_rsc_5_2_q <= yt_rsc_5_2_comp_q;
  yt_rsc_5_2_comp_radr <= yt_rsc_5_2_radr;
  yt_rsc_5_2_comp_wadr <= yt_rsc_5_2_wadr;

  yt_rsc_5_3_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_5_3_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_5_3_clkr_en,
      d => yt_rsc_5_3_comp_d,
      q => yt_rsc_5_3_comp_q,
      radr => yt_rsc_5_3_comp_radr,
      wadr => yt_rsc_5_3_comp_wadr,
      we => yt_rsc_5_3_we
    );
  yt_rsc_5_3_comp_d <= yt_rsc_5_3_d;
  yt_rsc_5_3_q <= yt_rsc_5_3_comp_q;
  yt_rsc_5_3_comp_radr <= yt_rsc_5_3_radr;
  yt_rsc_5_3_comp_wadr <= yt_rsc_5_3_wadr;

  yt_rsc_5_4_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_5_4_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_5_4_clkr_en,
      d => yt_rsc_5_4_comp_d,
      q => yt_rsc_5_4_comp_q,
      radr => yt_rsc_5_4_comp_radr,
      wadr => yt_rsc_5_4_comp_wadr,
      we => yt_rsc_5_4_we
    );
  yt_rsc_5_4_comp_d <= yt_rsc_5_4_d;
  yt_rsc_5_4_q <= yt_rsc_5_4_comp_q;
  yt_rsc_5_4_comp_radr <= yt_rsc_5_4_radr;
  yt_rsc_5_4_comp_wadr <= yt_rsc_5_4_wadr;

  yt_rsc_5_5_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_5_5_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_5_5_clkr_en,
      d => yt_rsc_5_5_comp_d,
      q => yt_rsc_5_5_comp_q,
      radr => yt_rsc_5_5_comp_radr,
      wadr => yt_rsc_5_5_comp_wadr,
      we => yt_rsc_5_5_we
    );
  yt_rsc_5_5_comp_d <= yt_rsc_5_5_d;
  yt_rsc_5_5_q <= yt_rsc_5_5_comp_q;
  yt_rsc_5_5_comp_radr <= yt_rsc_5_5_radr;
  yt_rsc_5_5_comp_wadr <= yt_rsc_5_5_wadr;

  yt_rsc_5_6_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_5_6_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_5_6_clkr_en,
      d => yt_rsc_5_6_comp_d,
      q => yt_rsc_5_6_comp_q,
      radr => yt_rsc_5_6_comp_radr,
      wadr => yt_rsc_5_6_comp_wadr,
      we => yt_rsc_5_6_we
    );
  yt_rsc_5_6_comp_d <= yt_rsc_5_6_d;
  yt_rsc_5_6_q <= yt_rsc_5_6_comp_q;
  yt_rsc_5_6_comp_radr <= yt_rsc_5_6_radr;
  yt_rsc_5_6_comp_wadr <= yt_rsc_5_6_wadr;

  yt_rsc_5_7_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_5_7_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_5_7_clkr_en,
      d => yt_rsc_5_7_comp_d,
      q => yt_rsc_5_7_comp_q,
      radr => yt_rsc_5_7_comp_radr,
      wadr => yt_rsc_5_7_comp_wadr,
      we => yt_rsc_5_7_we
    );
  yt_rsc_5_7_comp_d <= yt_rsc_5_7_d;
  yt_rsc_5_7_q <= yt_rsc_5_7_comp_q;
  yt_rsc_5_7_comp_radr <= yt_rsc_5_7_radr;
  yt_rsc_5_7_comp_wadr <= yt_rsc_5_7_wadr;

  yt_rsc_5_8_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_5_8_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_5_8_clkr_en,
      d => yt_rsc_5_8_comp_d,
      q => yt_rsc_5_8_comp_q,
      radr => yt_rsc_5_8_comp_radr,
      wadr => yt_rsc_5_8_comp_wadr,
      we => yt_rsc_5_8_we
    );
  yt_rsc_5_8_comp_d <= yt_rsc_5_8_d;
  yt_rsc_5_8_q <= yt_rsc_5_8_comp_q;
  yt_rsc_5_8_comp_radr <= yt_rsc_5_8_radr;
  yt_rsc_5_8_comp_wadr <= yt_rsc_5_8_wadr;

  yt_rsc_5_9_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_5_9_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_5_9_clkr_en,
      d => yt_rsc_5_9_comp_d,
      q => yt_rsc_5_9_comp_q,
      radr => yt_rsc_5_9_comp_radr,
      wadr => yt_rsc_5_9_comp_wadr,
      we => yt_rsc_5_9_we
    );
  yt_rsc_5_9_comp_d <= yt_rsc_5_9_d;
  yt_rsc_5_9_q <= yt_rsc_5_9_comp_q;
  yt_rsc_5_9_comp_radr <= yt_rsc_5_9_radr;
  yt_rsc_5_9_comp_wadr <= yt_rsc_5_9_wadr;

  yt_rsc_5_10_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_5_10_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_5_10_clkr_en,
      d => yt_rsc_5_10_comp_d,
      q => yt_rsc_5_10_comp_q,
      radr => yt_rsc_5_10_comp_radr,
      wadr => yt_rsc_5_10_comp_wadr,
      we => yt_rsc_5_10_we
    );
  yt_rsc_5_10_comp_d <= yt_rsc_5_10_d;
  yt_rsc_5_10_q <= yt_rsc_5_10_comp_q;
  yt_rsc_5_10_comp_radr <= yt_rsc_5_10_radr;
  yt_rsc_5_10_comp_wadr <= yt_rsc_5_10_wadr;

  yt_rsc_5_11_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_5_11_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_5_11_clkr_en,
      d => yt_rsc_5_11_comp_d,
      q => yt_rsc_5_11_comp_q,
      radr => yt_rsc_5_11_comp_radr,
      wadr => yt_rsc_5_11_comp_wadr,
      we => yt_rsc_5_11_we
    );
  yt_rsc_5_11_comp_d <= yt_rsc_5_11_d;
  yt_rsc_5_11_q <= yt_rsc_5_11_comp_q;
  yt_rsc_5_11_comp_radr <= yt_rsc_5_11_radr;
  yt_rsc_5_11_comp_wadr <= yt_rsc_5_11_wadr;

  yt_rsc_5_12_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_5_12_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_5_12_clkr_en,
      d => yt_rsc_5_12_comp_d,
      q => yt_rsc_5_12_comp_q,
      radr => yt_rsc_5_12_comp_radr,
      wadr => yt_rsc_5_12_comp_wadr,
      we => yt_rsc_5_12_we
    );
  yt_rsc_5_12_comp_d <= yt_rsc_5_12_d;
  yt_rsc_5_12_q <= yt_rsc_5_12_comp_q;
  yt_rsc_5_12_comp_radr <= yt_rsc_5_12_radr;
  yt_rsc_5_12_comp_wadr <= yt_rsc_5_12_wadr;

  yt_rsc_5_13_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_5_13_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_5_13_clkr_en,
      d => yt_rsc_5_13_comp_d,
      q => yt_rsc_5_13_comp_q,
      radr => yt_rsc_5_13_comp_radr,
      wadr => yt_rsc_5_13_comp_wadr,
      we => yt_rsc_5_13_we
    );
  yt_rsc_5_13_comp_d <= yt_rsc_5_13_d;
  yt_rsc_5_13_q <= yt_rsc_5_13_comp_q;
  yt_rsc_5_13_comp_radr <= yt_rsc_5_13_radr;
  yt_rsc_5_13_comp_wadr <= yt_rsc_5_13_wadr;

  yt_rsc_5_14_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_5_14_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_5_14_clkr_en,
      d => yt_rsc_5_14_comp_d,
      q => yt_rsc_5_14_comp_q,
      radr => yt_rsc_5_14_comp_radr,
      wadr => yt_rsc_5_14_comp_wadr,
      we => yt_rsc_5_14_we
    );
  yt_rsc_5_14_comp_d <= yt_rsc_5_14_d;
  yt_rsc_5_14_q <= yt_rsc_5_14_comp_q;
  yt_rsc_5_14_comp_radr <= yt_rsc_5_14_radr;
  yt_rsc_5_14_comp_wadr <= yt_rsc_5_14_wadr;

  yt_rsc_5_15_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_5_15_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_5_15_clkr_en,
      d => yt_rsc_5_15_comp_d,
      q => yt_rsc_5_15_comp_q,
      radr => yt_rsc_5_15_comp_radr,
      wadr => yt_rsc_5_15_comp_wadr,
      we => yt_rsc_5_15_we
    );
  yt_rsc_5_15_comp_d <= yt_rsc_5_15_d;
  yt_rsc_5_15_q <= yt_rsc_5_15_comp_q;
  yt_rsc_5_15_comp_radr <= yt_rsc_5_15_radr;
  yt_rsc_5_15_comp_wadr <= yt_rsc_5_15_wadr;

  yt_rsc_5_16_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_5_16_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_5_16_clkr_en,
      d => yt_rsc_5_16_comp_d,
      q => yt_rsc_5_16_comp_q,
      radr => yt_rsc_5_16_comp_radr,
      wadr => yt_rsc_5_16_comp_wadr,
      we => yt_rsc_5_16_we
    );
  yt_rsc_5_16_comp_d <= yt_rsc_5_16_d;
  yt_rsc_5_16_q <= yt_rsc_5_16_comp_q;
  yt_rsc_5_16_comp_radr <= yt_rsc_5_16_radr;
  yt_rsc_5_16_comp_wadr <= yt_rsc_5_16_wadr;

  yt_rsc_5_17_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_5_17_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_5_17_clkr_en,
      d => yt_rsc_5_17_comp_d,
      q => yt_rsc_5_17_comp_q,
      radr => yt_rsc_5_17_comp_radr,
      wadr => yt_rsc_5_17_comp_wadr,
      we => yt_rsc_5_17_we
    );
  yt_rsc_5_17_comp_d <= yt_rsc_5_17_d;
  yt_rsc_5_17_q <= yt_rsc_5_17_comp_q;
  yt_rsc_5_17_comp_radr <= yt_rsc_5_17_radr;
  yt_rsc_5_17_comp_wadr <= yt_rsc_5_17_wadr;

  yt_rsc_5_18_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_5_18_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_5_18_clkr_en,
      d => yt_rsc_5_18_comp_d,
      q => yt_rsc_5_18_comp_q,
      radr => yt_rsc_5_18_comp_radr,
      wadr => yt_rsc_5_18_comp_wadr,
      we => yt_rsc_5_18_we
    );
  yt_rsc_5_18_comp_d <= yt_rsc_5_18_d;
  yt_rsc_5_18_q <= yt_rsc_5_18_comp_q;
  yt_rsc_5_18_comp_radr <= yt_rsc_5_18_radr;
  yt_rsc_5_18_comp_wadr <= yt_rsc_5_18_wadr;

  yt_rsc_5_19_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_5_19_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_5_19_clkr_en,
      d => yt_rsc_5_19_comp_d,
      q => yt_rsc_5_19_comp_q,
      radr => yt_rsc_5_19_comp_radr,
      wadr => yt_rsc_5_19_comp_wadr,
      we => yt_rsc_5_19_we
    );
  yt_rsc_5_19_comp_d <= yt_rsc_5_19_d;
  yt_rsc_5_19_q <= yt_rsc_5_19_comp_q;
  yt_rsc_5_19_comp_radr <= yt_rsc_5_19_radr;
  yt_rsc_5_19_comp_wadr <= yt_rsc_5_19_wadr;

  yt_rsc_5_20_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_5_20_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_5_20_clkr_en,
      d => yt_rsc_5_20_comp_d,
      q => yt_rsc_5_20_comp_q,
      radr => yt_rsc_5_20_comp_radr,
      wadr => yt_rsc_5_20_comp_wadr,
      we => yt_rsc_5_20_we
    );
  yt_rsc_5_20_comp_d <= yt_rsc_5_20_d;
  yt_rsc_5_20_q <= yt_rsc_5_20_comp_q;
  yt_rsc_5_20_comp_radr <= yt_rsc_5_20_radr;
  yt_rsc_5_20_comp_wadr <= yt_rsc_5_20_wadr;

  yt_rsc_5_21_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_5_21_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_5_21_clkr_en,
      d => yt_rsc_5_21_comp_d,
      q => yt_rsc_5_21_comp_q,
      radr => yt_rsc_5_21_comp_radr,
      wadr => yt_rsc_5_21_comp_wadr,
      we => yt_rsc_5_21_we
    );
  yt_rsc_5_21_comp_d <= yt_rsc_5_21_d;
  yt_rsc_5_21_q <= yt_rsc_5_21_comp_q;
  yt_rsc_5_21_comp_radr <= yt_rsc_5_21_radr;
  yt_rsc_5_21_comp_wadr <= yt_rsc_5_21_wadr;

  yt_rsc_5_22_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_5_22_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_5_22_clkr_en,
      d => yt_rsc_5_22_comp_d,
      q => yt_rsc_5_22_comp_q,
      radr => yt_rsc_5_22_comp_radr,
      wadr => yt_rsc_5_22_comp_wadr,
      we => yt_rsc_5_22_we
    );
  yt_rsc_5_22_comp_d <= yt_rsc_5_22_d;
  yt_rsc_5_22_q <= yt_rsc_5_22_comp_q;
  yt_rsc_5_22_comp_radr <= yt_rsc_5_22_radr;
  yt_rsc_5_22_comp_wadr <= yt_rsc_5_22_wadr;

  yt_rsc_5_23_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_5_23_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_5_23_clkr_en,
      d => yt_rsc_5_23_comp_d,
      q => yt_rsc_5_23_comp_q,
      radr => yt_rsc_5_23_comp_radr,
      wadr => yt_rsc_5_23_comp_wadr,
      we => yt_rsc_5_23_we
    );
  yt_rsc_5_23_comp_d <= yt_rsc_5_23_d;
  yt_rsc_5_23_q <= yt_rsc_5_23_comp_q;
  yt_rsc_5_23_comp_radr <= yt_rsc_5_23_radr;
  yt_rsc_5_23_comp_wadr <= yt_rsc_5_23_wadr;

  yt_rsc_5_24_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_5_24_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_5_24_clkr_en,
      d => yt_rsc_5_24_comp_d,
      q => yt_rsc_5_24_comp_q,
      radr => yt_rsc_5_24_comp_radr,
      wadr => yt_rsc_5_24_comp_wadr,
      we => yt_rsc_5_24_we
    );
  yt_rsc_5_24_comp_d <= yt_rsc_5_24_d;
  yt_rsc_5_24_q <= yt_rsc_5_24_comp_q;
  yt_rsc_5_24_comp_radr <= yt_rsc_5_24_radr;
  yt_rsc_5_24_comp_wadr <= yt_rsc_5_24_wadr;

  yt_rsc_5_25_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_5_25_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_5_25_clkr_en,
      d => yt_rsc_5_25_comp_d,
      q => yt_rsc_5_25_comp_q,
      radr => yt_rsc_5_25_comp_radr,
      wadr => yt_rsc_5_25_comp_wadr,
      we => yt_rsc_5_25_we
    );
  yt_rsc_5_25_comp_d <= yt_rsc_5_25_d;
  yt_rsc_5_25_q <= yt_rsc_5_25_comp_q;
  yt_rsc_5_25_comp_radr <= yt_rsc_5_25_radr;
  yt_rsc_5_25_comp_wadr <= yt_rsc_5_25_wadr;

  yt_rsc_5_26_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_5_26_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_5_26_clkr_en,
      d => yt_rsc_5_26_comp_d,
      q => yt_rsc_5_26_comp_q,
      radr => yt_rsc_5_26_comp_radr,
      wadr => yt_rsc_5_26_comp_wadr,
      we => yt_rsc_5_26_we
    );
  yt_rsc_5_26_comp_d <= yt_rsc_5_26_d;
  yt_rsc_5_26_q <= yt_rsc_5_26_comp_q;
  yt_rsc_5_26_comp_radr <= yt_rsc_5_26_radr;
  yt_rsc_5_26_comp_wadr <= yt_rsc_5_26_wadr;

  yt_rsc_5_27_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_5_27_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_5_27_clkr_en,
      d => yt_rsc_5_27_comp_d,
      q => yt_rsc_5_27_comp_q,
      radr => yt_rsc_5_27_comp_radr,
      wadr => yt_rsc_5_27_comp_wadr,
      we => yt_rsc_5_27_we
    );
  yt_rsc_5_27_comp_d <= yt_rsc_5_27_d;
  yt_rsc_5_27_q <= yt_rsc_5_27_comp_q;
  yt_rsc_5_27_comp_radr <= yt_rsc_5_27_radr;
  yt_rsc_5_27_comp_wadr <= yt_rsc_5_27_wadr;

  yt_rsc_5_28_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_5_28_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_5_28_clkr_en,
      d => yt_rsc_5_28_comp_d,
      q => yt_rsc_5_28_comp_q,
      radr => yt_rsc_5_28_comp_radr,
      wadr => yt_rsc_5_28_comp_wadr,
      we => yt_rsc_5_28_we
    );
  yt_rsc_5_28_comp_d <= yt_rsc_5_28_d;
  yt_rsc_5_28_q <= yt_rsc_5_28_comp_q;
  yt_rsc_5_28_comp_radr <= yt_rsc_5_28_radr;
  yt_rsc_5_28_comp_wadr <= yt_rsc_5_28_wadr;

  yt_rsc_5_29_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_5_29_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_5_29_clkr_en,
      d => yt_rsc_5_29_comp_d,
      q => yt_rsc_5_29_comp_q,
      radr => yt_rsc_5_29_comp_radr,
      wadr => yt_rsc_5_29_comp_wadr,
      we => yt_rsc_5_29_we
    );
  yt_rsc_5_29_comp_d <= yt_rsc_5_29_d;
  yt_rsc_5_29_q <= yt_rsc_5_29_comp_q;
  yt_rsc_5_29_comp_radr <= yt_rsc_5_29_radr;
  yt_rsc_5_29_comp_wadr <= yt_rsc_5_29_wadr;

  yt_rsc_5_30_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_5_30_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_5_30_clkr_en,
      d => yt_rsc_5_30_comp_d,
      q => yt_rsc_5_30_comp_q,
      radr => yt_rsc_5_30_comp_radr,
      wadr => yt_rsc_5_30_comp_wadr,
      we => yt_rsc_5_30_we
    );
  yt_rsc_5_30_comp_d <= yt_rsc_5_30_d;
  yt_rsc_5_30_q <= yt_rsc_5_30_comp_q;
  yt_rsc_5_30_comp_radr <= yt_rsc_5_30_radr;
  yt_rsc_5_30_comp_wadr <= yt_rsc_5_30_wadr;

  yt_rsc_5_31_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_5_31_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_5_31_clkr_en,
      d => yt_rsc_5_31_comp_d,
      q => yt_rsc_5_31_comp_q,
      radr => yt_rsc_5_31_comp_radr,
      wadr => yt_rsc_5_31_comp_wadr,
      we => yt_rsc_5_31_we
    );
  yt_rsc_5_31_comp_d <= yt_rsc_5_31_d;
  yt_rsc_5_31_q <= yt_rsc_5_31_comp_q;
  yt_rsc_5_31_comp_radr <= yt_rsc_5_31_radr;
  yt_rsc_5_31_comp_wadr <= yt_rsc_5_31_wadr;

  yt_rsc_6_0_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_6_0_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_6_0_clkr_en,
      d => yt_rsc_6_0_comp_d,
      q => yt_rsc_6_0_comp_q,
      radr => yt_rsc_6_0_comp_radr,
      wadr => yt_rsc_6_0_comp_wadr,
      we => yt_rsc_6_0_we
    );
  yt_rsc_6_0_comp_d <= yt_rsc_6_0_d;
  yt_rsc_6_0_q <= yt_rsc_6_0_comp_q;
  yt_rsc_6_0_comp_radr <= yt_rsc_6_0_radr;
  yt_rsc_6_0_comp_wadr <= yt_rsc_6_0_wadr;

  yt_rsc_6_1_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_6_1_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_6_1_clkr_en,
      d => yt_rsc_6_1_comp_d,
      q => yt_rsc_6_1_comp_q,
      radr => yt_rsc_6_1_comp_radr,
      wadr => yt_rsc_6_1_comp_wadr,
      we => yt_rsc_6_1_we
    );
  yt_rsc_6_1_comp_d <= yt_rsc_6_1_d;
  yt_rsc_6_1_q <= yt_rsc_6_1_comp_q;
  yt_rsc_6_1_comp_radr <= yt_rsc_6_1_radr;
  yt_rsc_6_1_comp_wadr <= yt_rsc_6_1_wadr;

  yt_rsc_6_2_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_6_2_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_6_2_clkr_en,
      d => yt_rsc_6_2_comp_d,
      q => yt_rsc_6_2_comp_q,
      radr => yt_rsc_6_2_comp_radr,
      wadr => yt_rsc_6_2_comp_wadr,
      we => yt_rsc_6_2_we
    );
  yt_rsc_6_2_comp_d <= yt_rsc_6_2_d;
  yt_rsc_6_2_q <= yt_rsc_6_2_comp_q;
  yt_rsc_6_2_comp_radr <= yt_rsc_6_2_radr;
  yt_rsc_6_2_comp_wadr <= yt_rsc_6_2_wadr;

  yt_rsc_6_3_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_6_3_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_6_3_clkr_en,
      d => yt_rsc_6_3_comp_d,
      q => yt_rsc_6_3_comp_q,
      radr => yt_rsc_6_3_comp_radr,
      wadr => yt_rsc_6_3_comp_wadr,
      we => yt_rsc_6_3_we
    );
  yt_rsc_6_3_comp_d <= yt_rsc_6_3_d;
  yt_rsc_6_3_q <= yt_rsc_6_3_comp_q;
  yt_rsc_6_3_comp_radr <= yt_rsc_6_3_radr;
  yt_rsc_6_3_comp_wadr <= yt_rsc_6_3_wadr;

  yt_rsc_6_4_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_6_4_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_6_4_clkr_en,
      d => yt_rsc_6_4_comp_d,
      q => yt_rsc_6_4_comp_q,
      radr => yt_rsc_6_4_comp_radr,
      wadr => yt_rsc_6_4_comp_wadr,
      we => yt_rsc_6_4_we
    );
  yt_rsc_6_4_comp_d <= yt_rsc_6_4_d;
  yt_rsc_6_4_q <= yt_rsc_6_4_comp_q;
  yt_rsc_6_4_comp_radr <= yt_rsc_6_4_radr;
  yt_rsc_6_4_comp_wadr <= yt_rsc_6_4_wadr;

  yt_rsc_6_5_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_6_5_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_6_5_clkr_en,
      d => yt_rsc_6_5_comp_d,
      q => yt_rsc_6_5_comp_q,
      radr => yt_rsc_6_5_comp_radr,
      wadr => yt_rsc_6_5_comp_wadr,
      we => yt_rsc_6_5_we
    );
  yt_rsc_6_5_comp_d <= yt_rsc_6_5_d;
  yt_rsc_6_5_q <= yt_rsc_6_5_comp_q;
  yt_rsc_6_5_comp_radr <= yt_rsc_6_5_radr;
  yt_rsc_6_5_comp_wadr <= yt_rsc_6_5_wadr;

  yt_rsc_6_6_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_6_6_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_6_6_clkr_en,
      d => yt_rsc_6_6_comp_d,
      q => yt_rsc_6_6_comp_q,
      radr => yt_rsc_6_6_comp_radr,
      wadr => yt_rsc_6_6_comp_wadr,
      we => yt_rsc_6_6_we
    );
  yt_rsc_6_6_comp_d <= yt_rsc_6_6_d;
  yt_rsc_6_6_q <= yt_rsc_6_6_comp_q;
  yt_rsc_6_6_comp_radr <= yt_rsc_6_6_radr;
  yt_rsc_6_6_comp_wadr <= yt_rsc_6_6_wadr;

  yt_rsc_6_7_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_6_7_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_6_7_clkr_en,
      d => yt_rsc_6_7_comp_d,
      q => yt_rsc_6_7_comp_q,
      radr => yt_rsc_6_7_comp_radr,
      wadr => yt_rsc_6_7_comp_wadr,
      we => yt_rsc_6_7_we
    );
  yt_rsc_6_7_comp_d <= yt_rsc_6_7_d;
  yt_rsc_6_7_q <= yt_rsc_6_7_comp_q;
  yt_rsc_6_7_comp_radr <= yt_rsc_6_7_radr;
  yt_rsc_6_7_comp_wadr <= yt_rsc_6_7_wadr;

  yt_rsc_6_8_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_6_8_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_6_8_clkr_en,
      d => yt_rsc_6_8_comp_d,
      q => yt_rsc_6_8_comp_q,
      radr => yt_rsc_6_8_comp_radr,
      wadr => yt_rsc_6_8_comp_wadr,
      we => yt_rsc_6_8_we
    );
  yt_rsc_6_8_comp_d <= yt_rsc_6_8_d;
  yt_rsc_6_8_q <= yt_rsc_6_8_comp_q;
  yt_rsc_6_8_comp_radr <= yt_rsc_6_8_radr;
  yt_rsc_6_8_comp_wadr <= yt_rsc_6_8_wadr;

  yt_rsc_6_9_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_6_9_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_6_9_clkr_en,
      d => yt_rsc_6_9_comp_d,
      q => yt_rsc_6_9_comp_q,
      radr => yt_rsc_6_9_comp_radr,
      wadr => yt_rsc_6_9_comp_wadr,
      we => yt_rsc_6_9_we
    );
  yt_rsc_6_9_comp_d <= yt_rsc_6_9_d;
  yt_rsc_6_9_q <= yt_rsc_6_9_comp_q;
  yt_rsc_6_9_comp_radr <= yt_rsc_6_9_radr;
  yt_rsc_6_9_comp_wadr <= yt_rsc_6_9_wadr;

  yt_rsc_6_10_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_6_10_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_6_10_clkr_en,
      d => yt_rsc_6_10_comp_d,
      q => yt_rsc_6_10_comp_q,
      radr => yt_rsc_6_10_comp_radr,
      wadr => yt_rsc_6_10_comp_wadr,
      we => yt_rsc_6_10_we
    );
  yt_rsc_6_10_comp_d <= yt_rsc_6_10_d;
  yt_rsc_6_10_q <= yt_rsc_6_10_comp_q;
  yt_rsc_6_10_comp_radr <= yt_rsc_6_10_radr;
  yt_rsc_6_10_comp_wadr <= yt_rsc_6_10_wadr;

  yt_rsc_6_11_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_6_11_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_6_11_clkr_en,
      d => yt_rsc_6_11_comp_d,
      q => yt_rsc_6_11_comp_q,
      radr => yt_rsc_6_11_comp_radr,
      wadr => yt_rsc_6_11_comp_wadr,
      we => yt_rsc_6_11_we
    );
  yt_rsc_6_11_comp_d <= yt_rsc_6_11_d;
  yt_rsc_6_11_q <= yt_rsc_6_11_comp_q;
  yt_rsc_6_11_comp_radr <= yt_rsc_6_11_radr;
  yt_rsc_6_11_comp_wadr <= yt_rsc_6_11_wadr;

  yt_rsc_6_12_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_6_12_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_6_12_clkr_en,
      d => yt_rsc_6_12_comp_d,
      q => yt_rsc_6_12_comp_q,
      radr => yt_rsc_6_12_comp_radr,
      wadr => yt_rsc_6_12_comp_wadr,
      we => yt_rsc_6_12_we
    );
  yt_rsc_6_12_comp_d <= yt_rsc_6_12_d;
  yt_rsc_6_12_q <= yt_rsc_6_12_comp_q;
  yt_rsc_6_12_comp_radr <= yt_rsc_6_12_radr;
  yt_rsc_6_12_comp_wadr <= yt_rsc_6_12_wadr;

  yt_rsc_6_13_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_6_13_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_6_13_clkr_en,
      d => yt_rsc_6_13_comp_d,
      q => yt_rsc_6_13_comp_q,
      radr => yt_rsc_6_13_comp_radr,
      wadr => yt_rsc_6_13_comp_wadr,
      we => yt_rsc_6_13_we
    );
  yt_rsc_6_13_comp_d <= yt_rsc_6_13_d;
  yt_rsc_6_13_q <= yt_rsc_6_13_comp_q;
  yt_rsc_6_13_comp_radr <= yt_rsc_6_13_radr;
  yt_rsc_6_13_comp_wadr <= yt_rsc_6_13_wadr;

  yt_rsc_6_14_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_6_14_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_6_14_clkr_en,
      d => yt_rsc_6_14_comp_d,
      q => yt_rsc_6_14_comp_q,
      radr => yt_rsc_6_14_comp_radr,
      wadr => yt_rsc_6_14_comp_wadr,
      we => yt_rsc_6_14_we
    );
  yt_rsc_6_14_comp_d <= yt_rsc_6_14_d;
  yt_rsc_6_14_q <= yt_rsc_6_14_comp_q;
  yt_rsc_6_14_comp_radr <= yt_rsc_6_14_radr;
  yt_rsc_6_14_comp_wadr <= yt_rsc_6_14_wadr;

  yt_rsc_6_15_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_6_15_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_6_15_clkr_en,
      d => yt_rsc_6_15_comp_d,
      q => yt_rsc_6_15_comp_q,
      radr => yt_rsc_6_15_comp_radr,
      wadr => yt_rsc_6_15_comp_wadr,
      we => yt_rsc_6_15_we
    );
  yt_rsc_6_15_comp_d <= yt_rsc_6_15_d;
  yt_rsc_6_15_q <= yt_rsc_6_15_comp_q;
  yt_rsc_6_15_comp_radr <= yt_rsc_6_15_radr;
  yt_rsc_6_15_comp_wadr <= yt_rsc_6_15_wadr;

  yt_rsc_6_16_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_6_16_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_6_16_clkr_en,
      d => yt_rsc_6_16_comp_d,
      q => yt_rsc_6_16_comp_q,
      radr => yt_rsc_6_16_comp_radr,
      wadr => yt_rsc_6_16_comp_wadr,
      we => yt_rsc_6_16_we
    );
  yt_rsc_6_16_comp_d <= yt_rsc_6_16_d;
  yt_rsc_6_16_q <= yt_rsc_6_16_comp_q;
  yt_rsc_6_16_comp_radr <= yt_rsc_6_16_radr;
  yt_rsc_6_16_comp_wadr <= yt_rsc_6_16_wadr;

  yt_rsc_6_17_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_6_17_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_6_17_clkr_en,
      d => yt_rsc_6_17_comp_d,
      q => yt_rsc_6_17_comp_q,
      radr => yt_rsc_6_17_comp_radr,
      wadr => yt_rsc_6_17_comp_wadr,
      we => yt_rsc_6_17_we
    );
  yt_rsc_6_17_comp_d <= yt_rsc_6_17_d;
  yt_rsc_6_17_q <= yt_rsc_6_17_comp_q;
  yt_rsc_6_17_comp_radr <= yt_rsc_6_17_radr;
  yt_rsc_6_17_comp_wadr <= yt_rsc_6_17_wadr;

  yt_rsc_6_18_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_6_18_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_6_18_clkr_en,
      d => yt_rsc_6_18_comp_d,
      q => yt_rsc_6_18_comp_q,
      radr => yt_rsc_6_18_comp_radr,
      wadr => yt_rsc_6_18_comp_wadr,
      we => yt_rsc_6_18_we
    );
  yt_rsc_6_18_comp_d <= yt_rsc_6_18_d;
  yt_rsc_6_18_q <= yt_rsc_6_18_comp_q;
  yt_rsc_6_18_comp_radr <= yt_rsc_6_18_radr;
  yt_rsc_6_18_comp_wadr <= yt_rsc_6_18_wadr;

  yt_rsc_6_19_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_6_19_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_6_19_clkr_en,
      d => yt_rsc_6_19_comp_d,
      q => yt_rsc_6_19_comp_q,
      radr => yt_rsc_6_19_comp_radr,
      wadr => yt_rsc_6_19_comp_wadr,
      we => yt_rsc_6_19_we
    );
  yt_rsc_6_19_comp_d <= yt_rsc_6_19_d;
  yt_rsc_6_19_q <= yt_rsc_6_19_comp_q;
  yt_rsc_6_19_comp_radr <= yt_rsc_6_19_radr;
  yt_rsc_6_19_comp_wadr <= yt_rsc_6_19_wadr;

  yt_rsc_6_20_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_6_20_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_6_20_clkr_en,
      d => yt_rsc_6_20_comp_d,
      q => yt_rsc_6_20_comp_q,
      radr => yt_rsc_6_20_comp_radr,
      wadr => yt_rsc_6_20_comp_wadr,
      we => yt_rsc_6_20_we
    );
  yt_rsc_6_20_comp_d <= yt_rsc_6_20_d;
  yt_rsc_6_20_q <= yt_rsc_6_20_comp_q;
  yt_rsc_6_20_comp_radr <= yt_rsc_6_20_radr;
  yt_rsc_6_20_comp_wadr <= yt_rsc_6_20_wadr;

  yt_rsc_6_21_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_6_21_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_6_21_clkr_en,
      d => yt_rsc_6_21_comp_d,
      q => yt_rsc_6_21_comp_q,
      radr => yt_rsc_6_21_comp_radr,
      wadr => yt_rsc_6_21_comp_wadr,
      we => yt_rsc_6_21_we
    );
  yt_rsc_6_21_comp_d <= yt_rsc_6_21_d;
  yt_rsc_6_21_q <= yt_rsc_6_21_comp_q;
  yt_rsc_6_21_comp_radr <= yt_rsc_6_21_radr;
  yt_rsc_6_21_comp_wadr <= yt_rsc_6_21_wadr;

  yt_rsc_6_22_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_6_22_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_6_22_clkr_en,
      d => yt_rsc_6_22_comp_d,
      q => yt_rsc_6_22_comp_q,
      radr => yt_rsc_6_22_comp_radr,
      wadr => yt_rsc_6_22_comp_wadr,
      we => yt_rsc_6_22_we
    );
  yt_rsc_6_22_comp_d <= yt_rsc_6_22_d;
  yt_rsc_6_22_q <= yt_rsc_6_22_comp_q;
  yt_rsc_6_22_comp_radr <= yt_rsc_6_22_radr;
  yt_rsc_6_22_comp_wadr <= yt_rsc_6_22_wadr;

  yt_rsc_6_23_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_6_23_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_6_23_clkr_en,
      d => yt_rsc_6_23_comp_d,
      q => yt_rsc_6_23_comp_q,
      radr => yt_rsc_6_23_comp_radr,
      wadr => yt_rsc_6_23_comp_wadr,
      we => yt_rsc_6_23_we
    );
  yt_rsc_6_23_comp_d <= yt_rsc_6_23_d;
  yt_rsc_6_23_q <= yt_rsc_6_23_comp_q;
  yt_rsc_6_23_comp_radr <= yt_rsc_6_23_radr;
  yt_rsc_6_23_comp_wadr <= yt_rsc_6_23_wadr;

  yt_rsc_6_24_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_6_24_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_6_24_clkr_en,
      d => yt_rsc_6_24_comp_d,
      q => yt_rsc_6_24_comp_q,
      radr => yt_rsc_6_24_comp_radr,
      wadr => yt_rsc_6_24_comp_wadr,
      we => yt_rsc_6_24_we
    );
  yt_rsc_6_24_comp_d <= yt_rsc_6_24_d;
  yt_rsc_6_24_q <= yt_rsc_6_24_comp_q;
  yt_rsc_6_24_comp_radr <= yt_rsc_6_24_radr;
  yt_rsc_6_24_comp_wadr <= yt_rsc_6_24_wadr;

  yt_rsc_6_25_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_6_25_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_6_25_clkr_en,
      d => yt_rsc_6_25_comp_d,
      q => yt_rsc_6_25_comp_q,
      radr => yt_rsc_6_25_comp_radr,
      wadr => yt_rsc_6_25_comp_wadr,
      we => yt_rsc_6_25_we
    );
  yt_rsc_6_25_comp_d <= yt_rsc_6_25_d;
  yt_rsc_6_25_q <= yt_rsc_6_25_comp_q;
  yt_rsc_6_25_comp_radr <= yt_rsc_6_25_radr;
  yt_rsc_6_25_comp_wadr <= yt_rsc_6_25_wadr;

  yt_rsc_6_26_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_6_26_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_6_26_clkr_en,
      d => yt_rsc_6_26_comp_d,
      q => yt_rsc_6_26_comp_q,
      radr => yt_rsc_6_26_comp_radr,
      wadr => yt_rsc_6_26_comp_wadr,
      we => yt_rsc_6_26_we
    );
  yt_rsc_6_26_comp_d <= yt_rsc_6_26_d;
  yt_rsc_6_26_q <= yt_rsc_6_26_comp_q;
  yt_rsc_6_26_comp_radr <= yt_rsc_6_26_radr;
  yt_rsc_6_26_comp_wadr <= yt_rsc_6_26_wadr;

  yt_rsc_6_27_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_6_27_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_6_27_clkr_en,
      d => yt_rsc_6_27_comp_d,
      q => yt_rsc_6_27_comp_q,
      radr => yt_rsc_6_27_comp_radr,
      wadr => yt_rsc_6_27_comp_wadr,
      we => yt_rsc_6_27_we
    );
  yt_rsc_6_27_comp_d <= yt_rsc_6_27_d;
  yt_rsc_6_27_q <= yt_rsc_6_27_comp_q;
  yt_rsc_6_27_comp_radr <= yt_rsc_6_27_radr;
  yt_rsc_6_27_comp_wadr <= yt_rsc_6_27_wadr;

  yt_rsc_6_28_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_6_28_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_6_28_clkr_en,
      d => yt_rsc_6_28_comp_d,
      q => yt_rsc_6_28_comp_q,
      radr => yt_rsc_6_28_comp_radr,
      wadr => yt_rsc_6_28_comp_wadr,
      we => yt_rsc_6_28_we
    );
  yt_rsc_6_28_comp_d <= yt_rsc_6_28_d;
  yt_rsc_6_28_q <= yt_rsc_6_28_comp_q;
  yt_rsc_6_28_comp_radr <= yt_rsc_6_28_radr;
  yt_rsc_6_28_comp_wadr <= yt_rsc_6_28_wadr;

  yt_rsc_6_29_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_6_29_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_6_29_clkr_en,
      d => yt_rsc_6_29_comp_d,
      q => yt_rsc_6_29_comp_q,
      radr => yt_rsc_6_29_comp_radr,
      wadr => yt_rsc_6_29_comp_wadr,
      we => yt_rsc_6_29_we
    );
  yt_rsc_6_29_comp_d <= yt_rsc_6_29_d;
  yt_rsc_6_29_q <= yt_rsc_6_29_comp_q;
  yt_rsc_6_29_comp_radr <= yt_rsc_6_29_radr;
  yt_rsc_6_29_comp_wadr <= yt_rsc_6_29_wadr;

  yt_rsc_6_30_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_6_30_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_6_30_clkr_en,
      d => yt_rsc_6_30_comp_d,
      q => yt_rsc_6_30_comp_q,
      radr => yt_rsc_6_30_comp_radr,
      wadr => yt_rsc_6_30_comp_wadr,
      we => yt_rsc_6_30_we
    );
  yt_rsc_6_30_comp_d <= yt_rsc_6_30_d;
  yt_rsc_6_30_q <= yt_rsc_6_30_comp_q;
  yt_rsc_6_30_comp_radr <= yt_rsc_6_30_radr;
  yt_rsc_6_30_comp_wadr <= yt_rsc_6_30_wadr;

  yt_rsc_6_31_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_6_31_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_6_31_clkr_en,
      d => yt_rsc_6_31_comp_d,
      q => yt_rsc_6_31_comp_q,
      radr => yt_rsc_6_31_comp_radr,
      wadr => yt_rsc_6_31_comp_wadr,
      we => yt_rsc_6_31_we
    );
  yt_rsc_6_31_comp_d <= yt_rsc_6_31_d;
  yt_rsc_6_31_q <= yt_rsc_6_31_comp_q;
  yt_rsc_6_31_comp_radr <= yt_rsc_6_31_radr;
  yt_rsc_6_31_comp_wadr <= yt_rsc_6_31_wadr;

  yt_rsc_7_0_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_7_0_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_7_0_clkr_en,
      d => yt_rsc_7_0_comp_d,
      q => yt_rsc_7_0_comp_q,
      radr => yt_rsc_7_0_comp_radr,
      wadr => yt_rsc_7_0_comp_wadr,
      we => yt_rsc_7_0_we
    );
  yt_rsc_7_0_comp_d <= yt_rsc_7_0_d;
  yt_rsc_7_0_q <= yt_rsc_7_0_comp_q;
  yt_rsc_7_0_comp_radr <= yt_rsc_7_0_radr;
  yt_rsc_7_0_comp_wadr <= yt_rsc_7_0_wadr;

  yt_rsc_7_1_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_7_1_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_7_1_clkr_en,
      d => yt_rsc_7_1_comp_d,
      q => yt_rsc_7_1_comp_q,
      radr => yt_rsc_7_1_comp_radr,
      wadr => yt_rsc_7_1_comp_wadr,
      we => yt_rsc_7_1_we
    );
  yt_rsc_7_1_comp_d <= yt_rsc_7_1_d;
  yt_rsc_7_1_q <= yt_rsc_7_1_comp_q;
  yt_rsc_7_1_comp_radr <= yt_rsc_7_1_radr;
  yt_rsc_7_1_comp_wadr <= yt_rsc_7_1_wadr;

  yt_rsc_7_2_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_7_2_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_7_2_clkr_en,
      d => yt_rsc_7_2_comp_d,
      q => yt_rsc_7_2_comp_q,
      radr => yt_rsc_7_2_comp_radr,
      wadr => yt_rsc_7_2_comp_wadr,
      we => yt_rsc_7_2_we
    );
  yt_rsc_7_2_comp_d <= yt_rsc_7_2_d;
  yt_rsc_7_2_q <= yt_rsc_7_2_comp_q;
  yt_rsc_7_2_comp_radr <= yt_rsc_7_2_radr;
  yt_rsc_7_2_comp_wadr <= yt_rsc_7_2_wadr;

  yt_rsc_7_3_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_7_3_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_7_3_clkr_en,
      d => yt_rsc_7_3_comp_d,
      q => yt_rsc_7_3_comp_q,
      radr => yt_rsc_7_3_comp_radr,
      wadr => yt_rsc_7_3_comp_wadr,
      we => yt_rsc_7_3_we
    );
  yt_rsc_7_3_comp_d <= yt_rsc_7_3_d;
  yt_rsc_7_3_q <= yt_rsc_7_3_comp_q;
  yt_rsc_7_3_comp_radr <= yt_rsc_7_3_radr;
  yt_rsc_7_3_comp_wadr <= yt_rsc_7_3_wadr;

  yt_rsc_7_4_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_7_4_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_7_4_clkr_en,
      d => yt_rsc_7_4_comp_d,
      q => yt_rsc_7_4_comp_q,
      radr => yt_rsc_7_4_comp_radr,
      wadr => yt_rsc_7_4_comp_wadr,
      we => yt_rsc_7_4_we
    );
  yt_rsc_7_4_comp_d <= yt_rsc_7_4_d;
  yt_rsc_7_4_q <= yt_rsc_7_4_comp_q;
  yt_rsc_7_4_comp_radr <= yt_rsc_7_4_radr;
  yt_rsc_7_4_comp_wadr <= yt_rsc_7_4_wadr;

  yt_rsc_7_5_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_7_5_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_7_5_clkr_en,
      d => yt_rsc_7_5_comp_d,
      q => yt_rsc_7_5_comp_q,
      radr => yt_rsc_7_5_comp_radr,
      wadr => yt_rsc_7_5_comp_wadr,
      we => yt_rsc_7_5_we
    );
  yt_rsc_7_5_comp_d <= yt_rsc_7_5_d;
  yt_rsc_7_5_q <= yt_rsc_7_5_comp_q;
  yt_rsc_7_5_comp_radr <= yt_rsc_7_5_radr;
  yt_rsc_7_5_comp_wadr <= yt_rsc_7_5_wadr;

  yt_rsc_7_6_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_7_6_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_7_6_clkr_en,
      d => yt_rsc_7_6_comp_d,
      q => yt_rsc_7_6_comp_q,
      radr => yt_rsc_7_6_comp_radr,
      wadr => yt_rsc_7_6_comp_wadr,
      we => yt_rsc_7_6_we
    );
  yt_rsc_7_6_comp_d <= yt_rsc_7_6_d;
  yt_rsc_7_6_q <= yt_rsc_7_6_comp_q;
  yt_rsc_7_6_comp_radr <= yt_rsc_7_6_radr;
  yt_rsc_7_6_comp_wadr <= yt_rsc_7_6_wadr;

  yt_rsc_7_7_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_7_7_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_7_7_clkr_en,
      d => yt_rsc_7_7_comp_d,
      q => yt_rsc_7_7_comp_q,
      radr => yt_rsc_7_7_comp_radr,
      wadr => yt_rsc_7_7_comp_wadr,
      we => yt_rsc_7_7_we
    );
  yt_rsc_7_7_comp_d <= yt_rsc_7_7_d;
  yt_rsc_7_7_q <= yt_rsc_7_7_comp_q;
  yt_rsc_7_7_comp_radr <= yt_rsc_7_7_radr;
  yt_rsc_7_7_comp_wadr <= yt_rsc_7_7_wadr;

  yt_rsc_7_8_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_7_8_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_7_8_clkr_en,
      d => yt_rsc_7_8_comp_d,
      q => yt_rsc_7_8_comp_q,
      radr => yt_rsc_7_8_comp_radr,
      wadr => yt_rsc_7_8_comp_wadr,
      we => yt_rsc_7_8_we
    );
  yt_rsc_7_8_comp_d <= yt_rsc_7_8_d;
  yt_rsc_7_8_q <= yt_rsc_7_8_comp_q;
  yt_rsc_7_8_comp_radr <= yt_rsc_7_8_radr;
  yt_rsc_7_8_comp_wadr <= yt_rsc_7_8_wadr;

  yt_rsc_7_9_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_7_9_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_7_9_clkr_en,
      d => yt_rsc_7_9_comp_d,
      q => yt_rsc_7_9_comp_q,
      radr => yt_rsc_7_9_comp_radr,
      wadr => yt_rsc_7_9_comp_wadr,
      we => yt_rsc_7_9_we
    );
  yt_rsc_7_9_comp_d <= yt_rsc_7_9_d;
  yt_rsc_7_9_q <= yt_rsc_7_9_comp_q;
  yt_rsc_7_9_comp_radr <= yt_rsc_7_9_radr;
  yt_rsc_7_9_comp_wadr <= yt_rsc_7_9_wadr;

  yt_rsc_7_10_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_7_10_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_7_10_clkr_en,
      d => yt_rsc_7_10_comp_d,
      q => yt_rsc_7_10_comp_q,
      radr => yt_rsc_7_10_comp_radr,
      wadr => yt_rsc_7_10_comp_wadr,
      we => yt_rsc_7_10_we
    );
  yt_rsc_7_10_comp_d <= yt_rsc_7_10_d;
  yt_rsc_7_10_q <= yt_rsc_7_10_comp_q;
  yt_rsc_7_10_comp_radr <= yt_rsc_7_10_radr;
  yt_rsc_7_10_comp_wadr <= yt_rsc_7_10_wadr;

  yt_rsc_7_11_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_7_11_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_7_11_clkr_en,
      d => yt_rsc_7_11_comp_d,
      q => yt_rsc_7_11_comp_q,
      radr => yt_rsc_7_11_comp_radr,
      wadr => yt_rsc_7_11_comp_wadr,
      we => yt_rsc_7_11_we
    );
  yt_rsc_7_11_comp_d <= yt_rsc_7_11_d;
  yt_rsc_7_11_q <= yt_rsc_7_11_comp_q;
  yt_rsc_7_11_comp_radr <= yt_rsc_7_11_radr;
  yt_rsc_7_11_comp_wadr <= yt_rsc_7_11_wadr;

  yt_rsc_7_12_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_7_12_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_7_12_clkr_en,
      d => yt_rsc_7_12_comp_d,
      q => yt_rsc_7_12_comp_q,
      radr => yt_rsc_7_12_comp_radr,
      wadr => yt_rsc_7_12_comp_wadr,
      we => yt_rsc_7_12_we
    );
  yt_rsc_7_12_comp_d <= yt_rsc_7_12_d;
  yt_rsc_7_12_q <= yt_rsc_7_12_comp_q;
  yt_rsc_7_12_comp_radr <= yt_rsc_7_12_radr;
  yt_rsc_7_12_comp_wadr <= yt_rsc_7_12_wadr;

  yt_rsc_7_13_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_7_13_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_7_13_clkr_en,
      d => yt_rsc_7_13_comp_d,
      q => yt_rsc_7_13_comp_q,
      radr => yt_rsc_7_13_comp_radr,
      wadr => yt_rsc_7_13_comp_wadr,
      we => yt_rsc_7_13_we
    );
  yt_rsc_7_13_comp_d <= yt_rsc_7_13_d;
  yt_rsc_7_13_q <= yt_rsc_7_13_comp_q;
  yt_rsc_7_13_comp_radr <= yt_rsc_7_13_radr;
  yt_rsc_7_13_comp_wadr <= yt_rsc_7_13_wadr;

  yt_rsc_7_14_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_7_14_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_7_14_clkr_en,
      d => yt_rsc_7_14_comp_d,
      q => yt_rsc_7_14_comp_q,
      radr => yt_rsc_7_14_comp_radr,
      wadr => yt_rsc_7_14_comp_wadr,
      we => yt_rsc_7_14_we
    );
  yt_rsc_7_14_comp_d <= yt_rsc_7_14_d;
  yt_rsc_7_14_q <= yt_rsc_7_14_comp_q;
  yt_rsc_7_14_comp_radr <= yt_rsc_7_14_radr;
  yt_rsc_7_14_comp_wadr <= yt_rsc_7_14_wadr;

  yt_rsc_7_15_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_7_15_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_7_15_clkr_en,
      d => yt_rsc_7_15_comp_d,
      q => yt_rsc_7_15_comp_q,
      radr => yt_rsc_7_15_comp_radr,
      wadr => yt_rsc_7_15_comp_wadr,
      we => yt_rsc_7_15_we
    );
  yt_rsc_7_15_comp_d <= yt_rsc_7_15_d;
  yt_rsc_7_15_q <= yt_rsc_7_15_comp_q;
  yt_rsc_7_15_comp_radr <= yt_rsc_7_15_radr;
  yt_rsc_7_15_comp_wadr <= yt_rsc_7_15_wadr;

  yt_rsc_7_16_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_7_16_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_7_16_clkr_en,
      d => yt_rsc_7_16_comp_d,
      q => yt_rsc_7_16_comp_q,
      radr => yt_rsc_7_16_comp_radr,
      wadr => yt_rsc_7_16_comp_wadr,
      we => yt_rsc_7_16_we
    );
  yt_rsc_7_16_comp_d <= yt_rsc_7_16_d;
  yt_rsc_7_16_q <= yt_rsc_7_16_comp_q;
  yt_rsc_7_16_comp_radr <= yt_rsc_7_16_radr;
  yt_rsc_7_16_comp_wadr <= yt_rsc_7_16_wadr;

  yt_rsc_7_17_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_7_17_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_7_17_clkr_en,
      d => yt_rsc_7_17_comp_d,
      q => yt_rsc_7_17_comp_q,
      radr => yt_rsc_7_17_comp_radr,
      wadr => yt_rsc_7_17_comp_wadr,
      we => yt_rsc_7_17_we
    );
  yt_rsc_7_17_comp_d <= yt_rsc_7_17_d;
  yt_rsc_7_17_q <= yt_rsc_7_17_comp_q;
  yt_rsc_7_17_comp_radr <= yt_rsc_7_17_radr;
  yt_rsc_7_17_comp_wadr <= yt_rsc_7_17_wadr;

  yt_rsc_7_18_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_7_18_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_7_18_clkr_en,
      d => yt_rsc_7_18_comp_d,
      q => yt_rsc_7_18_comp_q,
      radr => yt_rsc_7_18_comp_radr,
      wadr => yt_rsc_7_18_comp_wadr,
      we => yt_rsc_7_18_we
    );
  yt_rsc_7_18_comp_d <= yt_rsc_7_18_d;
  yt_rsc_7_18_q <= yt_rsc_7_18_comp_q;
  yt_rsc_7_18_comp_radr <= yt_rsc_7_18_radr;
  yt_rsc_7_18_comp_wadr <= yt_rsc_7_18_wadr;

  yt_rsc_7_19_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_7_19_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_7_19_clkr_en,
      d => yt_rsc_7_19_comp_d,
      q => yt_rsc_7_19_comp_q,
      radr => yt_rsc_7_19_comp_radr,
      wadr => yt_rsc_7_19_comp_wadr,
      we => yt_rsc_7_19_we
    );
  yt_rsc_7_19_comp_d <= yt_rsc_7_19_d;
  yt_rsc_7_19_q <= yt_rsc_7_19_comp_q;
  yt_rsc_7_19_comp_radr <= yt_rsc_7_19_radr;
  yt_rsc_7_19_comp_wadr <= yt_rsc_7_19_wadr;

  yt_rsc_7_20_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_7_20_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_7_20_clkr_en,
      d => yt_rsc_7_20_comp_d,
      q => yt_rsc_7_20_comp_q,
      radr => yt_rsc_7_20_comp_radr,
      wadr => yt_rsc_7_20_comp_wadr,
      we => yt_rsc_7_20_we
    );
  yt_rsc_7_20_comp_d <= yt_rsc_7_20_d;
  yt_rsc_7_20_q <= yt_rsc_7_20_comp_q;
  yt_rsc_7_20_comp_radr <= yt_rsc_7_20_radr;
  yt_rsc_7_20_comp_wadr <= yt_rsc_7_20_wadr;

  yt_rsc_7_21_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_7_21_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_7_21_clkr_en,
      d => yt_rsc_7_21_comp_d,
      q => yt_rsc_7_21_comp_q,
      radr => yt_rsc_7_21_comp_radr,
      wadr => yt_rsc_7_21_comp_wadr,
      we => yt_rsc_7_21_we
    );
  yt_rsc_7_21_comp_d <= yt_rsc_7_21_d;
  yt_rsc_7_21_q <= yt_rsc_7_21_comp_q;
  yt_rsc_7_21_comp_radr <= yt_rsc_7_21_radr;
  yt_rsc_7_21_comp_wadr <= yt_rsc_7_21_wadr;

  yt_rsc_7_22_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_7_22_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_7_22_clkr_en,
      d => yt_rsc_7_22_comp_d,
      q => yt_rsc_7_22_comp_q,
      radr => yt_rsc_7_22_comp_radr,
      wadr => yt_rsc_7_22_comp_wadr,
      we => yt_rsc_7_22_we
    );
  yt_rsc_7_22_comp_d <= yt_rsc_7_22_d;
  yt_rsc_7_22_q <= yt_rsc_7_22_comp_q;
  yt_rsc_7_22_comp_radr <= yt_rsc_7_22_radr;
  yt_rsc_7_22_comp_wadr <= yt_rsc_7_22_wadr;

  yt_rsc_7_23_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_7_23_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_7_23_clkr_en,
      d => yt_rsc_7_23_comp_d,
      q => yt_rsc_7_23_comp_q,
      radr => yt_rsc_7_23_comp_radr,
      wadr => yt_rsc_7_23_comp_wadr,
      we => yt_rsc_7_23_we
    );
  yt_rsc_7_23_comp_d <= yt_rsc_7_23_d;
  yt_rsc_7_23_q <= yt_rsc_7_23_comp_q;
  yt_rsc_7_23_comp_radr <= yt_rsc_7_23_radr;
  yt_rsc_7_23_comp_wadr <= yt_rsc_7_23_wadr;

  yt_rsc_7_24_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_7_24_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_7_24_clkr_en,
      d => yt_rsc_7_24_comp_d,
      q => yt_rsc_7_24_comp_q,
      radr => yt_rsc_7_24_comp_radr,
      wadr => yt_rsc_7_24_comp_wadr,
      we => yt_rsc_7_24_we
    );
  yt_rsc_7_24_comp_d <= yt_rsc_7_24_d;
  yt_rsc_7_24_q <= yt_rsc_7_24_comp_q;
  yt_rsc_7_24_comp_radr <= yt_rsc_7_24_radr;
  yt_rsc_7_24_comp_wadr <= yt_rsc_7_24_wadr;

  yt_rsc_7_25_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_7_25_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_7_25_clkr_en,
      d => yt_rsc_7_25_comp_d,
      q => yt_rsc_7_25_comp_q,
      radr => yt_rsc_7_25_comp_radr,
      wadr => yt_rsc_7_25_comp_wadr,
      we => yt_rsc_7_25_we
    );
  yt_rsc_7_25_comp_d <= yt_rsc_7_25_d;
  yt_rsc_7_25_q <= yt_rsc_7_25_comp_q;
  yt_rsc_7_25_comp_radr <= yt_rsc_7_25_radr;
  yt_rsc_7_25_comp_wadr <= yt_rsc_7_25_wadr;

  yt_rsc_7_26_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_7_26_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_7_26_clkr_en,
      d => yt_rsc_7_26_comp_d,
      q => yt_rsc_7_26_comp_q,
      radr => yt_rsc_7_26_comp_radr,
      wadr => yt_rsc_7_26_comp_wadr,
      we => yt_rsc_7_26_we
    );
  yt_rsc_7_26_comp_d <= yt_rsc_7_26_d;
  yt_rsc_7_26_q <= yt_rsc_7_26_comp_q;
  yt_rsc_7_26_comp_radr <= yt_rsc_7_26_radr;
  yt_rsc_7_26_comp_wadr <= yt_rsc_7_26_wadr;

  yt_rsc_7_27_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_7_27_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_7_27_clkr_en,
      d => yt_rsc_7_27_comp_d,
      q => yt_rsc_7_27_comp_q,
      radr => yt_rsc_7_27_comp_radr,
      wadr => yt_rsc_7_27_comp_wadr,
      we => yt_rsc_7_27_we
    );
  yt_rsc_7_27_comp_d <= yt_rsc_7_27_d;
  yt_rsc_7_27_q <= yt_rsc_7_27_comp_q;
  yt_rsc_7_27_comp_radr <= yt_rsc_7_27_radr;
  yt_rsc_7_27_comp_wadr <= yt_rsc_7_27_wadr;

  yt_rsc_7_28_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_7_28_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_7_28_clkr_en,
      d => yt_rsc_7_28_comp_d,
      q => yt_rsc_7_28_comp_q,
      radr => yt_rsc_7_28_comp_radr,
      wadr => yt_rsc_7_28_comp_wadr,
      we => yt_rsc_7_28_we
    );
  yt_rsc_7_28_comp_d <= yt_rsc_7_28_d;
  yt_rsc_7_28_q <= yt_rsc_7_28_comp_q;
  yt_rsc_7_28_comp_radr <= yt_rsc_7_28_radr;
  yt_rsc_7_28_comp_wadr <= yt_rsc_7_28_wadr;

  yt_rsc_7_29_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_7_29_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_7_29_clkr_en,
      d => yt_rsc_7_29_comp_d,
      q => yt_rsc_7_29_comp_q,
      radr => yt_rsc_7_29_comp_radr,
      wadr => yt_rsc_7_29_comp_wadr,
      we => yt_rsc_7_29_we
    );
  yt_rsc_7_29_comp_d <= yt_rsc_7_29_d;
  yt_rsc_7_29_q <= yt_rsc_7_29_comp_q;
  yt_rsc_7_29_comp_radr <= yt_rsc_7_29_radr;
  yt_rsc_7_29_comp_wadr <= yt_rsc_7_29_wadr;

  yt_rsc_7_30_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_7_30_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_7_30_clkr_en,
      d => yt_rsc_7_30_comp_d,
      q => yt_rsc_7_30_comp_q,
      radr => yt_rsc_7_30_comp_radr,
      wadr => yt_rsc_7_30_comp_wadr,
      we => yt_rsc_7_30_we
    );
  yt_rsc_7_30_comp_d <= yt_rsc_7_30_d;
  yt_rsc_7_30_q <= yt_rsc_7_30_comp_q;
  yt_rsc_7_30_comp_radr <= yt_rsc_7_30_radr;
  yt_rsc_7_30_comp_wadr <= yt_rsc_7_30_wadr;

  yt_rsc_7_31_comp : work.block_1r1w_rbw_dual_pkg.BLOCK_1R1W_RBW_DUAL
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      clkr => clk,
      clkr_en => yt_rsc_7_31_clkr_en,
      clkw => clk,
      clkw_en => yt_rsc_7_31_clkr_en,
      d => yt_rsc_7_31_comp_d,
      q => yt_rsc_7_31_comp_q,
      radr => yt_rsc_7_31_comp_radr,
      wadr => yt_rsc_7_31_comp_wadr,
      we => yt_rsc_7_31_we
    );
  yt_rsc_7_31_comp_d <= yt_rsc_7_31_d;
  yt_rsc_7_31_q <= yt_rsc_7_31_comp_q;
  yt_rsc_7_31_comp_radr <= yt_rsc_7_31_radr;
  yt_rsc_7_31_comp_wadr <= yt_rsc_7_31_wadr;

  yt_rsc_0_0_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_7_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_0_0_clkr_en,
      clkw_en => yt_rsc_0_0_clkw_en,
      q => yt_rsc_0_0_i_q,
      radr => yt_rsc_0_0_i_radr,
      we => yt_rsc_0_0_we,
      d => yt_rsc_0_0_i_d,
      wadr => yt_rsc_0_0_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_0_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_0_0_i_clkr_en_d,
      d_d => yt_rsc_0_0_i_d_d,
      q_d => yt_rsc_0_0_i_q_d_1,
      radr_d => yt_rsc_0_0_i_radr_d,
      wadr_d => yt_rsc_0_0_i_wadr_d,
      we_d => yt_rsc_0_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_0_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_0_0_i_q <= yt_rsc_0_0_q;
  yt_rsc_0_0_radr <= yt_rsc_0_0_i_radr;
  yt_rsc_0_0_d <= yt_rsc_0_0_i_d;
  yt_rsc_0_0_wadr <= yt_rsc_0_0_i_wadr;
  yt_rsc_0_0_i_d_d <= yt_rsc_0_0_i_d_d_iff;
  yt_rsc_0_0_i_q_d <= yt_rsc_0_0_i_q_d_1;
  yt_rsc_0_0_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_0_0_i_wadr_d <= yt_rsc_0_0_i_wadr_d_iff;

  yt_rsc_0_1_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_8_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_0_1_clkr_en,
      clkw_en => yt_rsc_0_1_clkw_en,
      q => yt_rsc_0_1_i_q,
      radr => yt_rsc_0_1_i_radr,
      we => yt_rsc_0_1_we,
      d => yt_rsc_0_1_i_d,
      wadr => yt_rsc_0_1_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_0_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_0_0_i_clkr_en_d,
      d_d => yt_rsc_0_1_i_d_d,
      q_d => yt_rsc_0_1_i_q_d_1,
      radr_d => yt_rsc_0_1_i_radr_d,
      wadr_d => yt_rsc_0_1_i_wadr_d,
      we_d => yt_rsc_0_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_0_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_0_1_i_q <= yt_rsc_0_1_q;
  yt_rsc_0_1_radr <= yt_rsc_0_1_i_radr;
  yt_rsc_0_1_d <= yt_rsc_0_1_i_d;
  yt_rsc_0_1_wadr <= yt_rsc_0_1_i_wadr;
  yt_rsc_0_1_i_d_d <= yt_rsc_0_1_i_d_d_iff;
  yt_rsc_0_1_i_q_d <= yt_rsc_0_1_i_q_d_1;
  yt_rsc_0_1_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_0_1_i_wadr_d <= yt_rsc_0_1_i_wadr_d_iff;

  yt_rsc_0_2_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_9_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_0_2_clkr_en,
      clkw_en => yt_rsc_0_2_clkw_en,
      q => yt_rsc_0_2_i_q,
      radr => yt_rsc_0_2_i_radr,
      we => yt_rsc_0_2_we,
      d => yt_rsc_0_2_i_d,
      wadr => yt_rsc_0_2_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_0_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_0_0_i_clkr_en_d,
      d_d => yt_rsc_0_2_i_d_d,
      q_d => yt_rsc_0_2_i_q_d_1,
      radr_d => yt_rsc_0_2_i_radr_d,
      wadr_d => yt_rsc_0_2_i_wadr_d,
      we_d => yt_rsc_0_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_0_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_0_2_i_q <= yt_rsc_0_2_q;
  yt_rsc_0_2_radr <= yt_rsc_0_2_i_radr;
  yt_rsc_0_2_d <= yt_rsc_0_2_i_d;
  yt_rsc_0_2_wadr <= yt_rsc_0_2_i_wadr;
  yt_rsc_0_2_i_d_d <= yt_rsc_0_2_i_d_d_iff;
  yt_rsc_0_2_i_q_d <= yt_rsc_0_2_i_q_d_1;
  yt_rsc_0_2_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_0_2_i_wadr_d <= yt_rsc_0_2_i_wadr_d_iff;

  yt_rsc_0_3_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_10_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_0_3_clkr_en,
      clkw_en => yt_rsc_0_3_clkw_en,
      q => yt_rsc_0_3_i_q,
      radr => yt_rsc_0_3_i_radr,
      we => yt_rsc_0_3_we,
      d => yt_rsc_0_3_i_d,
      wadr => yt_rsc_0_3_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_0_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_0_0_i_clkr_en_d,
      d_d => yt_rsc_0_3_i_d_d,
      q_d => yt_rsc_0_3_i_q_d_1,
      radr_d => yt_rsc_0_3_i_radr_d,
      wadr_d => yt_rsc_0_3_i_wadr_d,
      we_d => yt_rsc_0_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_0_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_0_3_i_q <= yt_rsc_0_3_q;
  yt_rsc_0_3_radr <= yt_rsc_0_3_i_radr;
  yt_rsc_0_3_d <= yt_rsc_0_3_i_d;
  yt_rsc_0_3_wadr <= yt_rsc_0_3_i_wadr;
  yt_rsc_0_3_i_d_d <= yt_rsc_0_3_i_d_d_iff;
  yt_rsc_0_3_i_q_d <= yt_rsc_0_3_i_q_d_1;
  yt_rsc_0_3_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_0_3_i_wadr_d <= yt_rsc_0_3_i_wadr_d_iff;

  yt_rsc_0_4_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_11_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_0_4_clkr_en,
      clkw_en => yt_rsc_0_4_clkw_en,
      q => yt_rsc_0_4_i_q,
      radr => yt_rsc_0_4_i_radr,
      we => yt_rsc_0_4_we,
      d => yt_rsc_0_4_i_d,
      wadr => yt_rsc_0_4_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_0_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_0_0_i_clkr_en_d,
      d_d => yt_rsc_0_4_i_d_d,
      q_d => yt_rsc_0_4_i_q_d_1,
      radr_d => yt_rsc_0_4_i_radr_d,
      wadr_d => yt_rsc_0_4_i_wadr_d,
      we_d => yt_rsc_0_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_0_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_0_4_i_q <= yt_rsc_0_4_q;
  yt_rsc_0_4_radr <= yt_rsc_0_4_i_radr;
  yt_rsc_0_4_d <= yt_rsc_0_4_i_d;
  yt_rsc_0_4_wadr <= yt_rsc_0_4_i_wadr;
  yt_rsc_0_4_i_d_d <= yt_rsc_0_4_i_d_d_iff;
  yt_rsc_0_4_i_q_d <= yt_rsc_0_4_i_q_d_1;
  yt_rsc_0_4_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_0_4_i_wadr_d <= yt_rsc_0_4_i_wadr_d_iff;

  yt_rsc_0_5_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_12_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_0_5_clkr_en,
      clkw_en => yt_rsc_0_5_clkw_en,
      q => yt_rsc_0_5_i_q,
      radr => yt_rsc_0_5_i_radr,
      we => yt_rsc_0_5_we,
      d => yt_rsc_0_5_i_d,
      wadr => yt_rsc_0_5_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_0_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_0_0_i_clkr_en_d,
      d_d => yt_rsc_0_5_i_d_d,
      q_d => yt_rsc_0_5_i_q_d_1,
      radr_d => yt_rsc_0_5_i_radr_d,
      wadr_d => yt_rsc_0_5_i_wadr_d,
      we_d => yt_rsc_0_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_0_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_0_5_i_q <= yt_rsc_0_5_q;
  yt_rsc_0_5_radr <= yt_rsc_0_5_i_radr;
  yt_rsc_0_5_d <= yt_rsc_0_5_i_d;
  yt_rsc_0_5_wadr <= yt_rsc_0_5_i_wadr;
  yt_rsc_0_5_i_d_d <= yt_rsc_0_5_i_d_d_iff;
  yt_rsc_0_5_i_q_d <= yt_rsc_0_5_i_q_d_1;
  yt_rsc_0_5_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_0_5_i_wadr_d <= yt_rsc_0_5_i_wadr_d_iff;

  yt_rsc_0_6_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_13_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_0_6_clkr_en,
      clkw_en => yt_rsc_0_6_clkw_en,
      q => yt_rsc_0_6_i_q,
      radr => yt_rsc_0_6_i_radr,
      we => yt_rsc_0_6_we,
      d => yt_rsc_0_6_i_d,
      wadr => yt_rsc_0_6_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_0_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_0_0_i_clkr_en_d,
      d_d => yt_rsc_0_6_i_d_d,
      q_d => yt_rsc_0_6_i_q_d_1,
      radr_d => yt_rsc_0_6_i_radr_d,
      wadr_d => yt_rsc_0_6_i_wadr_d,
      we_d => yt_rsc_0_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_0_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_0_6_i_q <= yt_rsc_0_6_q;
  yt_rsc_0_6_radr <= yt_rsc_0_6_i_radr;
  yt_rsc_0_6_d <= yt_rsc_0_6_i_d;
  yt_rsc_0_6_wadr <= yt_rsc_0_6_i_wadr;
  yt_rsc_0_6_i_d_d <= yt_rsc_0_6_i_d_d_iff;
  yt_rsc_0_6_i_q_d <= yt_rsc_0_6_i_q_d_1;
  yt_rsc_0_6_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_0_6_i_wadr_d <= yt_rsc_0_6_i_wadr_d_iff;

  yt_rsc_0_7_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_14_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_0_7_clkr_en,
      clkw_en => yt_rsc_0_7_clkw_en,
      q => yt_rsc_0_7_i_q,
      radr => yt_rsc_0_7_i_radr,
      we => yt_rsc_0_7_we,
      d => yt_rsc_0_7_i_d,
      wadr => yt_rsc_0_7_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_0_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_0_0_i_clkr_en_d,
      d_d => yt_rsc_0_7_i_d_d,
      q_d => yt_rsc_0_7_i_q_d_1,
      radr_d => yt_rsc_0_7_i_radr_d,
      wadr_d => yt_rsc_0_7_i_wadr_d,
      we_d => yt_rsc_0_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_0_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_0_7_i_q <= yt_rsc_0_7_q;
  yt_rsc_0_7_radr <= yt_rsc_0_7_i_radr;
  yt_rsc_0_7_d <= yt_rsc_0_7_i_d;
  yt_rsc_0_7_wadr <= yt_rsc_0_7_i_wadr;
  yt_rsc_0_7_i_d_d <= yt_rsc_0_7_i_d_d_iff;
  yt_rsc_0_7_i_q_d <= yt_rsc_0_7_i_q_d_1;
  yt_rsc_0_7_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_0_7_i_wadr_d <= yt_rsc_0_0_i_wadr_d_iff;

  yt_rsc_0_8_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_15_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_0_8_clkr_en,
      clkw_en => yt_rsc_0_8_clkw_en,
      q => yt_rsc_0_8_i_q,
      radr => yt_rsc_0_8_i_radr,
      we => yt_rsc_0_8_we,
      d => yt_rsc_0_8_i_d,
      wadr => yt_rsc_0_8_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_0_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_0_0_i_clkr_en_d,
      d_d => yt_rsc_0_8_i_d_d,
      q_d => yt_rsc_0_8_i_q_d_1,
      radr_d => yt_rsc_0_8_i_radr_d,
      wadr_d => yt_rsc_0_8_i_wadr_d,
      we_d => yt_rsc_0_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_0_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_0_8_i_q <= yt_rsc_0_8_q;
  yt_rsc_0_8_radr <= yt_rsc_0_8_i_radr;
  yt_rsc_0_8_d <= yt_rsc_0_8_i_d;
  yt_rsc_0_8_wadr <= yt_rsc_0_8_i_wadr;
  yt_rsc_0_8_i_d_d <= yt_rsc_0_8_i_d_d_iff;
  yt_rsc_0_8_i_q_d <= yt_rsc_0_8_i_q_d_1;
  yt_rsc_0_8_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_0_8_i_wadr_d <= yt_rsc_0_1_i_wadr_d_iff;

  yt_rsc_0_9_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_16_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_0_9_clkr_en,
      clkw_en => yt_rsc_0_9_clkw_en,
      q => yt_rsc_0_9_i_q,
      radr => yt_rsc_0_9_i_radr,
      we => yt_rsc_0_9_we,
      d => yt_rsc_0_9_i_d,
      wadr => yt_rsc_0_9_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_0_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_0_0_i_clkr_en_d,
      d_d => yt_rsc_0_9_i_d_d,
      q_d => yt_rsc_0_9_i_q_d_1,
      radr_d => yt_rsc_0_9_i_radr_d,
      wadr_d => yt_rsc_0_9_i_wadr_d,
      we_d => yt_rsc_0_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_0_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_0_9_i_q <= yt_rsc_0_9_q;
  yt_rsc_0_9_radr <= yt_rsc_0_9_i_radr;
  yt_rsc_0_9_d <= yt_rsc_0_9_i_d;
  yt_rsc_0_9_wadr <= yt_rsc_0_9_i_wadr;
  yt_rsc_0_9_i_d_d <= yt_rsc_0_9_i_d_d_iff;
  yt_rsc_0_9_i_q_d <= yt_rsc_0_9_i_q_d_1;
  yt_rsc_0_9_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_0_9_i_wadr_d <= yt_rsc_0_2_i_wadr_d_iff;

  yt_rsc_0_10_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_17_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_0_10_clkr_en,
      clkw_en => yt_rsc_0_10_clkw_en,
      q => yt_rsc_0_10_i_q,
      radr => yt_rsc_0_10_i_radr,
      we => yt_rsc_0_10_we,
      d => yt_rsc_0_10_i_d,
      wadr => yt_rsc_0_10_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_0_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_0_0_i_clkr_en_d,
      d_d => yt_rsc_0_10_i_d_d,
      q_d => yt_rsc_0_10_i_q_d_1,
      radr_d => yt_rsc_0_10_i_radr_d,
      wadr_d => yt_rsc_0_10_i_wadr_d,
      we_d => yt_rsc_0_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_0_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_0_10_i_q <= yt_rsc_0_10_q;
  yt_rsc_0_10_radr <= yt_rsc_0_10_i_radr;
  yt_rsc_0_10_d <= yt_rsc_0_10_i_d;
  yt_rsc_0_10_wadr <= yt_rsc_0_10_i_wadr;
  yt_rsc_0_10_i_d_d <= yt_rsc_0_10_i_d_d_iff;
  yt_rsc_0_10_i_q_d <= yt_rsc_0_10_i_q_d_1;
  yt_rsc_0_10_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_0_10_i_wadr_d <= yt_rsc_0_10_i_wadr_d_iff;

  yt_rsc_0_11_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_18_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_0_11_clkr_en,
      clkw_en => yt_rsc_0_11_clkw_en,
      q => yt_rsc_0_11_i_q,
      radr => yt_rsc_0_11_i_radr,
      we => yt_rsc_0_11_we,
      d => yt_rsc_0_11_i_d,
      wadr => yt_rsc_0_11_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_0_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_0_0_i_clkr_en_d,
      d_d => yt_rsc_0_11_i_d_d,
      q_d => yt_rsc_0_11_i_q_d_1,
      radr_d => yt_rsc_0_11_i_radr_d,
      wadr_d => yt_rsc_0_11_i_wadr_d,
      we_d => yt_rsc_0_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_0_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_0_11_i_q <= yt_rsc_0_11_q;
  yt_rsc_0_11_radr <= yt_rsc_0_11_i_radr;
  yt_rsc_0_11_d <= yt_rsc_0_11_i_d;
  yt_rsc_0_11_wadr <= yt_rsc_0_11_i_wadr;
  yt_rsc_0_11_i_d_d <= yt_rsc_0_11_i_d_d_iff;
  yt_rsc_0_11_i_q_d <= yt_rsc_0_11_i_q_d_1;
  yt_rsc_0_11_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_0_11_i_wadr_d <= yt_rsc_0_11_i_wadr_d_iff;

  yt_rsc_0_12_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_19_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_0_12_clkr_en,
      clkw_en => yt_rsc_0_12_clkw_en,
      q => yt_rsc_0_12_i_q,
      radr => yt_rsc_0_12_i_radr,
      we => yt_rsc_0_12_we,
      d => yt_rsc_0_12_i_d,
      wadr => yt_rsc_0_12_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_0_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_0_0_i_clkr_en_d,
      d_d => yt_rsc_0_12_i_d_d,
      q_d => yt_rsc_0_12_i_q_d_1,
      radr_d => yt_rsc_0_12_i_radr_d,
      wadr_d => yt_rsc_0_12_i_wadr_d,
      we_d => yt_rsc_0_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_0_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_0_12_i_q <= yt_rsc_0_12_q;
  yt_rsc_0_12_radr <= yt_rsc_0_12_i_radr;
  yt_rsc_0_12_d <= yt_rsc_0_12_i_d;
  yt_rsc_0_12_wadr <= yt_rsc_0_12_i_wadr;
  yt_rsc_0_12_i_d_d <= yt_rsc_0_12_i_d_d_iff;
  yt_rsc_0_12_i_q_d <= yt_rsc_0_12_i_q_d_1;
  yt_rsc_0_12_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_0_12_i_wadr_d <= yt_rsc_0_3_i_wadr_d_iff;

  yt_rsc_0_13_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_20_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_0_13_clkr_en,
      clkw_en => yt_rsc_0_13_clkw_en,
      q => yt_rsc_0_13_i_q,
      radr => yt_rsc_0_13_i_radr,
      we => yt_rsc_0_13_we,
      d => yt_rsc_0_13_i_d,
      wadr => yt_rsc_0_13_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_0_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_0_0_i_clkr_en_d,
      d_d => yt_rsc_0_13_i_d_d,
      q_d => yt_rsc_0_13_i_q_d_1,
      radr_d => yt_rsc_0_13_i_radr_d,
      wadr_d => yt_rsc_0_13_i_wadr_d,
      we_d => yt_rsc_0_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_0_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_0_13_i_q <= yt_rsc_0_13_q;
  yt_rsc_0_13_radr <= yt_rsc_0_13_i_radr;
  yt_rsc_0_13_d <= yt_rsc_0_13_i_d;
  yt_rsc_0_13_wadr <= yt_rsc_0_13_i_wadr;
  yt_rsc_0_13_i_d_d <= yt_rsc_0_13_i_d_d_iff;
  yt_rsc_0_13_i_q_d <= yt_rsc_0_13_i_q_d_1;
  yt_rsc_0_13_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_0_13_i_wadr_d <= yt_rsc_0_4_i_wadr_d_iff;

  yt_rsc_0_14_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_21_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_0_14_clkr_en,
      clkw_en => yt_rsc_0_14_clkw_en,
      q => yt_rsc_0_14_i_q,
      radr => yt_rsc_0_14_i_radr,
      we => yt_rsc_0_14_we,
      d => yt_rsc_0_14_i_d,
      wadr => yt_rsc_0_14_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_0_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_0_0_i_clkr_en_d,
      d_d => yt_rsc_0_14_i_d_d,
      q_d => yt_rsc_0_14_i_q_d_1,
      radr_d => yt_rsc_0_14_i_radr_d,
      wadr_d => yt_rsc_0_14_i_wadr_d,
      we_d => yt_rsc_0_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_0_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_0_14_i_q <= yt_rsc_0_14_q;
  yt_rsc_0_14_radr <= yt_rsc_0_14_i_radr;
  yt_rsc_0_14_d <= yt_rsc_0_14_i_d;
  yt_rsc_0_14_wadr <= yt_rsc_0_14_i_wadr;
  yt_rsc_0_14_i_d_d <= yt_rsc_0_14_i_d_d_iff;
  yt_rsc_0_14_i_q_d <= yt_rsc_0_14_i_q_d_1;
  yt_rsc_0_14_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_0_14_i_wadr_d <= yt_rsc_0_5_i_wadr_d_iff;

  yt_rsc_0_15_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_22_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_0_15_clkr_en,
      clkw_en => yt_rsc_0_15_clkw_en,
      q => yt_rsc_0_15_i_q,
      radr => yt_rsc_0_15_i_radr,
      we => yt_rsc_0_15_we,
      d => yt_rsc_0_15_i_d,
      wadr => yt_rsc_0_15_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_0_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_0_0_i_clkr_en_d,
      d_d => yt_rsc_0_15_i_d_d,
      q_d => yt_rsc_0_15_i_q_d_1,
      radr_d => yt_rsc_0_15_i_radr_d,
      wadr_d => yt_rsc_0_15_i_wadr_d,
      we_d => yt_rsc_0_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_0_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_0_15_i_q <= yt_rsc_0_15_q;
  yt_rsc_0_15_radr <= yt_rsc_0_15_i_radr;
  yt_rsc_0_15_d <= yt_rsc_0_15_i_d;
  yt_rsc_0_15_wadr <= yt_rsc_0_15_i_wadr;
  yt_rsc_0_15_i_d_d <= yt_rsc_0_15_i_d_d_iff;
  yt_rsc_0_15_i_q_d <= yt_rsc_0_15_i_q_d_1;
  yt_rsc_0_15_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_0_15_i_wadr_d <= yt_rsc_0_6_i_wadr_d_iff;

  yt_rsc_0_16_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_23_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_0_16_clkr_en,
      clkw_en => yt_rsc_0_16_clkw_en,
      q => yt_rsc_0_16_i_q,
      radr => yt_rsc_0_16_i_radr,
      we => yt_rsc_0_16_we,
      d => yt_rsc_0_16_i_d,
      wadr => yt_rsc_0_16_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_0_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_0_16_i_clkr_en_d,
      d_d => yt_rsc_0_16_i_d_d,
      q_d => yt_rsc_0_16_i_q_d_1,
      radr_d => yt_rsc_0_16_i_radr_d,
      wadr_d => yt_rsc_0_16_i_wadr_d,
      we_d => yt_rsc_0_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_0_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_0_16_i_q <= yt_rsc_0_16_q;
  yt_rsc_0_16_radr <= yt_rsc_0_16_i_radr;
  yt_rsc_0_16_d <= yt_rsc_0_16_i_d;
  yt_rsc_0_16_wadr <= yt_rsc_0_16_i_wadr;
  yt_rsc_0_16_i_d_d <= yt_rsc_0_0_i_d_d_iff;
  yt_rsc_0_16_i_q_d <= yt_rsc_0_16_i_q_d_1;
  yt_rsc_0_16_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_0_16_i_wadr_d <= yt_rsc_0_0_i_wadr_d_iff;

  yt_rsc_0_17_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_24_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_0_17_clkr_en,
      clkw_en => yt_rsc_0_17_clkw_en,
      q => yt_rsc_0_17_i_q,
      radr => yt_rsc_0_17_i_radr,
      we => yt_rsc_0_17_we,
      d => yt_rsc_0_17_i_d,
      wadr => yt_rsc_0_17_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_0_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_0_16_i_clkr_en_d,
      d_d => yt_rsc_0_17_i_d_d,
      q_d => yt_rsc_0_17_i_q_d_1,
      radr_d => yt_rsc_0_17_i_radr_d,
      wadr_d => yt_rsc_0_17_i_wadr_d,
      we_d => yt_rsc_0_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_0_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_0_17_i_q <= yt_rsc_0_17_q;
  yt_rsc_0_17_radr <= yt_rsc_0_17_i_radr;
  yt_rsc_0_17_d <= yt_rsc_0_17_i_d;
  yt_rsc_0_17_wadr <= yt_rsc_0_17_i_wadr;
  yt_rsc_0_17_i_d_d <= yt_rsc_0_1_i_d_d_iff;
  yt_rsc_0_17_i_q_d <= yt_rsc_0_17_i_q_d_1;
  yt_rsc_0_17_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_0_17_i_wadr_d <= yt_rsc_0_1_i_wadr_d_iff;

  yt_rsc_0_18_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_25_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_0_18_clkr_en,
      clkw_en => yt_rsc_0_18_clkw_en,
      q => yt_rsc_0_18_i_q,
      radr => yt_rsc_0_18_i_radr,
      we => yt_rsc_0_18_we,
      d => yt_rsc_0_18_i_d,
      wadr => yt_rsc_0_18_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_0_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_0_16_i_clkr_en_d,
      d_d => yt_rsc_0_18_i_d_d,
      q_d => yt_rsc_0_18_i_q_d_1,
      radr_d => yt_rsc_0_18_i_radr_d,
      wadr_d => yt_rsc_0_18_i_wadr_d,
      we_d => yt_rsc_0_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_0_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_0_18_i_q <= yt_rsc_0_18_q;
  yt_rsc_0_18_radr <= yt_rsc_0_18_i_radr;
  yt_rsc_0_18_d <= yt_rsc_0_18_i_d;
  yt_rsc_0_18_wadr <= yt_rsc_0_18_i_wadr;
  yt_rsc_0_18_i_d_d <= yt_rsc_0_2_i_d_d_iff;
  yt_rsc_0_18_i_q_d <= yt_rsc_0_18_i_q_d_1;
  yt_rsc_0_18_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_0_18_i_wadr_d <= yt_rsc_0_2_i_wadr_d_iff;

  yt_rsc_0_19_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_26_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_0_19_clkr_en,
      clkw_en => yt_rsc_0_19_clkw_en,
      q => yt_rsc_0_19_i_q,
      radr => yt_rsc_0_19_i_radr,
      we => yt_rsc_0_19_we,
      d => yt_rsc_0_19_i_d,
      wadr => yt_rsc_0_19_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_0_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_0_16_i_clkr_en_d,
      d_d => yt_rsc_0_19_i_d_d,
      q_d => yt_rsc_0_19_i_q_d_1,
      radr_d => yt_rsc_0_19_i_radr_d,
      wadr_d => yt_rsc_0_19_i_wadr_d,
      we_d => yt_rsc_0_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_0_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_0_19_i_q <= yt_rsc_0_19_q;
  yt_rsc_0_19_radr <= yt_rsc_0_19_i_radr;
  yt_rsc_0_19_d <= yt_rsc_0_19_i_d;
  yt_rsc_0_19_wadr <= yt_rsc_0_19_i_wadr;
  yt_rsc_0_19_i_d_d <= yt_rsc_0_3_i_d_d_iff;
  yt_rsc_0_19_i_q_d <= yt_rsc_0_19_i_q_d_1;
  yt_rsc_0_19_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_0_19_i_wadr_d <= yt_rsc_0_3_i_wadr_d_iff;

  yt_rsc_0_20_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_27_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_0_20_clkr_en,
      clkw_en => yt_rsc_0_20_clkw_en,
      q => yt_rsc_0_20_i_q,
      radr => yt_rsc_0_20_i_radr,
      we => yt_rsc_0_20_we,
      d => yt_rsc_0_20_i_d,
      wadr => yt_rsc_0_20_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_0_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_0_16_i_clkr_en_d,
      d_d => yt_rsc_0_20_i_d_d,
      q_d => yt_rsc_0_20_i_q_d_1,
      radr_d => yt_rsc_0_20_i_radr_d,
      wadr_d => yt_rsc_0_20_i_wadr_d,
      we_d => yt_rsc_0_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_0_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_0_20_i_q <= yt_rsc_0_20_q;
  yt_rsc_0_20_radr <= yt_rsc_0_20_i_radr;
  yt_rsc_0_20_d <= yt_rsc_0_20_i_d;
  yt_rsc_0_20_wadr <= yt_rsc_0_20_i_wadr;
  yt_rsc_0_20_i_d_d <= yt_rsc_0_4_i_d_d_iff;
  yt_rsc_0_20_i_q_d <= yt_rsc_0_20_i_q_d_1;
  yt_rsc_0_20_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_0_20_i_wadr_d <= yt_rsc_0_4_i_wadr_d_iff;

  yt_rsc_0_21_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_28_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_0_21_clkr_en,
      clkw_en => yt_rsc_0_21_clkw_en,
      q => yt_rsc_0_21_i_q,
      radr => yt_rsc_0_21_i_radr,
      we => yt_rsc_0_21_we,
      d => yt_rsc_0_21_i_d,
      wadr => yt_rsc_0_21_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_0_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_0_16_i_clkr_en_d,
      d_d => yt_rsc_0_21_i_d_d,
      q_d => yt_rsc_0_21_i_q_d_1,
      radr_d => yt_rsc_0_21_i_radr_d,
      wadr_d => yt_rsc_0_21_i_wadr_d,
      we_d => yt_rsc_0_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_0_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_0_21_i_q <= yt_rsc_0_21_q;
  yt_rsc_0_21_radr <= yt_rsc_0_21_i_radr;
  yt_rsc_0_21_d <= yt_rsc_0_21_i_d;
  yt_rsc_0_21_wadr <= yt_rsc_0_21_i_wadr;
  yt_rsc_0_21_i_d_d <= yt_rsc_0_5_i_d_d_iff;
  yt_rsc_0_21_i_q_d <= yt_rsc_0_21_i_q_d_1;
  yt_rsc_0_21_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_0_21_i_wadr_d <= yt_rsc_0_5_i_wadr_d_iff;

  yt_rsc_0_22_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_29_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_0_22_clkr_en,
      clkw_en => yt_rsc_0_22_clkw_en,
      q => yt_rsc_0_22_i_q,
      radr => yt_rsc_0_22_i_radr,
      we => yt_rsc_0_22_we,
      d => yt_rsc_0_22_i_d,
      wadr => yt_rsc_0_22_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_0_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_0_16_i_clkr_en_d,
      d_d => yt_rsc_0_22_i_d_d,
      q_d => yt_rsc_0_22_i_q_d_1,
      radr_d => yt_rsc_0_22_i_radr_d,
      wadr_d => yt_rsc_0_22_i_wadr_d,
      we_d => yt_rsc_0_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_0_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_0_22_i_q <= yt_rsc_0_22_q;
  yt_rsc_0_22_radr <= yt_rsc_0_22_i_radr;
  yt_rsc_0_22_d <= yt_rsc_0_22_i_d;
  yt_rsc_0_22_wadr <= yt_rsc_0_22_i_wadr;
  yt_rsc_0_22_i_d_d <= yt_rsc_0_6_i_d_d_iff;
  yt_rsc_0_22_i_q_d <= yt_rsc_0_22_i_q_d_1;
  yt_rsc_0_22_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_0_22_i_wadr_d <= yt_rsc_0_6_i_wadr_d_iff;

  yt_rsc_0_23_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_30_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_0_23_clkr_en,
      clkw_en => yt_rsc_0_23_clkw_en,
      q => yt_rsc_0_23_i_q,
      radr => yt_rsc_0_23_i_radr,
      we => yt_rsc_0_23_we,
      d => yt_rsc_0_23_i_d,
      wadr => yt_rsc_0_23_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_0_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_0_16_i_clkr_en_d,
      d_d => yt_rsc_0_23_i_d_d,
      q_d => yt_rsc_0_23_i_q_d_1,
      radr_d => yt_rsc_0_23_i_radr_d,
      wadr_d => yt_rsc_0_23_i_wadr_d,
      we_d => yt_rsc_0_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_0_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_0_23_i_q <= yt_rsc_0_23_q;
  yt_rsc_0_23_radr <= yt_rsc_0_23_i_radr;
  yt_rsc_0_23_d <= yt_rsc_0_23_i_d;
  yt_rsc_0_23_wadr <= yt_rsc_0_23_i_wadr;
  yt_rsc_0_23_i_d_d <= yt_rsc_0_7_i_d_d_iff;
  yt_rsc_0_23_i_q_d <= yt_rsc_0_23_i_q_d_1;
  yt_rsc_0_23_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_0_23_i_wadr_d <= yt_rsc_0_0_i_wadr_d_iff;

  yt_rsc_0_24_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_31_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_0_24_clkr_en,
      clkw_en => yt_rsc_0_24_clkw_en,
      q => yt_rsc_0_24_i_q,
      radr => yt_rsc_0_24_i_radr,
      we => yt_rsc_0_24_we,
      d => yt_rsc_0_24_i_d,
      wadr => yt_rsc_0_24_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_0_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_0_16_i_clkr_en_d,
      d_d => yt_rsc_0_24_i_d_d,
      q_d => yt_rsc_0_24_i_q_d_1,
      radr_d => yt_rsc_0_24_i_radr_d,
      wadr_d => yt_rsc_0_24_i_wadr_d,
      we_d => yt_rsc_0_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_0_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_0_24_i_q <= yt_rsc_0_24_q;
  yt_rsc_0_24_radr <= yt_rsc_0_24_i_radr;
  yt_rsc_0_24_d <= yt_rsc_0_24_i_d;
  yt_rsc_0_24_wadr <= yt_rsc_0_24_i_wadr;
  yt_rsc_0_24_i_d_d <= yt_rsc_0_8_i_d_d_iff;
  yt_rsc_0_24_i_q_d <= yt_rsc_0_24_i_q_d_1;
  yt_rsc_0_24_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_0_24_i_wadr_d <= yt_rsc_0_1_i_wadr_d_iff;

  yt_rsc_0_25_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_32_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_0_25_clkr_en,
      clkw_en => yt_rsc_0_25_clkw_en,
      q => yt_rsc_0_25_i_q,
      radr => yt_rsc_0_25_i_radr,
      we => yt_rsc_0_25_we,
      d => yt_rsc_0_25_i_d,
      wadr => yt_rsc_0_25_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_0_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_0_16_i_clkr_en_d,
      d_d => yt_rsc_0_25_i_d_d,
      q_d => yt_rsc_0_25_i_q_d_1,
      radr_d => yt_rsc_0_25_i_radr_d,
      wadr_d => yt_rsc_0_25_i_wadr_d,
      we_d => yt_rsc_0_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_0_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_0_25_i_q <= yt_rsc_0_25_q;
  yt_rsc_0_25_radr <= yt_rsc_0_25_i_radr;
  yt_rsc_0_25_d <= yt_rsc_0_25_i_d;
  yt_rsc_0_25_wadr <= yt_rsc_0_25_i_wadr;
  yt_rsc_0_25_i_d_d <= yt_rsc_0_9_i_d_d_iff;
  yt_rsc_0_25_i_q_d <= yt_rsc_0_25_i_q_d_1;
  yt_rsc_0_25_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_0_25_i_wadr_d <= yt_rsc_0_2_i_wadr_d_iff;

  yt_rsc_0_26_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_33_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_0_26_clkr_en,
      clkw_en => yt_rsc_0_26_clkw_en,
      q => yt_rsc_0_26_i_q,
      radr => yt_rsc_0_26_i_radr,
      we => yt_rsc_0_26_we,
      d => yt_rsc_0_26_i_d,
      wadr => yt_rsc_0_26_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_0_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_0_16_i_clkr_en_d,
      d_d => yt_rsc_0_26_i_d_d,
      q_d => yt_rsc_0_26_i_q_d_1,
      radr_d => yt_rsc_0_26_i_radr_d,
      wadr_d => yt_rsc_0_26_i_wadr_d,
      we_d => yt_rsc_0_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_0_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_0_26_i_q <= yt_rsc_0_26_q;
  yt_rsc_0_26_radr <= yt_rsc_0_26_i_radr;
  yt_rsc_0_26_d <= yt_rsc_0_26_i_d;
  yt_rsc_0_26_wadr <= yt_rsc_0_26_i_wadr;
  yt_rsc_0_26_i_d_d <= yt_rsc_0_10_i_d_d_iff;
  yt_rsc_0_26_i_q_d <= yt_rsc_0_26_i_q_d_1;
  yt_rsc_0_26_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_0_26_i_wadr_d <= yt_rsc_0_10_i_wadr_d_iff;

  yt_rsc_0_27_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_34_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_0_27_clkr_en,
      clkw_en => yt_rsc_0_27_clkw_en,
      q => yt_rsc_0_27_i_q,
      radr => yt_rsc_0_27_i_radr,
      we => yt_rsc_0_27_we,
      d => yt_rsc_0_27_i_d,
      wadr => yt_rsc_0_27_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_0_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_0_16_i_clkr_en_d,
      d_d => yt_rsc_0_27_i_d_d,
      q_d => yt_rsc_0_27_i_q_d_1,
      radr_d => yt_rsc_0_27_i_radr_d,
      wadr_d => yt_rsc_0_27_i_wadr_d,
      we_d => yt_rsc_0_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_0_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_0_27_i_q <= yt_rsc_0_27_q;
  yt_rsc_0_27_radr <= yt_rsc_0_27_i_radr;
  yt_rsc_0_27_d <= yt_rsc_0_27_i_d;
  yt_rsc_0_27_wadr <= yt_rsc_0_27_i_wadr;
  yt_rsc_0_27_i_d_d <= yt_rsc_0_11_i_d_d_iff;
  yt_rsc_0_27_i_q_d <= yt_rsc_0_27_i_q_d_1;
  yt_rsc_0_27_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_0_27_i_wadr_d <= yt_rsc_0_11_i_wadr_d_iff;

  yt_rsc_0_28_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_35_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_0_28_clkr_en,
      clkw_en => yt_rsc_0_28_clkw_en,
      q => yt_rsc_0_28_i_q,
      radr => yt_rsc_0_28_i_radr,
      we => yt_rsc_0_28_we,
      d => yt_rsc_0_28_i_d,
      wadr => yt_rsc_0_28_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_0_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_0_16_i_clkr_en_d,
      d_d => yt_rsc_0_28_i_d_d,
      q_d => yt_rsc_0_28_i_q_d_1,
      radr_d => yt_rsc_0_28_i_radr_d,
      wadr_d => yt_rsc_0_28_i_wadr_d,
      we_d => yt_rsc_0_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_0_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_0_28_i_q <= yt_rsc_0_28_q;
  yt_rsc_0_28_radr <= yt_rsc_0_28_i_radr;
  yt_rsc_0_28_d <= yt_rsc_0_28_i_d;
  yt_rsc_0_28_wadr <= yt_rsc_0_28_i_wadr;
  yt_rsc_0_28_i_d_d <= yt_rsc_0_12_i_d_d_iff;
  yt_rsc_0_28_i_q_d <= yt_rsc_0_28_i_q_d_1;
  yt_rsc_0_28_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_0_28_i_wadr_d <= yt_rsc_0_3_i_wadr_d_iff;

  yt_rsc_0_29_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_36_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_0_29_clkr_en,
      clkw_en => yt_rsc_0_29_clkw_en,
      q => yt_rsc_0_29_i_q,
      radr => yt_rsc_0_29_i_radr,
      we => yt_rsc_0_29_we,
      d => yt_rsc_0_29_i_d,
      wadr => yt_rsc_0_29_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_0_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_0_16_i_clkr_en_d,
      d_d => yt_rsc_0_29_i_d_d,
      q_d => yt_rsc_0_29_i_q_d_1,
      radr_d => yt_rsc_0_29_i_radr_d,
      wadr_d => yt_rsc_0_29_i_wadr_d,
      we_d => yt_rsc_0_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_0_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_0_29_i_q <= yt_rsc_0_29_q;
  yt_rsc_0_29_radr <= yt_rsc_0_29_i_radr;
  yt_rsc_0_29_d <= yt_rsc_0_29_i_d;
  yt_rsc_0_29_wadr <= yt_rsc_0_29_i_wadr;
  yt_rsc_0_29_i_d_d <= yt_rsc_0_13_i_d_d_iff;
  yt_rsc_0_29_i_q_d <= yt_rsc_0_29_i_q_d_1;
  yt_rsc_0_29_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_0_29_i_wadr_d <= yt_rsc_0_4_i_wadr_d_iff;

  yt_rsc_0_30_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_37_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_0_30_clkr_en,
      clkw_en => yt_rsc_0_30_clkw_en,
      q => yt_rsc_0_30_i_q,
      radr => yt_rsc_0_30_i_radr,
      we => yt_rsc_0_30_we,
      d => yt_rsc_0_30_i_d,
      wadr => yt_rsc_0_30_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_0_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_0_16_i_clkr_en_d,
      d_d => yt_rsc_0_30_i_d_d,
      q_d => yt_rsc_0_30_i_q_d_1,
      radr_d => yt_rsc_0_30_i_radr_d,
      wadr_d => yt_rsc_0_30_i_wadr_d,
      we_d => yt_rsc_0_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_0_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_0_30_i_q <= yt_rsc_0_30_q;
  yt_rsc_0_30_radr <= yt_rsc_0_30_i_radr;
  yt_rsc_0_30_d <= yt_rsc_0_30_i_d;
  yt_rsc_0_30_wadr <= yt_rsc_0_30_i_wadr;
  yt_rsc_0_30_i_d_d <= yt_rsc_0_14_i_d_d_iff;
  yt_rsc_0_30_i_q_d <= yt_rsc_0_30_i_q_d_1;
  yt_rsc_0_30_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_0_30_i_wadr_d <= yt_rsc_0_5_i_wadr_d_iff;

  yt_rsc_0_31_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_38_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_0_31_clkr_en,
      clkw_en => yt_rsc_0_31_clkw_en,
      q => yt_rsc_0_31_i_q,
      radr => yt_rsc_0_31_i_radr,
      we => yt_rsc_0_31_we,
      d => yt_rsc_0_31_i_d,
      wadr => yt_rsc_0_31_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_0_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_0_16_i_clkr_en_d,
      d_d => yt_rsc_0_31_i_d_d,
      q_d => yt_rsc_0_31_i_q_d_1,
      radr_d => yt_rsc_0_31_i_radr_d,
      wadr_d => yt_rsc_0_31_i_wadr_d,
      we_d => yt_rsc_0_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_0_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_0_31_i_q <= yt_rsc_0_31_q;
  yt_rsc_0_31_radr <= yt_rsc_0_31_i_radr;
  yt_rsc_0_31_d <= yt_rsc_0_31_i_d;
  yt_rsc_0_31_wadr <= yt_rsc_0_31_i_wadr;
  yt_rsc_0_31_i_d_d <= yt_rsc_0_15_i_d_d_iff;
  yt_rsc_0_31_i_q_d <= yt_rsc_0_31_i_q_d_1;
  yt_rsc_0_31_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_0_31_i_wadr_d <= yt_rsc_0_6_i_wadr_d_iff;

  yt_rsc_1_0_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_39_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_1_0_clkr_en,
      clkw_en => yt_rsc_1_0_clkw_en,
      q => yt_rsc_1_0_i_q,
      radr => yt_rsc_1_0_i_radr,
      we => yt_rsc_1_0_we,
      d => yt_rsc_1_0_i_d,
      wadr => yt_rsc_1_0_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_1_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_1_0_i_clkr_en_d,
      d_d => yt_rsc_1_0_i_d_d,
      q_d => yt_rsc_1_0_i_q_d_1,
      radr_d => yt_rsc_1_0_i_radr_d,
      wadr_d => yt_rsc_1_0_i_wadr_d,
      we_d => yt_rsc_1_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_1_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_1_0_i_q <= yt_rsc_1_0_q;
  yt_rsc_1_0_radr <= yt_rsc_1_0_i_radr;
  yt_rsc_1_0_d <= yt_rsc_1_0_i_d;
  yt_rsc_1_0_wadr <= yt_rsc_1_0_i_wadr;
  yt_rsc_1_0_i_d_d <= yt_rsc_0_0_i_d_d_iff;
  yt_rsc_1_0_i_q_d <= yt_rsc_1_0_i_q_d_1;
  yt_rsc_1_0_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_1_0_i_wadr_d <= yt_rsc_0_0_i_wadr_d_iff;

  yt_rsc_1_1_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_40_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_1_1_clkr_en,
      clkw_en => yt_rsc_1_1_clkw_en,
      q => yt_rsc_1_1_i_q,
      radr => yt_rsc_1_1_i_radr,
      we => yt_rsc_1_1_we,
      d => yt_rsc_1_1_i_d,
      wadr => yt_rsc_1_1_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_1_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_1_0_i_clkr_en_d,
      d_d => yt_rsc_1_1_i_d_d,
      q_d => yt_rsc_1_1_i_q_d_1,
      radr_d => yt_rsc_1_1_i_radr_d,
      wadr_d => yt_rsc_1_1_i_wadr_d,
      we_d => yt_rsc_1_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_1_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_1_1_i_q <= yt_rsc_1_1_q;
  yt_rsc_1_1_radr <= yt_rsc_1_1_i_radr;
  yt_rsc_1_1_d <= yt_rsc_1_1_i_d;
  yt_rsc_1_1_wadr <= yt_rsc_1_1_i_wadr;
  yt_rsc_1_1_i_d_d <= yt_rsc_0_1_i_d_d_iff;
  yt_rsc_1_1_i_q_d <= yt_rsc_1_1_i_q_d_1;
  yt_rsc_1_1_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_1_1_i_wadr_d <= yt_rsc_0_1_i_wadr_d_iff;

  yt_rsc_1_2_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_41_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_1_2_clkr_en,
      clkw_en => yt_rsc_1_2_clkw_en,
      q => yt_rsc_1_2_i_q,
      radr => yt_rsc_1_2_i_radr,
      we => yt_rsc_1_2_we,
      d => yt_rsc_1_2_i_d,
      wadr => yt_rsc_1_2_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_1_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_1_0_i_clkr_en_d,
      d_d => yt_rsc_1_2_i_d_d,
      q_d => yt_rsc_1_2_i_q_d_1,
      radr_d => yt_rsc_1_2_i_radr_d,
      wadr_d => yt_rsc_1_2_i_wadr_d,
      we_d => yt_rsc_1_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_1_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_1_2_i_q <= yt_rsc_1_2_q;
  yt_rsc_1_2_radr <= yt_rsc_1_2_i_radr;
  yt_rsc_1_2_d <= yt_rsc_1_2_i_d;
  yt_rsc_1_2_wadr <= yt_rsc_1_2_i_wadr;
  yt_rsc_1_2_i_d_d <= yt_rsc_0_2_i_d_d_iff;
  yt_rsc_1_2_i_q_d <= yt_rsc_1_2_i_q_d_1;
  yt_rsc_1_2_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_1_2_i_wadr_d <= yt_rsc_0_2_i_wadr_d_iff;

  yt_rsc_1_3_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_42_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_1_3_clkr_en,
      clkw_en => yt_rsc_1_3_clkw_en,
      q => yt_rsc_1_3_i_q,
      radr => yt_rsc_1_3_i_radr,
      we => yt_rsc_1_3_we,
      d => yt_rsc_1_3_i_d,
      wadr => yt_rsc_1_3_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_1_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_1_0_i_clkr_en_d,
      d_d => yt_rsc_1_3_i_d_d,
      q_d => yt_rsc_1_3_i_q_d_1,
      radr_d => yt_rsc_1_3_i_radr_d,
      wadr_d => yt_rsc_1_3_i_wadr_d,
      we_d => yt_rsc_1_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_1_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_1_3_i_q <= yt_rsc_1_3_q;
  yt_rsc_1_3_radr <= yt_rsc_1_3_i_radr;
  yt_rsc_1_3_d <= yt_rsc_1_3_i_d;
  yt_rsc_1_3_wadr <= yt_rsc_1_3_i_wadr;
  yt_rsc_1_3_i_d_d <= yt_rsc_0_3_i_d_d_iff;
  yt_rsc_1_3_i_q_d <= yt_rsc_1_3_i_q_d_1;
  yt_rsc_1_3_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_1_3_i_wadr_d <= yt_rsc_0_3_i_wadr_d_iff;

  yt_rsc_1_4_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_43_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_1_4_clkr_en,
      clkw_en => yt_rsc_1_4_clkw_en,
      q => yt_rsc_1_4_i_q,
      radr => yt_rsc_1_4_i_radr,
      we => yt_rsc_1_4_we,
      d => yt_rsc_1_4_i_d,
      wadr => yt_rsc_1_4_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_1_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_1_0_i_clkr_en_d,
      d_d => yt_rsc_1_4_i_d_d,
      q_d => yt_rsc_1_4_i_q_d_1,
      radr_d => yt_rsc_1_4_i_radr_d,
      wadr_d => yt_rsc_1_4_i_wadr_d,
      we_d => yt_rsc_1_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_1_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_1_4_i_q <= yt_rsc_1_4_q;
  yt_rsc_1_4_radr <= yt_rsc_1_4_i_radr;
  yt_rsc_1_4_d <= yt_rsc_1_4_i_d;
  yt_rsc_1_4_wadr <= yt_rsc_1_4_i_wadr;
  yt_rsc_1_4_i_d_d <= yt_rsc_0_4_i_d_d_iff;
  yt_rsc_1_4_i_q_d <= yt_rsc_1_4_i_q_d_1;
  yt_rsc_1_4_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_1_4_i_wadr_d <= yt_rsc_0_4_i_wadr_d_iff;

  yt_rsc_1_5_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_44_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_1_5_clkr_en,
      clkw_en => yt_rsc_1_5_clkw_en,
      q => yt_rsc_1_5_i_q,
      radr => yt_rsc_1_5_i_radr,
      we => yt_rsc_1_5_we,
      d => yt_rsc_1_5_i_d,
      wadr => yt_rsc_1_5_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_1_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_1_0_i_clkr_en_d,
      d_d => yt_rsc_1_5_i_d_d,
      q_d => yt_rsc_1_5_i_q_d_1,
      radr_d => yt_rsc_1_5_i_radr_d,
      wadr_d => yt_rsc_1_5_i_wadr_d,
      we_d => yt_rsc_1_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_1_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_1_5_i_q <= yt_rsc_1_5_q;
  yt_rsc_1_5_radr <= yt_rsc_1_5_i_radr;
  yt_rsc_1_5_d <= yt_rsc_1_5_i_d;
  yt_rsc_1_5_wadr <= yt_rsc_1_5_i_wadr;
  yt_rsc_1_5_i_d_d <= yt_rsc_0_5_i_d_d_iff;
  yt_rsc_1_5_i_q_d <= yt_rsc_1_5_i_q_d_1;
  yt_rsc_1_5_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_1_5_i_wadr_d <= yt_rsc_0_5_i_wadr_d_iff;

  yt_rsc_1_6_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_45_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_1_6_clkr_en,
      clkw_en => yt_rsc_1_6_clkw_en,
      q => yt_rsc_1_6_i_q,
      radr => yt_rsc_1_6_i_radr,
      we => yt_rsc_1_6_we,
      d => yt_rsc_1_6_i_d,
      wadr => yt_rsc_1_6_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_1_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_1_0_i_clkr_en_d,
      d_d => yt_rsc_1_6_i_d_d,
      q_d => yt_rsc_1_6_i_q_d_1,
      radr_d => yt_rsc_1_6_i_radr_d,
      wadr_d => yt_rsc_1_6_i_wadr_d,
      we_d => yt_rsc_1_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_1_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_1_6_i_q <= yt_rsc_1_6_q;
  yt_rsc_1_6_radr <= yt_rsc_1_6_i_radr;
  yt_rsc_1_6_d <= yt_rsc_1_6_i_d;
  yt_rsc_1_6_wadr <= yt_rsc_1_6_i_wadr;
  yt_rsc_1_6_i_d_d <= yt_rsc_0_6_i_d_d_iff;
  yt_rsc_1_6_i_q_d <= yt_rsc_1_6_i_q_d_1;
  yt_rsc_1_6_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_1_6_i_wadr_d <= yt_rsc_0_6_i_wadr_d_iff;

  yt_rsc_1_7_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_46_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_1_7_clkr_en,
      clkw_en => yt_rsc_1_7_clkw_en,
      q => yt_rsc_1_7_i_q,
      radr => yt_rsc_1_7_i_radr,
      we => yt_rsc_1_7_we,
      d => yt_rsc_1_7_i_d,
      wadr => yt_rsc_1_7_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_1_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_1_0_i_clkr_en_d,
      d_d => yt_rsc_1_7_i_d_d,
      q_d => yt_rsc_1_7_i_q_d_1,
      radr_d => yt_rsc_1_7_i_radr_d,
      wadr_d => yt_rsc_1_7_i_wadr_d,
      we_d => yt_rsc_1_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_1_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_1_7_i_q <= yt_rsc_1_7_q;
  yt_rsc_1_7_radr <= yt_rsc_1_7_i_radr;
  yt_rsc_1_7_d <= yt_rsc_1_7_i_d;
  yt_rsc_1_7_wadr <= yt_rsc_1_7_i_wadr;
  yt_rsc_1_7_i_d_d <= yt_rsc_0_7_i_d_d_iff;
  yt_rsc_1_7_i_q_d <= yt_rsc_1_7_i_q_d_1;
  yt_rsc_1_7_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_1_7_i_wadr_d <= yt_rsc_0_0_i_wadr_d_iff;

  yt_rsc_1_8_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_47_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_1_8_clkr_en,
      clkw_en => yt_rsc_1_8_clkw_en,
      q => yt_rsc_1_8_i_q,
      radr => yt_rsc_1_8_i_radr,
      we => yt_rsc_1_8_we,
      d => yt_rsc_1_8_i_d,
      wadr => yt_rsc_1_8_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_1_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_1_0_i_clkr_en_d,
      d_d => yt_rsc_1_8_i_d_d,
      q_d => yt_rsc_1_8_i_q_d_1,
      radr_d => yt_rsc_1_8_i_radr_d,
      wadr_d => yt_rsc_1_8_i_wadr_d,
      we_d => yt_rsc_1_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_1_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_1_8_i_q <= yt_rsc_1_8_q;
  yt_rsc_1_8_radr <= yt_rsc_1_8_i_radr;
  yt_rsc_1_8_d <= yt_rsc_1_8_i_d;
  yt_rsc_1_8_wadr <= yt_rsc_1_8_i_wadr;
  yt_rsc_1_8_i_d_d <= yt_rsc_0_8_i_d_d_iff;
  yt_rsc_1_8_i_q_d <= yt_rsc_1_8_i_q_d_1;
  yt_rsc_1_8_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_1_8_i_wadr_d <= yt_rsc_0_1_i_wadr_d_iff;

  yt_rsc_1_9_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_48_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_1_9_clkr_en,
      clkw_en => yt_rsc_1_9_clkw_en,
      q => yt_rsc_1_9_i_q,
      radr => yt_rsc_1_9_i_radr,
      we => yt_rsc_1_9_we,
      d => yt_rsc_1_9_i_d,
      wadr => yt_rsc_1_9_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_1_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_1_0_i_clkr_en_d,
      d_d => yt_rsc_1_9_i_d_d,
      q_d => yt_rsc_1_9_i_q_d_1,
      radr_d => yt_rsc_1_9_i_radr_d,
      wadr_d => yt_rsc_1_9_i_wadr_d,
      we_d => yt_rsc_1_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_1_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_1_9_i_q <= yt_rsc_1_9_q;
  yt_rsc_1_9_radr <= yt_rsc_1_9_i_radr;
  yt_rsc_1_9_d <= yt_rsc_1_9_i_d;
  yt_rsc_1_9_wadr <= yt_rsc_1_9_i_wadr;
  yt_rsc_1_9_i_d_d <= yt_rsc_0_9_i_d_d_iff;
  yt_rsc_1_9_i_q_d <= yt_rsc_1_9_i_q_d_1;
  yt_rsc_1_9_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_1_9_i_wadr_d <= yt_rsc_0_2_i_wadr_d_iff;

  yt_rsc_1_10_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_49_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_1_10_clkr_en,
      clkw_en => yt_rsc_1_10_clkw_en,
      q => yt_rsc_1_10_i_q,
      radr => yt_rsc_1_10_i_radr,
      we => yt_rsc_1_10_we,
      d => yt_rsc_1_10_i_d,
      wadr => yt_rsc_1_10_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_1_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_1_0_i_clkr_en_d,
      d_d => yt_rsc_1_10_i_d_d,
      q_d => yt_rsc_1_10_i_q_d_1,
      radr_d => yt_rsc_1_10_i_radr_d,
      wadr_d => yt_rsc_1_10_i_wadr_d,
      we_d => yt_rsc_1_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_1_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_1_10_i_q <= yt_rsc_1_10_q;
  yt_rsc_1_10_radr <= yt_rsc_1_10_i_radr;
  yt_rsc_1_10_d <= yt_rsc_1_10_i_d;
  yt_rsc_1_10_wadr <= yt_rsc_1_10_i_wadr;
  yt_rsc_1_10_i_d_d <= yt_rsc_0_10_i_d_d_iff;
  yt_rsc_1_10_i_q_d <= yt_rsc_1_10_i_q_d_1;
  yt_rsc_1_10_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_1_10_i_wadr_d <= yt_rsc_0_10_i_wadr_d_iff;

  yt_rsc_1_11_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_50_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_1_11_clkr_en,
      clkw_en => yt_rsc_1_11_clkw_en,
      q => yt_rsc_1_11_i_q,
      radr => yt_rsc_1_11_i_radr,
      we => yt_rsc_1_11_we,
      d => yt_rsc_1_11_i_d,
      wadr => yt_rsc_1_11_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_1_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_1_0_i_clkr_en_d,
      d_d => yt_rsc_1_11_i_d_d,
      q_d => yt_rsc_1_11_i_q_d_1,
      radr_d => yt_rsc_1_11_i_radr_d,
      wadr_d => yt_rsc_1_11_i_wadr_d,
      we_d => yt_rsc_1_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_1_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_1_11_i_q <= yt_rsc_1_11_q;
  yt_rsc_1_11_radr <= yt_rsc_1_11_i_radr;
  yt_rsc_1_11_d <= yt_rsc_1_11_i_d;
  yt_rsc_1_11_wadr <= yt_rsc_1_11_i_wadr;
  yt_rsc_1_11_i_d_d <= yt_rsc_0_11_i_d_d_iff;
  yt_rsc_1_11_i_q_d <= yt_rsc_1_11_i_q_d_1;
  yt_rsc_1_11_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_1_11_i_wadr_d <= yt_rsc_0_11_i_wadr_d_iff;

  yt_rsc_1_12_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_51_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_1_12_clkr_en,
      clkw_en => yt_rsc_1_12_clkw_en,
      q => yt_rsc_1_12_i_q,
      radr => yt_rsc_1_12_i_radr,
      we => yt_rsc_1_12_we,
      d => yt_rsc_1_12_i_d,
      wadr => yt_rsc_1_12_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_1_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_1_0_i_clkr_en_d,
      d_d => yt_rsc_1_12_i_d_d,
      q_d => yt_rsc_1_12_i_q_d_1,
      radr_d => yt_rsc_1_12_i_radr_d,
      wadr_d => yt_rsc_1_12_i_wadr_d,
      we_d => yt_rsc_1_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_1_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_1_12_i_q <= yt_rsc_1_12_q;
  yt_rsc_1_12_radr <= yt_rsc_1_12_i_radr;
  yt_rsc_1_12_d <= yt_rsc_1_12_i_d;
  yt_rsc_1_12_wadr <= yt_rsc_1_12_i_wadr;
  yt_rsc_1_12_i_d_d <= yt_rsc_0_12_i_d_d_iff;
  yt_rsc_1_12_i_q_d <= yt_rsc_1_12_i_q_d_1;
  yt_rsc_1_12_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_1_12_i_wadr_d <= yt_rsc_0_3_i_wadr_d_iff;

  yt_rsc_1_13_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_52_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_1_13_clkr_en,
      clkw_en => yt_rsc_1_13_clkw_en,
      q => yt_rsc_1_13_i_q,
      radr => yt_rsc_1_13_i_radr,
      we => yt_rsc_1_13_we,
      d => yt_rsc_1_13_i_d,
      wadr => yt_rsc_1_13_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_1_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_1_0_i_clkr_en_d,
      d_d => yt_rsc_1_13_i_d_d,
      q_d => yt_rsc_1_13_i_q_d_1,
      radr_d => yt_rsc_1_13_i_radr_d,
      wadr_d => yt_rsc_1_13_i_wadr_d,
      we_d => yt_rsc_1_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_1_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_1_13_i_q <= yt_rsc_1_13_q;
  yt_rsc_1_13_radr <= yt_rsc_1_13_i_radr;
  yt_rsc_1_13_d <= yt_rsc_1_13_i_d;
  yt_rsc_1_13_wadr <= yt_rsc_1_13_i_wadr;
  yt_rsc_1_13_i_d_d <= yt_rsc_0_13_i_d_d_iff;
  yt_rsc_1_13_i_q_d <= yt_rsc_1_13_i_q_d_1;
  yt_rsc_1_13_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_1_13_i_wadr_d <= yt_rsc_0_4_i_wadr_d_iff;

  yt_rsc_1_14_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_53_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_1_14_clkr_en,
      clkw_en => yt_rsc_1_14_clkw_en,
      q => yt_rsc_1_14_i_q,
      radr => yt_rsc_1_14_i_radr,
      we => yt_rsc_1_14_we,
      d => yt_rsc_1_14_i_d,
      wadr => yt_rsc_1_14_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_1_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_1_0_i_clkr_en_d,
      d_d => yt_rsc_1_14_i_d_d,
      q_d => yt_rsc_1_14_i_q_d_1,
      radr_d => yt_rsc_1_14_i_radr_d,
      wadr_d => yt_rsc_1_14_i_wadr_d,
      we_d => yt_rsc_1_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_1_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_1_14_i_q <= yt_rsc_1_14_q;
  yt_rsc_1_14_radr <= yt_rsc_1_14_i_radr;
  yt_rsc_1_14_d <= yt_rsc_1_14_i_d;
  yt_rsc_1_14_wadr <= yt_rsc_1_14_i_wadr;
  yt_rsc_1_14_i_d_d <= yt_rsc_0_14_i_d_d_iff;
  yt_rsc_1_14_i_q_d <= yt_rsc_1_14_i_q_d_1;
  yt_rsc_1_14_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_1_14_i_wadr_d <= yt_rsc_0_5_i_wadr_d_iff;

  yt_rsc_1_15_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_54_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_1_15_clkr_en,
      clkw_en => yt_rsc_1_15_clkw_en,
      q => yt_rsc_1_15_i_q,
      radr => yt_rsc_1_15_i_radr,
      we => yt_rsc_1_15_we,
      d => yt_rsc_1_15_i_d,
      wadr => yt_rsc_1_15_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_1_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_1_0_i_clkr_en_d,
      d_d => yt_rsc_1_15_i_d_d,
      q_d => yt_rsc_1_15_i_q_d_1,
      radr_d => yt_rsc_1_15_i_radr_d,
      wadr_d => yt_rsc_1_15_i_wadr_d,
      we_d => yt_rsc_1_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_1_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_1_15_i_q <= yt_rsc_1_15_q;
  yt_rsc_1_15_radr <= yt_rsc_1_15_i_radr;
  yt_rsc_1_15_d <= yt_rsc_1_15_i_d;
  yt_rsc_1_15_wadr <= yt_rsc_1_15_i_wadr;
  yt_rsc_1_15_i_d_d <= yt_rsc_0_15_i_d_d_iff;
  yt_rsc_1_15_i_q_d <= yt_rsc_1_15_i_q_d_1;
  yt_rsc_1_15_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_1_15_i_wadr_d <= yt_rsc_0_6_i_wadr_d_iff;

  yt_rsc_1_16_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_55_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_1_16_clkr_en,
      clkw_en => yt_rsc_1_16_clkw_en,
      q => yt_rsc_1_16_i_q,
      radr => yt_rsc_1_16_i_radr,
      we => yt_rsc_1_16_we,
      d => yt_rsc_1_16_i_d,
      wadr => yt_rsc_1_16_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_1_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_1_16_i_clkr_en_d,
      d_d => yt_rsc_1_16_i_d_d,
      q_d => yt_rsc_1_16_i_q_d_1,
      radr_d => yt_rsc_1_16_i_radr_d,
      wadr_d => yt_rsc_1_16_i_wadr_d,
      we_d => yt_rsc_1_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_1_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_1_16_i_q <= yt_rsc_1_16_q;
  yt_rsc_1_16_radr <= yt_rsc_1_16_i_radr;
  yt_rsc_1_16_d <= yt_rsc_1_16_i_d;
  yt_rsc_1_16_wadr <= yt_rsc_1_16_i_wadr;
  yt_rsc_1_16_i_d_d <= yt_rsc_0_0_i_d_d_iff;
  yt_rsc_1_16_i_q_d <= yt_rsc_1_16_i_q_d_1;
  yt_rsc_1_16_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_1_16_i_wadr_d <= yt_rsc_0_0_i_wadr_d_iff;

  yt_rsc_1_17_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_56_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_1_17_clkr_en,
      clkw_en => yt_rsc_1_17_clkw_en,
      q => yt_rsc_1_17_i_q,
      radr => yt_rsc_1_17_i_radr,
      we => yt_rsc_1_17_we,
      d => yt_rsc_1_17_i_d,
      wadr => yt_rsc_1_17_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_1_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_1_16_i_clkr_en_d,
      d_d => yt_rsc_1_17_i_d_d,
      q_d => yt_rsc_1_17_i_q_d_1,
      radr_d => yt_rsc_1_17_i_radr_d,
      wadr_d => yt_rsc_1_17_i_wadr_d,
      we_d => yt_rsc_1_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_1_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_1_17_i_q <= yt_rsc_1_17_q;
  yt_rsc_1_17_radr <= yt_rsc_1_17_i_radr;
  yt_rsc_1_17_d <= yt_rsc_1_17_i_d;
  yt_rsc_1_17_wadr <= yt_rsc_1_17_i_wadr;
  yt_rsc_1_17_i_d_d <= yt_rsc_0_1_i_d_d_iff;
  yt_rsc_1_17_i_q_d <= yt_rsc_1_17_i_q_d_1;
  yt_rsc_1_17_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_1_17_i_wadr_d <= yt_rsc_0_1_i_wadr_d_iff;

  yt_rsc_1_18_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_57_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_1_18_clkr_en,
      clkw_en => yt_rsc_1_18_clkw_en,
      q => yt_rsc_1_18_i_q,
      radr => yt_rsc_1_18_i_radr,
      we => yt_rsc_1_18_we,
      d => yt_rsc_1_18_i_d,
      wadr => yt_rsc_1_18_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_1_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_1_16_i_clkr_en_d,
      d_d => yt_rsc_1_18_i_d_d,
      q_d => yt_rsc_1_18_i_q_d_1,
      radr_d => yt_rsc_1_18_i_radr_d,
      wadr_d => yt_rsc_1_18_i_wadr_d,
      we_d => yt_rsc_1_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_1_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_1_18_i_q <= yt_rsc_1_18_q;
  yt_rsc_1_18_radr <= yt_rsc_1_18_i_radr;
  yt_rsc_1_18_d <= yt_rsc_1_18_i_d;
  yt_rsc_1_18_wadr <= yt_rsc_1_18_i_wadr;
  yt_rsc_1_18_i_d_d <= yt_rsc_0_2_i_d_d_iff;
  yt_rsc_1_18_i_q_d <= yt_rsc_1_18_i_q_d_1;
  yt_rsc_1_18_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_1_18_i_wadr_d <= yt_rsc_0_2_i_wadr_d_iff;

  yt_rsc_1_19_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_58_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_1_19_clkr_en,
      clkw_en => yt_rsc_1_19_clkw_en,
      q => yt_rsc_1_19_i_q,
      radr => yt_rsc_1_19_i_radr,
      we => yt_rsc_1_19_we,
      d => yt_rsc_1_19_i_d,
      wadr => yt_rsc_1_19_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_1_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_1_16_i_clkr_en_d,
      d_d => yt_rsc_1_19_i_d_d,
      q_d => yt_rsc_1_19_i_q_d_1,
      radr_d => yt_rsc_1_19_i_radr_d,
      wadr_d => yt_rsc_1_19_i_wadr_d,
      we_d => yt_rsc_1_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_1_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_1_19_i_q <= yt_rsc_1_19_q;
  yt_rsc_1_19_radr <= yt_rsc_1_19_i_radr;
  yt_rsc_1_19_d <= yt_rsc_1_19_i_d;
  yt_rsc_1_19_wadr <= yt_rsc_1_19_i_wadr;
  yt_rsc_1_19_i_d_d <= yt_rsc_0_3_i_d_d_iff;
  yt_rsc_1_19_i_q_d <= yt_rsc_1_19_i_q_d_1;
  yt_rsc_1_19_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_1_19_i_wadr_d <= yt_rsc_0_3_i_wadr_d_iff;

  yt_rsc_1_20_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_59_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_1_20_clkr_en,
      clkw_en => yt_rsc_1_20_clkw_en,
      q => yt_rsc_1_20_i_q,
      radr => yt_rsc_1_20_i_radr,
      we => yt_rsc_1_20_we,
      d => yt_rsc_1_20_i_d,
      wadr => yt_rsc_1_20_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_1_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_1_16_i_clkr_en_d,
      d_d => yt_rsc_1_20_i_d_d,
      q_d => yt_rsc_1_20_i_q_d_1,
      radr_d => yt_rsc_1_20_i_radr_d,
      wadr_d => yt_rsc_1_20_i_wadr_d,
      we_d => yt_rsc_1_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_1_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_1_20_i_q <= yt_rsc_1_20_q;
  yt_rsc_1_20_radr <= yt_rsc_1_20_i_radr;
  yt_rsc_1_20_d <= yt_rsc_1_20_i_d;
  yt_rsc_1_20_wadr <= yt_rsc_1_20_i_wadr;
  yt_rsc_1_20_i_d_d <= yt_rsc_0_4_i_d_d_iff;
  yt_rsc_1_20_i_q_d <= yt_rsc_1_20_i_q_d_1;
  yt_rsc_1_20_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_1_20_i_wadr_d <= yt_rsc_0_4_i_wadr_d_iff;

  yt_rsc_1_21_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_60_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_1_21_clkr_en,
      clkw_en => yt_rsc_1_21_clkw_en,
      q => yt_rsc_1_21_i_q,
      radr => yt_rsc_1_21_i_radr,
      we => yt_rsc_1_21_we,
      d => yt_rsc_1_21_i_d,
      wadr => yt_rsc_1_21_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_1_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_1_16_i_clkr_en_d,
      d_d => yt_rsc_1_21_i_d_d,
      q_d => yt_rsc_1_21_i_q_d_1,
      radr_d => yt_rsc_1_21_i_radr_d,
      wadr_d => yt_rsc_1_21_i_wadr_d,
      we_d => yt_rsc_1_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_1_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_1_21_i_q <= yt_rsc_1_21_q;
  yt_rsc_1_21_radr <= yt_rsc_1_21_i_radr;
  yt_rsc_1_21_d <= yt_rsc_1_21_i_d;
  yt_rsc_1_21_wadr <= yt_rsc_1_21_i_wadr;
  yt_rsc_1_21_i_d_d <= yt_rsc_0_5_i_d_d_iff;
  yt_rsc_1_21_i_q_d <= yt_rsc_1_21_i_q_d_1;
  yt_rsc_1_21_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_1_21_i_wadr_d <= yt_rsc_0_5_i_wadr_d_iff;

  yt_rsc_1_22_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_61_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_1_22_clkr_en,
      clkw_en => yt_rsc_1_22_clkw_en,
      q => yt_rsc_1_22_i_q,
      radr => yt_rsc_1_22_i_radr,
      we => yt_rsc_1_22_we,
      d => yt_rsc_1_22_i_d,
      wadr => yt_rsc_1_22_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_1_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_1_16_i_clkr_en_d,
      d_d => yt_rsc_1_22_i_d_d,
      q_d => yt_rsc_1_22_i_q_d_1,
      radr_d => yt_rsc_1_22_i_radr_d,
      wadr_d => yt_rsc_1_22_i_wadr_d,
      we_d => yt_rsc_1_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_1_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_1_22_i_q <= yt_rsc_1_22_q;
  yt_rsc_1_22_radr <= yt_rsc_1_22_i_radr;
  yt_rsc_1_22_d <= yt_rsc_1_22_i_d;
  yt_rsc_1_22_wadr <= yt_rsc_1_22_i_wadr;
  yt_rsc_1_22_i_d_d <= yt_rsc_0_6_i_d_d_iff;
  yt_rsc_1_22_i_q_d <= yt_rsc_1_22_i_q_d_1;
  yt_rsc_1_22_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_1_22_i_wadr_d <= yt_rsc_0_6_i_wadr_d_iff;

  yt_rsc_1_23_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_62_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_1_23_clkr_en,
      clkw_en => yt_rsc_1_23_clkw_en,
      q => yt_rsc_1_23_i_q,
      radr => yt_rsc_1_23_i_radr,
      we => yt_rsc_1_23_we,
      d => yt_rsc_1_23_i_d,
      wadr => yt_rsc_1_23_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_1_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_1_16_i_clkr_en_d,
      d_d => yt_rsc_1_23_i_d_d,
      q_d => yt_rsc_1_23_i_q_d_1,
      radr_d => yt_rsc_1_23_i_radr_d,
      wadr_d => yt_rsc_1_23_i_wadr_d,
      we_d => yt_rsc_1_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_1_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_1_23_i_q <= yt_rsc_1_23_q;
  yt_rsc_1_23_radr <= yt_rsc_1_23_i_radr;
  yt_rsc_1_23_d <= yt_rsc_1_23_i_d;
  yt_rsc_1_23_wadr <= yt_rsc_1_23_i_wadr;
  yt_rsc_1_23_i_d_d <= yt_rsc_0_7_i_d_d_iff;
  yt_rsc_1_23_i_q_d <= yt_rsc_1_23_i_q_d_1;
  yt_rsc_1_23_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_1_23_i_wadr_d <= yt_rsc_0_0_i_wadr_d_iff;

  yt_rsc_1_24_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_63_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_1_24_clkr_en,
      clkw_en => yt_rsc_1_24_clkw_en,
      q => yt_rsc_1_24_i_q,
      radr => yt_rsc_1_24_i_radr,
      we => yt_rsc_1_24_we,
      d => yt_rsc_1_24_i_d,
      wadr => yt_rsc_1_24_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_1_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_1_16_i_clkr_en_d,
      d_d => yt_rsc_1_24_i_d_d,
      q_d => yt_rsc_1_24_i_q_d_1,
      radr_d => yt_rsc_1_24_i_radr_d,
      wadr_d => yt_rsc_1_24_i_wadr_d,
      we_d => yt_rsc_1_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_1_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_1_24_i_q <= yt_rsc_1_24_q;
  yt_rsc_1_24_radr <= yt_rsc_1_24_i_radr;
  yt_rsc_1_24_d <= yt_rsc_1_24_i_d;
  yt_rsc_1_24_wadr <= yt_rsc_1_24_i_wadr;
  yt_rsc_1_24_i_d_d <= yt_rsc_0_8_i_d_d_iff;
  yt_rsc_1_24_i_q_d <= yt_rsc_1_24_i_q_d_1;
  yt_rsc_1_24_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_1_24_i_wadr_d <= yt_rsc_0_1_i_wadr_d_iff;

  yt_rsc_1_25_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_64_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_1_25_clkr_en,
      clkw_en => yt_rsc_1_25_clkw_en,
      q => yt_rsc_1_25_i_q,
      radr => yt_rsc_1_25_i_radr,
      we => yt_rsc_1_25_we,
      d => yt_rsc_1_25_i_d,
      wadr => yt_rsc_1_25_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_1_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_1_16_i_clkr_en_d,
      d_d => yt_rsc_1_25_i_d_d,
      q_d => yt_rsc_1_25_i_q_d_1,
      radr_d => yt_rsc_1_25_i_radr_d,
      wadr_d => yt_rsc_1_25_i_wadr_d,
      we_d => yt_rsc_1_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_1_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_1_25_i_q <= yt_rsc_1_25_q;
  yt_rsc_1_25_radr <= yt_rsc_1_25_i_radr;
  yt_rsc_1_25_d <= yt_rsc_1_25_i_d;
  yt_rsc_1_25_wadr <= yt_rsc_1_25_i_wadr;
  yt_rsc_1_25_i_d_d <= yt_rsc_0_9_i_d_d_iff;
  yt_rsc_1_25_i_q_d <= yt_rsc_1_25_i_q_d_1;
  yt_rsc_1_25_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_1_25_i_wadr_d <= yt_rsc_0_2_i_wadr_d_iff;

  yt_rsc_1_26_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_65_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_1_26_clkr_en,
      clkw_en => yt_rsc_1_26_clkw_en,
      q => yt_rsc_1_26_i_q,
      radr => yt_rsc_1_26_i_radr,
      we => yt_rsc_1_26_we,
      d => yt_rsc_1_26_i_d,
      wadr => yt_rsc_1_26_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_1_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_1_16_i_clkr_en_d,
      d_d => yt_rsc_1_26_i_d_d,
      q_d => yt_rsc_1_26_i_q_d_1,
      radr_d => yt_rsc_1_26_i_radr_d,
      wadr_d => yt_rsc_1_26_i_wadr_d,
      we_d => yt_rsc_1_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_1_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_1_26_i_q <= yt_rsc_1_26_q;
  yt_rsc_1_26_radr <= yt_rsc_1_26_i_radr;
  yt_rsc_1_26_d <= yt_rsc_1_26_i_d;
  yt_rsc_1_26_wadr <= yt_rsc_1_26_i_wadr;
  yt_rsc_1_26_i_d_d <= yt_rsc_0_10_i_d_d_iff;
  yt_rsc_1_26_i_q_d <= yt_rsc_1_26_i_q_d_1;
  yt_rsc_1_26_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_1_26_i_wadr_d <= yt_rsc_0_10_i_wadr_d_iff;

  yt_rsc_1_27_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_66_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_1_27_clkr_en,
      clkw_en => yt_rsc_1_27_clkw_en,
      q => yt_rsc_1_27_i_q,
      radr => yt_rsc_1_27_i_radr,
      we => yt_rsc_1_27_we,
      d => yt_rsc_1_27_i_d,
      wadr => yt_rsc_1_27_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_1_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_1_16_i_clkr_en_d,
      d_d => yt_rsc_1_27_i_d_d,
      q_d => yt_rsc_1_27_i_q_d_1,
      radr_d => yt_rsc_1_27_i_radr_d,
      wadr_d => yt_rsc_1_27_i_wadr_d,
      we_d => yt_rsc_1_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_1_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_1_27_i_q <= yt_rsc_1_27_q;
  yt_rsc_1_27_radr <= yt_rsc_1_27_i_radr;
  yt_rsc_1_27_d <= yt_rsc_1_27_i_d;
  yt_rsc_1_27_wadr <= yt_rsc_1_27_i_wadr;
  yt_rsc_1_27_i_d_d <= yt_rsc_0_11_i_d_d_iff;
  yt_rsc_1_27_i_q_d <= yt_rsc_1_27_i_q_d_1;
  yt_rsc_1_27_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_1_27_i_wadr_d <= yt_rsc_0_11_i_wadr_d_iff;

  yt_rsc_1_28_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_67_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_1_28_clkr_en,
      clkw_en => yt_rsc_1_28_clkw_en,
      q => yt_rsc_1_28_i_q,
      radr => yt_rsc_1_28_i_radr,
      we => yt_rsc_1_28_we,
      d => yt_rsc_1_28_i_d,
      wadr => yt_rsc_1_28_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_1_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_1_16_i_clkr_en_d,
      d_d => yt_rsc_1_28_i_d_d,
      q_d => yt_rsc_1_28_i_q_d_1,
      radr_d => yt_rsc_1_28_i_radr_d,
      wadr_d => yt_rsc_1_28_i_wadr_d,
      we_d => yt_rsc_1_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_1_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_1_28_i_q <= yt_rsc_1_28_q;
  yt_rsc_1_28_radr <= yt_rsc_1_28_i_radr;
  yt_rsc_1_28_d <= yt_rsc_1_28_i_d;
  yt_rsc_1_28_wadr <= yt_rsc_1_28_i_wadr;
  yt_rsc_1_28_i_d_d <= yt_rsc_0_12_i_d_d_iff;
  yt_rsc_1_28_i_q_d <= yt_rsc_1_28_i_q_d_1;
  yt_rsc_1_28_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_1_28_i_wadr_d <= yt_rsc_0_3_i_wadr_d_iff;

  yt_rsc_1_29_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_68_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_1_29_clkr_en,
      clkw_en => yt_rsc_1_29_clkw_en,
      q => yt_rsc_1_29_i_q,
      radr => yt_rsc_1_29_i_radr,
      we => yt_rsc_1_29_we,
      d => yt_rsc_1_29_i_d,
      wadr => yt_rsc_1_29_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_1_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_1_16_i_clkr_en_d,
      d_d => yt_rsc_1_29_i_d_d,
      q_d => yt_rsc_1_29_i_q_d_1,
      radr_d => yt_rsc_1_29_i_radr_d,
      wadr_d => yt_rsc_1_29_i_wadr_d,
      we_d => yt_rsc_1_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_1_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_1_29_i_q <= yt_rsc_1_29_q;
  yt_rsc_1_29_radr <= yt_rsc_1_29_i_radr;
  yt_rsc_1_29_d <= yt_rsc_1_29_i_d;
  yt_rsc_1_29_wadr <= yt_rsc_1_29_i_wadr;
  yt_rsc_1_29_i_d_d <= yt_rsc_0_13_i_d_d_iff;
  yt_rsc_1_29_i_q_d <= yt_rsc_1_29_i_q_d_1;
  yt_rsc_1_29_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_1_29_i_wadr_d <= yt_rsc_0_4_i_wadr_d_iff;

  yt_rsc_1_30_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_69_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_1_30_clkr_en,
      clkw_en => yt_rsc_1_30_clkw_en,
      q => yt_rsc_1_30_i_q,
      radr => yt_rsc_1_30_i_radr,
      we => yt_rsc_1_30_we,
      d => yt_rsc_1_30_i_d,
      wadr => yt_rsc_1_30_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_1_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_1_16_i_clkr_en_d,
      d_d => yt_rsc_1_30_i_d_d,
      q_d => yt_rsc_1_30_i_q_d_1,
      radr_d => yt_rsc_1_30_i_radr_d,
      wadr_d => yt_rsc_1_30_i_wadr_d,
      we_d => yt_rsc_1_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_1_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_1_30_i_q <= yt_rsc_1_30_q;
  yt_rsc_1_30_radr <= yt_rsc_1_30_i_radr;
  yt_rsc_1_30_d <= yt_rsc_1_30_i_d;
  yt_rsc_1_30_wadr <= yt_rsc_1_30_i_wadr;
  yt_rsc_1_30_i_d_d <= yt_rsc_0_14_i_d_d_iff;
  yt_rsc_1_30_i_q_d <= yt_rsc_1_30_i_q_d_1;
  yt_rsc_1_30_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_1_30_i_wadr_d <= yt_rsc_0_5_i_wadr_d_iff;

  yt_rsc_1_31_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_70_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_1_31_clkr_en,
      clkw_en => yt_rsc_1_31_clkw_en,
      q => yt_rsc_1_31_i_q,
      radr => yt_rsc_1_31_i_radr,
      we => yt_rsc_1_31_we,
      d => yt_rsc_1_31_i_d,
      wadr => yt_rsc_1_31_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_1_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_1_16_i_clkr_en_d,
      d_d => yt_rsc_1_31_i_d_d,
      q_d => yt_rsc_1_31_i_q_d_1,
      radr_d => yt_rsc_1_31_i_radr_d,
      wadr_d => yt_rsc_1_31_i_wadr_d,
      we_d => yt_rsc_1_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_1_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_1_31_i_q <= yt_rsc_1_31_q;
  yt_rsc_1_31_radr <= yt_rsc_1_31_i_radr;
  yt_rsc_1_31_d <= yt_rsc_1_31_i_d;
  yt_rsc_1_31_wadr <= yt_rsc_1_31_i_wadr;
  yt_rsc_1_31_i_d_d <= yt_rsc_0_15_i_d_d_iff;
  yt_rsc_1_31_i_q_d <= yt_rsc_1_31_i_q_d_1;
  yt_rsc_1_31_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_1_31_i_wadr_d <= yt_rsc_0_6_i_wadr_d_iff;

  yt_rsc_2_0_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_71_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_2_0_clkr_en,
      clkw_en => yt_rsc_2_0_clkw_en,
      q => yt_rsc_2_0_i_q,
      radr => yt_rsc_2_0_i_radr,
      we => yt_rsc_2_0_we,
      d => yt_rsc_2_0_i_d,
      wadr => yt_rsc_2_0_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_2_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_2_0_i_clkr_en_d,
      d_d => yt_rsc_2_0_i_d_d,
      q_d => yt_rsc_2_0_i_q_d_1,
      radr_d => yt_rsc_2_0_i_radr_d,
      wadr_d => yt_rsc_2_0_i_wadr_d,
      we_d => yt_rsc_2_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_2_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_2_0_i_q <= yt_rsc_2_0_q;
  yt_rsc_2_0_radr <= yt_rsc_2_0_i_radr;
  yt_rsc_2_0_d <= yt_rsc_2_0_i_d;
  yt_rsc_2_0_wadr <= yt_rsc_2_0_i_wadr;
  yt_rsc_2_0_i_d_d <= yt_rsc_0_0_i_d_d_iff;
  yt_rsc_2_0_i_q_d <= yt_rsc_2_0_i_q_d_1;
  yt_rsc_2_0_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_2_0_i_wadr_d <= yt_rsc_0_0_i_wadr_d_iff;

  yt_rsc_2_1_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_72_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_2_1_clkr_en,
      clkw_en => yt_rsc_2_1_clkw_en,
      q => yt_rsc_2_1_i_q,
      radr => yt_rsc_2_1_i_radr,
      we => yt_rsc_2_1_we,
      d => yt_rsc_2_1_i_d,
      wadr => yt_rsc_2_1_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_2_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_2_0_i_clkr_en_d,
      d_d => yt_rsc_2_1_i_d_d,
      q_d => yt_rsc_2_1_i_q_d_1,
      radr_d => yt_rsc_2_1_i_radr_d,
      wadr_d => yt_rsc_2_1_i_wadr_d,
      we_d => yt_rsc_2_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_2_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_2_1_i_q <= yt_rsc_2_1_q;
  yt_rsc_2_1_radr <= yt_rsc_2_1_i_radr;
  yt_rsc_2_1_d <= yt_rsc_2_1_i_d;
  yt_rsc_2_1_wadr <= yt_rsc_2_1_i_wadr;
  yt_rsc_2_1_i_d_d <= yt_rsc_0_1_i_d_d_iff;
  yt_rsc_2_1_i_q_d <= yt_rsc_2_1_i_q_d_1;
  yt_rsc_2_1_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_2_1_i_wadr_d <= yt_rsc_0_1_i_wadr_d_iff;

  yt_rsc_2_2_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_73_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_2_2_clkr_en,
      clkw_en => yt_rsc_2_2_clkw_en,
      q => yt_rsc_2_2_i_q,
      radr => yt_rsc_2_2_i_radr,
      we => yt_rsc_2_2_we,
      d => yt_rsc_2_2_i_d,
      wadr => yt_rsc_2_2_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_2_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_2_0_i_clkr_en_d,
      d_d => yt_rsc_2_2_i_d_d,
      q_d => yt_rsc_2_2_i_q_d_1,
      radr_d => yt_rsc_2_2_i_radr_d,
      wadr_d => yt_rsc_2_2_i_wadr_d,
      we_d => yt_rsc_2_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_2_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_2_2_i_q <= yt_rsc_2_2_q;
  yt_rsc_2_2_radr <= yt_rsc_2_2_i_radr;
  yt_rsc_2_2_d <= yt_rsc_2_2_i_d;
  yt_rsc_2_2_wadr <= yt_rsc_2_2_i_wadr;
  yt_rsc_2_2_i_d_d <= yt_rsc_0_2_i_d_d_iff;
  yt_rsc_2_2_i_q_d <= yt_rsc_2_2_i_q_d_1;
  yt_rsc_2_2_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_2_2_i_wadr_d <= yt_rsc_0_2_i_wadr_d_iff;

  yt_rsc_2_3_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_74_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_2_3_clkr_en,
      clkw_en => yt_rsc_2_3_clkw_en,
      q => yt_rsc_2_3_i_q,
      radr => yt_rsc_2_3_i_radr,
      we => yt_rsc_2_3_we,
      d => yt_rsc_2_3_i_d,
      wadr => yt_rsc_2_3_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_2_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_2_0_i_clkr_en_d,
      d_d => yt_rsc_2_3_i_d_d,
      q_d => yt_rsc_2_3_i_q_d_1,
      radr_d => yt_rsc_2_3_i_radr_d,
      wadr_d => yt_rsc_2_3_i_wadr_d,
      we_d => yt_rsc_2_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_2_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_2_3_i_q <= yt_rsc_2_3_q;
  yt_rsc_2_3_radr <= yt_rsc_2_3_i_radr;
  yt_rsc_2_3_d <= yt_rsc_2_3_i_d;
  yt_rsc_2_3_wadr <= yt_rsc_2_3_i_wadr;
  yt_rsc_2_3_i_d_d <= yt_rsc_0_3_i_d_d_iff;
  yt_rsc_2_3_i_q_d <= yt_rsc_2_3_i_q_d_1;
  yt_rsc_2_3_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_2_3_i_wadr_d <= yt_rsc_0_3_i_wadr_d_iff;

  yt_rsc_2_4_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_75_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_2_4_clkr_en,
      clkw_en => yt_rsc_2_4_clkw_en,
      q => yt_rsc_2_4_i_q,
      radr => yt_rsc_2_4_i_radr,
      we => yt_rsc_2_4_we,
      d => yt_rsc_2_4_i_d,
      wadr => yt_rsc_2_4_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_2_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_2_0_i_clkr_en_d,
      d_d => yt_rsc_2_4_i_d_d,
      q_d => yt_rsc_2_4_i_q_d_1,
      radr_d => yt_rsc_2_4_i_radr_d,
      wadr_d => yt_rsc_2_4_i_wadr_d,
      we_d => yt_rsc_2_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_2_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_2_4_i_q <= yt_rsc_2_4_q;
  yt_rsc_2_4_radr <= yt_rsc_2_4_i_radr;
  yt_rsc_2_4_d <= yt_rsc_2_4_i_d;
  yt_rsc_2_4_wadr <= yt_rsc_2_4_i_wadr;
  yt_rsc_2_4_i_d_d <= yt_rsc_0_4_i_d_d_iff;
  yt_rsc_2_4_i_q_d <= yt_rsc_2_4_i_q_d_1;
  yt_rsc_2_4_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_2_4_i_wadr_d <= yt_rsc_0_4_i_wadr_d_iff;

  yt_rsc_2_5_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_76_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_2_5_clkr_en,
      clkw_en => yt_rsc_2_5_clkw_en,
      q => yt_rsc_2_5_i_q,
      radr => yt_rsc_2_5_i_radr,
      we => yt_rsc_2_5_we,
      d => yt_rsc_2_5_i_d,
      wadr => yt_rsc_2_5_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_2_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_2_0_i_clkr_en_d,
      d_d => yt_rsc_2_5_i_d_d,
      q_d => yt_rsc_2_5_i_q_d_1,
      radr_d => yt_rsc_2_5_i_radr_d,
      wadr_d => yt_rsc_2_5_i_wadr_d,
      we_d => yt_rsc_2_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_2_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_2_5_i_q <= yt_rsc_2_5_q;
  yt_rsc_2_5_radr <= yt_rsc_2_5_i_radr;
  yt_rsc_2_5_d <= yt_rsc_2_5_i_d;
  yt_rsc_2_5_wadr <= yt_rsc_2_5_i_wadr;
  yt_rsc_2_5_i_d_d <= yt_rsc_0_5_i_d_d_iff;
  yt_rsc_2_5_i_q_d <= yt_rsc_2_5_i_q_d_1;
  yt_rsc_2_5_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_2_5_i_wadr_d <= yt_rsc_0_5_i_wadr_d_iff;

  yt_rsc_2_6_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_77_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_2_6_clkr_en,
      clkw_en => yt_rsc_2_6_clkw_en,
      q => yt_rsc_2_6_i_q,
      radr => yt_rsc_2_6_i_radr,
      we => yt_rsc_2_6_we,
      d => yt_rsc_2_6_i_d,
      wadr => yt_rsc_2_6_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_2_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_2_0_i_clkr_en_d,
      d_d => yt_rsc_2_6_i_d_d,
      q_d => yt_rsc_2_6_i_q_d_1,
      radr_d => yt_rsc_2_6_i_radr_d,
      wadr_d => yt_rsc_2_6_i_wadr_d,
      we_d => yt_rsc_2_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_2_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_2_6_i_q <= yt_rsc_2_6_q;
  yt_rsc_2_6_radr <= yt_rsc_2_6_i_radr;
  yt_rsc_2_6_d <= yt_rsc_2_6_i_d;
  yt_rsc_2_6_wadr <= yt_rsc_2_6_i_wadr;
  yt_rsc_2_6_i_d_d <= yt_rsc_0_6_i_d_d_iff;
  yt_rsc_2_6_i_q_d <= yt_rsc_2_6_i_q_d_1;
  yt_rsc_2_6_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_2_6_i_wadr_d <= yt_rsc_0_6_i_wadr_d_iff;

  yt_rsc_2_7_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_78_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_2_7_clkr_en,
      clkw_en => yt_rsc_2_7_clkw_en,
      q => yt_rsc_2_7_i_q,
      radr => yt_rsc_2_7_i_radr,
      we => yt_rsc_2_7_we,
      d => yt_rsc_2_7_i_d,
      wadr => yt_rsc_2_7_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_2_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_2_0_i_clkr_en_d,
      d_d => yt_rsc_2_7_i_d_d,
      q_d => yt_rsc_2_7_i_q_d_1,
      radr_d => yt_rsc_2_7_i_radr_d,
      wadr_d => yt_rsc_2_7_i_wadr_d,
      we_d => yt_rsc_2_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_2_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_2_7_i_q <= yt_rsc_2_7_q;
  yt_rsc_2_7_radr <= yt_rsc_2_7_i_radr;
  yt_rsc_2_7_d <= yt_rsc_2_7_i_d;
  yt_rsc_2_7_wadr <= yt_rsc_2_7_i_wadr;
  yt_rsc_2_7_i_d_d <= yt_rsc_0_7_i_d_d_iff;
  yt_rsc_2_7_i_q_d <= yt_rsc_2_7_i_q_d_1;
  yt_rsc_2_7_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_2_7_i_wadr_d <= yt_rsc_0_0_i_wadr_d_iff;

  yt_rsc_2_8_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_79_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_2_8_clkr_en,
      clkw_en => yt_rsc_2_8_clkw_en,
      q => yt_rsc_2_8_i_q,
      radr => yt_rsc_2_8_i_radr,
      we => yt_rsc_2_8_we,
      d => yt_rsc_2_8_i_d,
      wadr => yt_rsc_2_8_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_2_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_2_0_i_clkr_en_d,
      d_d => yt_rsc_2_8_i_d_d,
      q_d => yt_rsc_2_8_i_q_d_1,
      radr_d => yt_rsc_2_8_i_radr_d,
      wadr_d => yt_rsc_2_8_i_wadr_d,
      we_d => yt_rsc_2_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_2_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_2_8_i_q <= yt_rsc_2_8_q;
  yt_rsc_2_8_radr <= yt_rsc_2_8_i_radr;
  yt_rsc_2_8_d <= yt_rsc_2_8_i_d;
  yt_rsc_2_8_wadr <= yt_rsc_2_8_i_wadr;
  yt_rsc_2_8_i_d_d <= yt_rsc_0_8_i_d_d_iff;
  yt_rsc_2_8_i_q_d <= yt_rsc_2_8_i_q_d_1;
  yt_rsc_2_8_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_2_8_i_wadr_d <= yt_rsc_0_1_i_wadr_d_iff;

  yt_rsc_2_9_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_80_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_2_9_clkr_en,
      clkw_en => yt_rsc_2_9_clkw_en,
      q => yt_rsc_2_9_i_q,
      radr => yt_rsc_2_9_i_radr,
      we => yt_rsc_2_9_we,
      d => yt_rsc_2_9_i_d,
      wadr => yt_rsc_2_9_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_2_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_2_0_i_clkr_en_d,
      d_d => yt_rsc_2_9_i_d_d,
      q_d => yt_rsc_2_9_i_q_d_1,
      radr_d => yt_rsc_2_9_i_radr_d,
      wadr_d => yt_rsc_2_9_i_wadr_d,
      we_d => yt_rsc_2_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_2_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_2_9_i_q <= yt_rsc_2_9_q;
  yt_rsc_2_9_radr <= yt_rsc_2_9_i_radr;
  yt_rsc_2_9_d <= yt_rsc_2_9_i_d;
  yt_rsc_2_9_wadr <= yt_rsc_2_9_i_wadr;
  yt_rsc_2_9_i_d_d <= yt_rsc_0_9_i_d_d_iff;
  yt_rsc_2_9_i_q_d <= yt_rsc_2_9_i_q_d_1;
  yt_rsc_2_9_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_2_9_i_wadr_d <= yt_rsc_0_2_i_wadr_d_iff;

  yt_rsc_2_10_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_81_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_2_10_clkr_en,
      clkw_en => yt_rsc_2_10_clkw_en,
      q => yt_rsc_2_10_i_q,
      radr => yt_rsc_2_10_i_radr,
      we => yt_rsc_2_10_we,
      d => yt_rsc_2_10_i_d,
      wadr => yt_rsc_2_10_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_2_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_2_0_i_clkr_en_d,
      d_d => yt_rsc_2_10_i_d_d,
      q_d => yt_rsc_2_10_i_q_d_1,
      radr_d => yt_rsc_2_10_i_radr_d,
      wadr_d => yt_rsc_2_10_i_wadr_d,
      we_d => yt_rsc_2_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_2_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_2_10_i_q <= yt_rsc_2_10_q;
  yt_rsc_2_10_radr <= yt_rsc_2_10_i_radr;
  yt_rsc_2_10_d <= yt_rsc_2_10_i_d;
  yt_rsc_2_10_wadr <= yt_rsc_2_10_i_wadr;
  yt_rsc_2_10_i_d_d <= yt_rsc_0_10_i_d_d_iff;
  yt_rsc_2_10_i_q_d <= yt_rsc_2_10_i_q_d_1;
  yt_rsc_2_10_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_2_10_i_wadr_d <= yt_rsc_0_10_i_wadr_d_iff;

  yt_rsc_2_11_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_82_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_2_11_clkr_en,
      clkw_en => yt_rsc_2_11_clkw_en,
      q => yt_rsc_2_11_i_q,
      radr => yt_rsc_2_11_i_radr,
      we => yt_rsc_2_11_we,
      d => yt_rsc_2_11_i_d,
      wadr => yt_rsc_2_11_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_2_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_2_0_i_clkr_en_d,
      d_d => yt_rsc_2_11_i_d_d,
      q_d => yt_rsc_2_11_i_q_d_1,
      radr_d => yt_rsc_2_11_i_radr_d,
      wadr_d => yt_rsc_2_11_i_wadr_d,
      we_d => yt_rsc_2_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_2_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_2_11_i_q <= yt_rsc_2_11_q;
  yt_rsc_2_11_radr <= yt_rsc_2_11_i_radr;
  yt_rsc_2_11_d <= yt_rsc_2_11_i_d;
  yt_rsc_2_11_wadr <= yt_rsc_2_11_i_wadr;
  yt_rsc_2_11_i_d_d <= yt_rsc_0_11_i_d_d_iff;
  yt_rsc_2_11_i_q_d <= yt_rsc_2_11_i_q_d_1;
  yt_rsc_2_11_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_2_11_i_wadr_d <= yt_rsc_0_11_i_wadr_d_iff;

  yt_rsc_2_12_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_83_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_2_12_clkr_en,
      clkw_en => yt_rsc_2_12_clkw_en,
      q => yt_rsc_2_12_i_q,
      radr => yt_rsc_2_12_i_radr,
      we => yt_rsc_2_12_we,
      d => yt_rsc_2_12_i_d,
      wadr => yt_rsc_2_12_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_2_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_2_0_i_clkr_en_d,
      d_d => yt_rsc_2_12_i_d_d,
      q_d => yt_rsc_2_12_i_q_d_1,
      radr_d => yt_rsc_2_12_i_radr_d,
      wadr_d => yt_rsc_2_12_i_wadr_d,
      we_d => yt_rsc_2_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_2_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_2_12_i_q <= yt_rsc_2_12_q;
  yt_rsc_2_12_radr <= yt_rsc_2_12_i_radr;
  yt_rsc_2_12_d <= yt_rsc_2_12_i_d;
  yt_rsc_2_12_wadr <= yt_rsc_2_12_i_wadr;
  yt_rsc_2_12_i_d_d <= yt_rsc_0_12_i_d_d_iff;
  yt_rsc_2_12_i_q_d <= yt_rsc_2_12_i_q_d_1;
  yt_rsc_2_12_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_2_12_i_wadr_d <= yt_rsc_0_3_i_wadr_d_iff;

  yt_rsc_2_13_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_84_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_2_13_clkr_en,
      clkw_en => yt_rsc_2_13_clkw_en,
      q => yt_rsc_2_13_i_q,
      radr => yt_rsc_2_13_i_radr,
      we => yt_rsc_2_13_we,
      d => yt_rsc_2_13_i_d,
      wadr => yt_rsc_2_13_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_2_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_2_0_i_clkr_en_d,
      d_d => yt_rsc_2_13_i_d_d,
      q_d => yt_rsc_2_13_i_q_d_1,
      radr_d => yt_rsc_2_13_i_radr_d,
      wadr_d => yt_rsc_2_13_i_wadr_d,
      we_d => yt_rsc_2_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_2_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_2_13_i_q <= yt_rsc_2_13_q;
  yt_rsc_2_13_radr <= yt_rsc_2_13_i_radr;
  yt_rsc_2_13_d <= yt_rsc_2_13_i_d;
  yt_rsc_2_13_wadr <= yt_rsc_2_13_i_wadr;
  yt_rsc_2_13_i_d_d <= yt_rsc_0_13_i_d_d_iff;
  yt_rsc_2_13_i_q_d <= yt_rsc_2_13_i_q_d_1;
  yt_rsc_2_13_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_2_13_i_wadr_d <= yt_rsc_0_4_i_wadr_d_iff;

  yt_rsc_2_14_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_85_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_2_14_clkr_en,
      clkw_en => yt_rsc_2_14_clkw_en,
      q => yt_rsc_2_14_i_q,
      radr => yt_rsc_2_14_i_radr,
      we => yt_rsc_2_14_we,
      d => yt_rsc_2_14_i_d,
      wadr => yt_rsc_2_14_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_2_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_2_0_i_clkr_en_d,
      d_d => yt_rsc_2_14_i_d_d,
      q_d => yt_rsc_2_14_i_q_d_1,
      radr_d => yt_rsc_2_14_i_radr_d,
      wadr_d => yt_rsc_2_14_i_wadr_d,
      we_d => yt_rsc_2_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_2_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_2_14_i_q <= yt_rsc_2_14_q;
  yt_rsc_2_14_radr <= yt_rsc_2_14_i_radr;
  yt_rsc_2_14_d <= yt_rsc_2_14_i_d;
  yt_rsc_2_14_wadr <= yt_rsc_2_14_i_wadr;
  yt_rsc_2_14_i_d_d <= yt_rsc_0_14_i_d_d_iff;
  yt_rsc_2_14_i_q_d <= yt_rsc_2_14_i_q_d_1;
  yt_rsc_2_14_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_2_14_i_wadr_d <= yt_rsc_0_5_i_wadr_d_iff;

  yt_rsc_2_15_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_86_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_2_15_clkr_en,
      clkw_en => yt_rsc_2_15_clkw_en,
      q => yt_rsc_2_15_i_q,
      radr => yt_rsc_2_15_i_radr,
      we => yt_rsc_2_15_we,
      d => yt_rsc_2_15_i_d,
      wadr => yt_rsc_2_15_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_2_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_2_0_i_clkr_en_d,
      d_d => yt_rsc_2_15_i_d_d,
      q_d => yt_rsc_2_15_i_q_d_1,
      radr_d => yt_rsc_2_15_i_radr_d,
      wadr_d => yt_rsc_2_15_i_wadr_d,
      we_d => yt_rsc_2_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_2_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_2_15_i_q <= yt_rsc_2_15_q;
  yt_rsc_2_15_radr <= yt_rsc_2_15_i_radr;
  yt_rsc_2_15_d <= yt_rsc_2_15_i_d;
  yt_rsc_2_15_wadr <= yt_rsc_2_15_i_wadr;
  yt_rsc_2_15_i_d_d <= yt_rsc_0_15_i_d_d_iff;
  yt_rsc_2_15_i_q_d <= yt_rsc_2_15_i_q_d_1;
  yt_rsc_2_15_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_2_15_i_wadr_d <= yt_rsc_0_6_i_wadr_d_iff;

  yt_rsc_2_16_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_87_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_2_16_clkr_en,
      clkw_en => yt_rsc_2_16_clkw_en,
      q => yt_rsc_2_16_i_q,
      radr => yt_rsc_2_16_i_radr,
      we => yt_rsc_2_16_we,
      d => yt_rsc_2_16_i_d,
      wadr => yt_rsc_2_16_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_2_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_2_16_i_clkr_en_d,
      d_d => yt_rsc_2_16_i_d_d,
      q_d => yt_rsc_2_16_i_q_d_1,
      radr_d => yt_rsc_2_16_i_radr_d,
      wadr_d => yt_rsc_2_16_i_wadr_d,
      we_d => yt_rsc_2_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_2_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_2_16_i_q <= yt_rsc_2_16_q;
  yt_rsc_2_16_radr <= yt_rsc_2_16_i_radr;
  yt_rsc_2_16_d <= yt_rsc_2_16_i_d;
  yt_rsc_2_16_wadr <= yt_rsc_2_16_i_wadr;
  yt_rsc_2_16_i_d_d <= yt_rsc_0_0_i_d_d_iff;
  yt_rsc_2_16_i_q_d <= yt_rsc_2_16_i_q_d_1;
  yt_rsc_2_16_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_2_16_i_wadr_d <= yt_rsc_0_0_i_wadr_d_iff;

  yt_rsc_2_17_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_88_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_2_17_clkr_en,
      clkw_en => yt_rsc_2_17_clkw_en,
      q => yt_rsc_2_17_i_q,
      radr => yt_rsc_2_17_i_radr,
      we => yt_rsc_2_17_we,
      d => yt_rsc_2_17_i_d,
      wadr => yt_rsc_2_17_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_2_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_2_16_i_clkr_en_d,
      d_d => yt_rsc_2_17_i_d_d,
      q_d => yt_rsc_2_17_i_q_d_1,
      radr_d => yt_rsc_2_17_i_radr_d,
      wadr_d => yt_rsc_2_17_i_wadr_d,
      we_d => yt_rsc_2_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_2_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_2_17_i_q <= yt_rsc_2_17_q;
  yt_rsc_2_17_radr <= yt_rsc_2_17_i_radr;
  yt_rsc_2_17_d <= yt_rsc_2_17_i_d;
  yt_rsc_2_17_wadr <= yt_rsc_2_17_i_wadr;
  yt_rsc_2_17_i_d_d <= yt_rsc_0_1_i_d_d_iff;
  yt_rsc_2_17_i_q_d <= yt_rsc_2_17_i_q_d_1;
  yt_rsc_2_17_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_2_17_i_wadr_d <= yt_rsc_0_1_i_wadr_d_iff;

  yt_rsc_2_18_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_89_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_2_18_clkr_en,
      clkw_en => yt_rsc_2_18_clkw_en,
      q => yt_rsc_2_18_i_q,
      radr => yt_rsc_2_18_i_radr,
      we => yt_rsc_2_18_we,
      d => yt_rsc_2_18_i_d,
      wadr => yt_rsc_2_18_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_2_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_2_16_i_clkr_en_d,
      d_d => yt_rsc_2_18_i_d_d,
      q_d => yt_rsc_2_18_i_q_d_1,
      radr_d => yt_rsc_2_18_i_radr_d,
      wadr_d => yt_rsc_2_18_i_wadr_d,
      we_d => yt_rsc_2_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_2_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_2_18_i_q <= yt_rsc_2_18_q;
  yt_rsc_2_18_radr <= yt_rsc_2_18_i_radr;
  yt_rsc_2_18_d <= yt_rsc_2_18_i_d;
  yt_rsc_2_18_wadr <= yt_rsc_2_18_i_wadr;
  yt_rsc_2_18_i_d_d <= yt_rsc_0_2_i_d_d_iff;
  yt_rsc_2_18_i_q_d <= yt_rsc_2_18_i_q_d_1;
  yt_rsc_2_18_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_2_18_i_wadr_d <= yt_rsc_0_2_i_wadr_d_iff;

  yt_rsc_2_19_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_90_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_2_19_clkr_en,
      clkw_en => yt_rsc_2_19_clkw_en,
      q => yt_rsc_2_19_i_q,
      radr => yt_rsc_2_19_i_radr,
      we => yt_rsc_2_19_we,
      d => yt_rsc_2_19_i_d,
      wadr => yt_rsc_2_19_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_2_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_2_16_i_clkr_en_d,
      d_d => yt_rsc_2_19_i_d_d,
      q_d => yt_rsc_2_19_i_q_d_1,
      radr_d => yt_rsc_2_19_i_radr_d,
      wadr_d => yt_rsc_2_19_i_wadr_d,
      we_d => yt_rsc_2_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_2_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_2_19_i_q <= yt_rsc_2_19_q;
  yt_rsc_2_19_radr <= yt_rsc_2_19_i_radr;
  yt_rsc_2_19_d <= yt_rsc_2_19_i_d;
  yt_rsc_2_19_wadr <= yt_rsc_2_19_i_wadr;
  yt_rsc_2_19_i_d_d <= yt_rsc_0_3_i_d_d_iff;
  yt_rsc_2_19_i_q_d <= yt_rsc_2_19_i_q_d_1;
  yt_rsc_2_19_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_2_19_i_wadr_d <= yt_rsc_0_3_i_wadr_d_iff;

  yt_rsc_2_20_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_91_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_2_20_clkr_en,
      clkw_en => yt_rsc_2_20_clkw_en,
      q => yt_rsc_2_20_i_q,
      radr => yt_rsc_2_20_i_radr,
      we => yt_rsc_2_20_we,
      d => yt_rsc_2_20_i_d,
      wadr => yt_rsc_2_20_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_2_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_2_16_i_clkr_en_d,
      d_d => yt_rsc_2_20_i_d_d,
      q_d => yt_rsc_2_20_i_q_d_1,
      radr_d => yt_rsc_2_20_i_radr_d,
      wadr_d => yt_rsc_2_20_i_wadr_d,
      we_d => yt_rsc_2_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_2_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_2_20_i_q <= yt_rsc_2_20_q;
  yt_rsc_2_20_radr <= yt_rsc_2_20_i_radr;
  yt_rsc_2_20_d <= yt_rsc_2_20_i_d;
  yt_rsc_2_20_wadr <= yt_rsc_2_20_i_wadr;
  yt_rsc_2_20_i_d_d <= yt_rsc_0_4_i_d_d_iff;
  yt_rsc_2_20_i_q_d <= yt_rsc_2_20_i_q_d_1;
  yt_rsc_2_20_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_2_20_i_wadr_d <= yt_rsc_0_4_i_wadr_d_iff;

  yt_rsc_2_21_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_92_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_2_21_clkr_en,
      clkw_en => yt_rsc_2_21_clkw_en,
      q => yt_rsc_2_21_i_q,
      radr => yt_rsc_2_21_i_radr,
      we => yt_rsc_2_21_we,
      d => yt_rsc_2_21_i_d,
      wadr => yt_rsc_2_21_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_2_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_2_16_i_clkr_en_d,
      d_d => yt_rsc_2_21_i_d_d,
      q_d => yt_rsc_2_21_i_q_d_1,
      radr_d => yt_rsc_2_21_i_radr_d,
      wadr_d => yt_rsc_2_21_i_wadr_d,
      we_d => yt_rsc_2_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_2_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_2_21_i_q <= yt_rsc_2_21_q;
  yt_rsc_2_21_radr <= yt_rsc_2_21_i_radr;
  yt_rsc_2_21_d <= yt_rsc_2_21_i_d;
  yt_rsc_2_21_wadr <= yt_rsc_2_21_i_wadr;
  yt_rsc_2_21_i_d_d <= yt_rsc_0_5_i_d_d_iff;
  yt_rsc_2_21_i_q_d <= yt_rsc_2_21_i_q_d_1;
  yt_rsc_2_21_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_2_21_i_wadr_d <= yt_rsc_0_5_i_wadr_d_iff;

  yt_rsc_2_22_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_93_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_2_22_clkr_en,
      clkw_en => yt_rsc_2_22_clkw_en,
      q => yt_rsc_2_22_i_q,
      radr => yt_rsc_2_22_i_radr,
      we => yt_rsc_2_22_we,
      d => yt_rsc_2_22_i_d,
      wadr => yt_rsc_2_22_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_2_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_2_16_i_clkr_en_d,
      d_d => yt_rsc_2_22_i_d_d,
      q_d => yt_rsc_2_22_i_q_d_1,
      radr_d => yt_rsc_2_22_i_radr_d,
      wadr_d => yt_rsc_2_22_i_wadr_d,
      we_d => yt_rsc_2_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_2_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_2_22_i_q <= yt_rsc_2_22_q;
  yt_rsc_2_22_radr <= yt_rsc_2_22_i_radr;
  yt_rsc_2_22_d <= yt_rsc_2_22_i_d;
  yt_rsc_2_22_wadr <= yt_rsc_2_22_i_wadr;
  yt_rsc_2_22_i_d_d <= yt_rsc_0_6_i_d_d_iff;
  yt_rsc_2_22_i_q_d <= yt_rsc_2_22_i_q_d_1;
  yt_rsc_2_22_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_2_22_i_wadr_d <= yt_rsc_0_6_i_wadr_d_iff;

  yt_rsc_2_23_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_94_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_2_23_clkr_en,
      clkw_en => yt_rsc_2_23_clkw_en,
      q => yt_rsc_2_23_i_q,
      radr => yt_rsc_2_23_i_radr,
      we => yt_rsc_2_23_we,
      d => yt_rsc_2_23_i_d,
      wadr => yt_rsc_2_23_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_2_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_2_16_i_clkr_en_d,
      d_d => yt_rsc_2_23_i_d_d,
      q_d => yt_rsc_2_23_i_q_d_1,
      radr_d => yt_rsc_2_23_i_radr_d,
      wadr_d => yt_rsc_2_23_i_wadr_d,
      we_d => yt_rsc_2_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_2_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_2_23_i_q <= yt_rsc_2_23_q;
  yt_rsc_2_23_radr <= yt_rsc_2_23_i_radr;
  yt_rsc_2_23_d <= yt_rsc_2_23_i_d;
  yt_rsc_2_23_wadr <= yt_rsc_2_23_i_wadr;
  yt_rsc_2_23_i_d_d <= yt_rsc_0_7_i_d_d_iff;
  yt_rsc_2_23_i_q_d <= yt_rsc_2_23_i_q_d_1;
  yt_rsc_2_23_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_2_23_i_wadr_d <= yt_rsc_0_0_i_wadr_d_iff;

  yt_rsc_2_24_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_95_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_2_24_clkr_en,
      clkw_en => yt_rsc_2_24_clkw_en,
      q => yt_rsc_2_24_i_q,
      radr => yt_rsc_2_24_i_radr,
      we => yt_rsc_2_24_we,
      d => yt_rsc_2_24_i_d,
      wadr => yt_rsc_2_24_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_2_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_2_16_i_clkr_en_d,
      d_d => yt_rsc_2_24_i_d_d,
      q_d => yt_rsc_2_24_i_q_d_1,
      radr_d => yt_rsc_2_24_i_radr_d,
      wadr_d => yt_rsc_2_24_i_wadr_d,
      we_d => yt_rsc_2_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_2_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_2_24_i_q <= yt_rsc_2_24_q;
  yt_rsc_2_24_radr <= yt_rsc_2_24_i_radr;
  yt_rsc_2_24_d <= yt_rsc_2_24_i_d;
  yt_rsc_2_24_wadr <= yt_rsc_2_24_i_wadr;
  yt_rsc_2_24_i_d_d <= yt_rsc_0_8_i_d_d_iff;
  yt_rsc_2_24_i_q_d <= yt_rsc_2_24_i_q_d_1;
  yt_rsc_2_24_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_2_24_i_wadr_d <= yt_rsc_0_1_i_wadr_d_iff;

  yt_rsc_2_25_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_96_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_2_25_clkr_en,
      clkw_en => yt_rsc_2_25_clkw_en,
      q => yt_rsc_2_25_i_q,
      radr => yt_rsc_2_25_i_radr,
      we => yt_rsc_2_25_we,
      d => yt_rsc_2_25_i_d,
      wadr => yt_rsc_2_25_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_2_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_2_16_i_clkr_en_d,
      d_d => yt_rsc_2_25_i_d_d,
      q_d => yt_rsc_2_25_i_q_d_1,
      radr_d => yt_rsc_2_25_i_radr_d,
      wadr_d => yt_rsc_2_25_i_wadr_d,
      we_d => yt_rsc_2_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_2_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_2_25_i_q <= yt_rsc_2_25_q;
  yt_rsc_2_25_radr <= yt_rsc_2_25_i_radr;
  yt_rsc_2_25_d <= yt_rsc_2_25_i_d;
  yt_rsc_2_25_wadr <= yt_rsc_2_25_i_wadr;
  yt_rsc_2_25_i_d_d <= yt_rsc_0_9_i_d_d_iff;
  yt_rsc_2_25_i_q_d <= yt_rsc_2_25_i_q_d_1;
  yt_rsc_2_25_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_2_25_i_wadr_d <= yt_rsc_0_2_i_wadr_d_iff;

  yt_rsc_2_26_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_97_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_2_26_clkr_en,
      clkw_en => yt_rsc_2_26_clkw_en,
      q => yt_rsc_2_26_i_q,
      radr => yt_rsc_2_26_i_radr,
      we => yt_rsc_2_26_we,
      d => yt_rsc_2_26_i_d,
      wadr => yt_rsc_2_26_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_2_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_2_16_i_clkr_en_d,
      d_d => yt_rsc_2_26_i_d_d,
      q_d => yt_rsc_2_26_i_q_d_1,
      radr_d => yt_rsc_2_26_i_radr_d,
      wadr_d => yt_rsc_2_26_i_wadr_d,
      we_d => yt_rsc_2_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_2_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_2_26_i_q <= yt_rsc_2_26_q;
  yt_rsc_2_26_radr <= yt_rsc_2_26_i_radr;
  yt_rsc_2_26_d <= yt_rsc_2_26_i_d;
  yt_rsc_2_26_wadr <= yt_rsc_2_26_i_wadr;
  yt_rsc_2_26_i_d_d <= yt_rsc_0_10_i_d_d_iff;
  yt_rsc_2_26_i_q_d <= yt_rsc_2_26_i_q_d_1;
  yt_rsc_2_26_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_2_26_i_wadr_d <= yt_rsc_0_10_i_wadr_d_iff;

  yt_rsc_2_27_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_98_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_2_27_clkr_en,
      clkw_en => yt_rsc_2_27_clkw_en,
      q => yt_rsc_2_27_i_q,
      radr => yt_rsc_2_27_i_radr,
      we => yt_rsc_2_27_we,
      d => yt_rsc_2_27_i_d,
      wadr => yt_rsc_2_27_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_2_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_2_16_i_clkr_en_d,
      d_d => yt_rsc_2_27_i_d_d,
      q_d => yt_rsc_2_27_i_q_d_1,
      radr_d => yt_rsc_2_27_i_radr_d,
      wadr_d => yt_rsc_2_27_i_wadr_d,
      we_d => yt_rsc_2_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_2_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_2_27_i_q <= yt_rsc_2_27_q;
  yt_rsc_2_27_radr <= yt_rsc_2_27_i_radr;
  yt_rsc_2_27_d <= yt_rsc_2_27_i_d;
  yt_rsc_2_27_wadr <= yt_rsc_2_27_i_wadr;
  yt_rsc_2_27_i_d_d <= yt_rsc_0_11_i_d_d_iff;
  yt_rsc_2_27_i_q_d <= yt_rsc_2_27_i_q_d_1;
  yt_rsc_2_27_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_2_27_i_wadr_d <= yt_rsc_0_11_i_wadr_d_iff;

  yt_rsc_2_28_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_99_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_2_28_clkr_en,
      clkw_en => yt_rsc_2_28_clkw_en,
      q => yt_rsc_2_28_i_q,
      radr => yt_rsc_2_28_i_radr,
      we => yt_rsc_2_28_we,
      d => yt_rsc_2_28_i_d,
      wadr => yt_rsc_2_28_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_2_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_2_16_i_clkr_en_d,
      d_d => yt_rsc_2_28_i_d_d,
      q_d => yt_rsc_2_28_i_q_d_1,
      radr_d => yt_rsc_2_28_i_radr_d,
      wadr_d => yt_rsc_2_28_i_wadr_d,
      we_d => yt_rsc_2_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_2_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_2_28_i_q <= yt_rsc_2_28_q;
  yt_rsc_2_28_radr <= yt_rsc_2_28_i_radr;
  yt_rsc_2_28_d <= yt_rsc_2_28_i_d;
  yt_rsc_2_28_wadr <= yt_rsc_2_28_i_wadr;
  yt_rsc_2_28_i_d_d <= yt_rsc_0_12_i_d_d_iff;
  yt_rsc_2_28_i_q_d <= yt_rsc_2_28_i_q_d_1;
  yt_rsc_2_28_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_2_28_i_wadr_d <= yt_rsc_0_3_i_wadr_d_iff;

  yt_rsc_2_29_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_100_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_2_29_clkr_en,
      clkw_en => yt_rsc_2_29_clkw_en,
      q => yt_rsc_2_29_i_q,
      radr => yt_rsc_2_29_i_radr,
      we => yt_rsc_2_29_we,
      d => yt_rsc_2_29_i_d,
      wadr => yt_rsc_2_29_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_2_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_2_16_i_clkr_en_d,
      d_d => yt_rsc_2_29_i_d_d,
      q_d => yt_rsc_2_29_i_q_d_1,
      radr_d => yt_rsc_2_29_i_radr_d,
      wadr_d => yt_rsc_2_29_i_wadr_d,
      we_d => yt_rsc_2_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_2_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_2_29_i_q <= yt_rsc_2_29_q;
  yt_rsc_2_29_radr <= yt_rsc_2_29_i_radr;
  yt_rsc_2_29_d <= yt_rsc_2_29_i_d;
  yt_rsc_2_29_wadr <= yt_rsc_2_29_i_wadr;
  yt_rsc_2_29_i_d_d <= yt_rsc_0_13_i_d_d_iff;
  yt_rsc_2_29_i_q_d <= yt_rsc_2_29_i_q_d_1;
  yt_rsc_2_29_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_2_29_i_wadr_d <= yt_rsc_0_4_i_wadr_d_iff;

  yt_rsc_2_30_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_101_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_2_30_clkr_en,
      clkw_en => yt_rsc_2_30_clkw_en,
      q => yt_rsc_2_30_i_q,
      radr => yt_rsc_2_30_i_radr,
      we => yt_rsc_2_30_we,
      d => yt_rsc_2_30_i_d,
      wadr => yt_rsc_2_30_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_2_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_2_16_i_clkr_en_d,
      d_d => yt_rsc_2_30_i_d_d,
      q_d => yt_rsc_2_30_i_q_d_1,
      radr_d => yt_rsc_2_30_i_radr_d,
      wadr_d => yt_rsc_2_30_i_wadr_d,
      we_d => yt_rsc_2_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_2_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_2_30_i_q <= yt_rsc_2_30_q;
  yt_rsc_2_30_radr <= yt_rsc_2_30_i_radr;
  yt_rsc_2_30_d <= yt_rsc_2_30_i_d;
  yt_rsc_2_30_wadr <= yt_rsc_2_30_i_wadr;
  yt_rsc_2_30_i_d_d <= yt_rsc_0_14_i_d_d_iff;
  yt_rsc_2_30_i_q_d <= yt_rsc_2_30_i_q_d_1;
  yt_rsc_2_30_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_2_30_i_wadr_d <= yt_rsc_0_5_i_wadr_d_iff;

  yt_rsc_2_31_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_102_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_2_31_clkr_en,
      clkw_en => yt_rsc_2_31_clkw_en,
      q => yt_rsc_2_31_i_q,
      radr => yt_rsc_2_31_i_radr,
      we => yt_rsc_2_31_we,
      d => yt_rsc_2_31_i_d,
      wadr => yt_rsc_2_31_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_2_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_2_16_i_clkr_en_d,
      d_d => yt_rsc_2_31_i_d_d,
      q_d => yt_rsc_2_31_i_q_d_1,
      radr_d => yt_rsc_2_31_i_radr_d,
      wadr_d => yt_rsc_2_31_i_wadr_d,
      we_d => yt_rsc_2_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_2_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_2_31_i_q <= yt_rsc_2_31_q;
  yt_rsc_2_31_radr <= yt_rsc_2_31_i_radr;
  yt_rsc_2_31_d <= yt_rsc_2_31_i_d;
  yt_rsc_2_31_wadr <= yt_rsc_2_31_i_wadr;
  yt_rsc_2_31_i_d_d <= yt_rsc_0_15_i_d_d_iff;
  yt_rsc_2_31_i_q_d <= yt_rsc_2_31_i_q_d_1;
  yt_rsc_2_31_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_2_31_i_wadr_d <= yt_rsc_0_6_i_wadr_d_iff;

  yt_rsc_3_0_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_103_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_3_0_clkr_en,
      clkw_en => yt_rsc_3_0_clkw_en,
      q => yt_rsc_3_0_i_q,
      radr => yt_rsc_3_0_i_radr,
      we => yt_rsc_3_0_we,
      d => yt_rsc_3_0_i_d,
      wadr => yt_rsc_3_0_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_3_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_3_0_i_clkr_en_d,
      d_d => yt_rsc_3_0_i_d_d,
      q_d => yt_rsc_3_0_i_q_d_1,
      radr_d => yt_rsc_3_0_i_radr_d,
      wadr_d => yt_rsc_3_0_i_wadr_d,
      we_d => yt_rsc_3_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_3_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_3_0_i_q <= yt_rsc_3_0_q;
  yt_rsc_3_0_radr <= yt_rsc_3_0_i_radr;
  yt_rsc_3_0_d <= yt_rsc_3_0_i_d;
  yt_rsc_3_0_wadr <= yt_rsc_3_0_i_wadr;
  yt_rsc_3_0_i_d_d <= yt_rsc_0_0_i_d_d_iff;
  yt_rsc_3_0_i_q_d <= yt_rsc_3_0_i_q_d_1;
  yt_rsc_3_0_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_3_0_i_wadr_d <= yt_rsc_0_0_i_wadr_d_iff;

  yt_rsc_3_1_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_104_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_3_1_clkr_en,
      clkw_en => yt_rsc_3_1_clkw_en,
      q => yt_rsc_3_1_i_q,
      radr => yt_rsc_3_1_i_radr,
      we => yt_rsc_3_1_we,
      d => yt_rsc_3_1_i_d,
      wadr => yt_rsc_3_1_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_3_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_3_0_i_clkr_en_d,
      d_d => yt_rsc_3_1_i_d_d,
      q_d => yt_rsc_3_1_i_q_d_1,
      radr_d => yt_rsc_3_1_i_radr_d,
      wadr_d => yt_rsc_3_1_i_wadr_d,
      we_d => yt_rsc_3_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_3_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_3_1_i_q <= yt_rsc_3_1_q;
  yt_rsc_3_1_radr <= yt_rsc_3_1_i_radr;
  yt_rsc_3_1_d <= yt_rsc_3_1_i_d;
  yt_rsc_3_1_wadr <= yt_rsc_3_1_i_wadr;
  yt_rsc_3_1_i_d_d <= yt_rsc_0_1_i_d_d_iff;
  yt_rsc_3_1_i_q_d <= yt_rsc_3_1_i_q_d_1;
  yt_rsc_3_1_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_3_1_i_wadr_d <= yt_rsc_0_1_i_wadr_d_iff;

  yt_rsc_3_2_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_105_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_3_2_clkr_en,
      clkw_en => yt_rsc_3_2_clkw_en,
      q => yt_rsc_3_2_i_q,
      radr => yt_rsc_3_2_i_radr,
      we => yt_rsc_3_2_we,
      d => yt_rsc_3_2_i_d,
      wadr => yt_rsc_3_2_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_3_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_3_0_i_clkr_en_d,
      d_d => yt_rsc_3_2_i_d_d,
      q_d => yt_rsc_3_2_i_q_d_1,
      radr_d => yt_rsc_3_2_i_radr_d,
      wadr_d => yt_rsc_3_2_i_wadr_d,
      we_d => yt_rsc_3_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_3_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_3_2_i_q <= yt_rsc_3_2_q;
  yt_rsc_3_2_radr <= yt_rsc_3_2_i_radr;
  yt_rsc_3_2_d <= yt_rsc_3_2_i_d;
  yt_rsc_3_2_wadr <= yt_rsc_3_2_i_wadr;
  yt_rsc_3_2_i_d_d <= yt_rsc_0_2_i_d_d_iff;
  yt_rsc_3_2_i_q_d <= yt_rsc_3_2_i_q_d_1;
  yt_rsc_3_2_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_3_2_i_wadr_d <= yt_rsc_0_2_i_wadr_d_iff;

  yt_rsc_3_3_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_106_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_3_3_clkr_en,
      clkw_en => yt_rsc_3_3_clkw_en,
      q => yt_rsc_3_3_i_q,
      radr => yt_rsc_3_3_i_radr,
      we => yt_rsc_3_3_we,
      d => yt_rsc_3_3_i_d,
      wadr => yt_rsc_3_3_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_3_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_3_0_i_clkr_en_d,
      d_d => yt_rsc_3_3_i_d_d,
      q_d => yt_rsc_3_3_i_q_d_1,
      radr_d => yt_rsc_3_3_i_radr_d,
      wadr_d => yt_rsc_3_3_i_wadr_d,
      we_d => yt_rsc_3_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_3_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_3_3_i_q <= yt_rsc_3_3_q;
  yt_rsc_3_3_radr <= yt_rsc_3_3_i_radr;
  yt_rsc_3_3_d <= yt_rsc_3_3_i_d;
  yt_rsc_3_3_wadr <= yt_rsc_3_3_i_wadr;
  yt_rsc_3_3_i_d_d <= yt_rsc_0_3_i_d_d_iff;
  yt_rsc_3_3_i_q_d <= yt_rsc_3_3_i_q_d_1;
  yt_rsc_3_3_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_3_3_i_wadr_d <= yt_rsc_0_3_i_wadr_d_iff;

  yt_rsc_3_4_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_107_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_3_4_clkr_en,
      clkw_en => yt_rsc_3_4_clkw_en,
      q => yt_rsc_3_4_i_q,
      radr => yt_rsc_3_4_i_radr,
      we => yt_rsc_3_4_we,
      d => yt_rsc_3_4_i_d,
      wadr => yt_rsc_3_4_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_3_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_3_0_i_clkr_en_d,
      d_d => yt_rsc_3_4_i_d_d,
      q_d => yt_rsc_3_4_i_q_d_1,
      radr_d => yt_rsc_3_4_i_radr_d,
      wadr_d => yt_rsc_3_4_i_wadr_d,
      we_d => yt_rsc_3_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_3_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_3_4_i_q <= yt_rsc_3_4_q;
  yt_rsc_3_4_radr <= yt_rsc_3_4_i_radr;
  yt_rsc_3_4_d <= yt_rsc_3_4_i_d;
  yt_rsc_3_4_wadr <= yt_rsc_3_4_i_wadr;
  yt_rsc_3_4_i_d_d <= yt_rsc_0_4_i_d_d_iff;
  yt_rsc_3_4_i_q_d <= yt_rsc_3_4_i_q_d_1;
  yt_rsc_3_4_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_3_4_i_wadr_d <= yt_rsc_0_4_i_wadr_d_iff;

  yt_rsc_3_5_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_108_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_3_5_clkr_en,
      clkw_en => yt_rsc_3_5_clkw_en,
      q => yt_rsc_3_5_i_q,
      radr => yt_rsc_3_5_i_radr,
      we => yt_rsc_3_5_we,
      d => yt_rsc_3_5_i_d,
      wadr => yt_rsc_3_5_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_3_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_3_0_i_clkr_en_d,
      d_d => yt_rsc_3_5_i_d_d,
      q_d => yt_rsc_3_5_i_q_d_1,
      radr_d => yt_rsc_3_5_i_radr_d,
      wadr_d => yt_rsc_3_5_i_wadr_d,
      we_d => yt_rsc_3_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_3_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_3_5_i_q <= yt_rsc_3_5_q;
  yt_rsc_3_5_radr <= yt_rsc_3_5_i_radr;
  yt_rsc_3_5_d <= yt_rsc_3_5_i_d;
  yt_rsc_3_5_wadr <= yt_rsc_3_5_i_wadr;
  yt_rsc_3_5_i_d_d <= yt_rsc_0_5_i_d_d_iff;
  yt_rsc_3_5_i_q_d <= yt_rsc_3_5_i_q_d_1;
  yt_rsc_3_5_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_3_5_i_wadr_d <= yt_rsc_0_5_i_wadr_d_iff;

  yt_rsc_3_6_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_109_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_3_6_clkr_en,
      clkw_en => yt_rsc_3_6_clkw_en,
      q => yt_rsc_3_6_i_q,
      radr => yt_rsc_3_6_i_radr,
      we => yt_rsc_3_6_we,
      d => yt_rsc_3_6_i_d,
      wadr => yt_rsc_3_6_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_3_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_3_0_i_clkr_en_d,
      d_d => yt_rsc_3_6_i_d_d,
      q_d => yt_rsc_3_6_i_q_d_1,
      radr_d => yt_rsc_3_6_i_radr_d,
      wadr_d => yt_rsc_3_6_i_wadr_d,
      we_d => yt_rsc_3_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_3_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_3_6_i_q <= yt_rsc_3_6_q;
  yt_rsc_3_6_radr <= yt_rsc_3_6_i_radr;
  yt_rsc_3_6_d <= yt_rsc_3_6_i_d;
  yt_rsc_3_6_wadr <= yt_rsc_3_6_i_wadr;
  yt_rsc_3_6_i_d_d <= yt_rsc_0_6_i_d_d_iff;
  yt_rsc_3_6_i_q_d <= yt_rsc_3_6_i_q_d_1;
  yt_rsc_3_6_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_3_6_i_wadr_d <= yt_rsc_0_6_i_wadr_d_iff;

  yt_rsc_3_7_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_110_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_3_7_clkr_en,
      clkw_en => yt_rsc_3_7_clkw_en,
      q => yt_rsc_3_7_i_q,
      radr => yt_rsc_3_7_i_radr,
      we => yt_rsc_3_7_we,
      d => yt_rsc_3_7_i_d,
      wadr => yt_rsc_3_7_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_3_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_3_0_i_clkr_en_d,
      d_d => yt_rsc_3_7_i_d_d,
      q_d => yt_rsc_3_7_i_q_d_1,
      radr_d => yt_rsc_3_7_i_radr_d,
      wadr_d => yt_rsc_3_7_i_wadr_d,
      we_d => yt_rsc_3_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_3_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_3_7_i_q <= yt_rsc_3_7_q;
  yt_rsc_3_7_radr <= yt_rsc_3_7_i_radr;
  yt_rsc_3_7_d <= yt_rsc_3_7_i_d;
  yt_rsc_3_7_wadr <= yt_rsc_3_7_i_wadr;
  yt_rsc_3_7_i_d_d <= yt_rsc_0_7_i_d_d_iff;
  yt_rsc_3_7_i_q_d <= yt_rsc_3_7_i_q_d_1;
  yt_rsc_3_7_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_3_7_i_wadr_d <= yt_rsc_0_0_i_wadr_d_iff;

  yt_rsc_3_8_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_111_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_3_8_clkr_en,
      clkw_en => yt_rsc_3_8_clkw_en,
      q => yt_rsc_3_8_i_q,
      radr => yt_rsc_3_8_i_radr,
      we => yt_rsc_3_8_we,
      d => yt_rsc_3_8_i_d,
      wadr => yt_rsc_3_8_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_3_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_3_0_i_clkr_en_d,
      d_d => yt_rsc_3_8_i_d_d,
      q_d => yt_rsc_3_8_i_q_d_1,
      radr_d => yt_rsc_3_8_i_radr_d,
      wadr_d => yt_rsc_3_8_i_wadr_d,
      we_d => yt_rsc_3_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_3_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_3_8_i_q <= yt_rsc_3_8_q;
  yt_rsc_3_8_radr <= yt_rsc_3_8_i_radr;
  yt_rsc_3_8_d <= yt_rsc_3_8_i_d;
  yt_rsc_3_8_wadr <= yt_rsc_3_8_i_wadr;
  yt_rsc_3_8_i_d_d <= yt_rsc_0_8_i_d_d_iff;
  yt_rsc_3_8_i_q_d <= yt_rsc_3_8_i_q_d_1;
  yt_rsc_3_8_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_3_8_i_wadr_d <= yt_rsc_0_1_i_wadr_d_iff;

  yt_rsc_3_9_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_112_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_3_9_clkr_en,
      clkw_en => yt_rsc_3_9_clkw_en,
      q => yt_rsc_3_9_i_q,
      radr => yt_rsc_3_9_i_radr,
      we => yt_rsc_3_9_we,
      d => yt_rsc_3_9_i_d,
      wadr => yt_rsc_3_9_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_3_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_3_0_i_clkr_en_d,
      d_d => yt_rsc_3_9_i_d_d,
      q_d => yt_rsc_3_9_i_q_d_1,
      radr_d => yt_rsc_3_9_i_radr_d,
      wadr_d => yt_rsc_3_9_i_wadr_d,
      we_d => yt_rsc_3_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_3_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_3_9_i_q <= yt_rsc_3_9_q;
  yt_rsc_3_9_radr <= yt_rsc_3_9_i_radr;
  yt_rsc_3_9_d <= yt_rsc_3_9_i_d;
  yt_rsc_3_9_wadr <= yt_rsc_3_9_i_wadr;
  yt_rsc_3_9_i_d_d <= yt_rsc_0_9_i_d_d_iff;
  yt_rsc_3_9_i_q_d <= yt_rsc_3_9_i_q_d_1;
  yt_rsc_3_9_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_3_9_i_wadr_d <= yt_rsc_0_2_i_wadr_d_iff;

  yt_rsc_3_10_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_113_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_3_10_clkr_en,
      clkw_en => yt_rsc_3_10_clkw_en,
      q => yt_rsc_3_10_i_q,
      radr => yt_rsc_3_10_i_radr,
      we => yt_rsc_3_10_we,
      d => yt_rsc_3_10_i_d,
      wadr => yt_rsc_3_10_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_3_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_3_0_i_clkr_en_d,
      d_d => yt_rsc_3_10_i_d_d,
      q_d => yt_rsc_3_10_i_q_d_1,
      radr_d => yt_rsc_3_10_i_radr_d,
      wadr_d => yt_rsc_3_10_i_wadr_d,
      we_d => yt_rsc_3_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_3_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_3_10_i_q <= yt_rsc_3_10_q;
  yt_rsc_3_10_radr <= yt_rsc_3_10_i_radr;
  yt_rsc_3_10_d <= yt_rsc_3_10_i_d;
  yt_rsc_3_10_wadr <= yt_rsc_3_10_i_wadr;
  yt_rsc_3_10_i_d_d <= yt_rsc_0_10_i_d_d_iff;
  yt_rsc_3_10_i_q_d <= yt_rsc_3_10_i_q_d_1;
  yt_rsc_3_10_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_3_10_i_wadr_d <= yt_rsc_0_10_i_wadr_d_iff;

  yt_rsc_3_11_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_114_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_3_11_clkr_en,
      clkw_en => yt_rsc_3_11_clkw_en,
      q => yt_rsc_3_11_i_q,
      radr => yt_rsc_3_11_i_radr,
      we => yt_rsc_3_11_we,
      d => yt_rsc_3_11_i_d,
      wadr => yt_rsc_3_11_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_3_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_3_0_i_clkr_en_d,
      d_d => yt_rsc_3_11_i_d_d,
      q_d => yt_rsc_3_11_i_q_d_1,
      radr_d => yt_rsc_3_11_i_radr_d,
      wadr_d => yt_rsc_3_11_i_wadr_d,
      we_d => yt_rsc_3_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_3_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_3_11_i_q <= yt_rsc_3_11_q;
  yt_rsc_3_11_radr <= yt_rsc_3_11_i_radr;
  yt_rsc_3_11_d <= yt_rsc_3_11_i_d;
  yt_rsc_3_11_wadr <= yt_rsc_3_11_i_wadr;
  yt_rsc_3_11_i_d_d <= yt_rsc_0_11_i_d_d_iff;
  yt_rsc_3_11_i_q_d <= yt_rsc_3_11_i_q_d_1;
  yt_rsc_3_11_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_3_11_i_wadr_d <= yt_rsc_0_11_i_wadr_d_iff;

  yt_rsc_3_12_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_115_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_3_12_clkr_en,
      clkw_en => yt_rsc_3_12_clkw_en,
      q => yt_rsc_3_12_i_q,
      radr => yt_rsc_3_12_i_radr,
      we => yt_rsc_3_12_we,
      d => yt_rsc_3_12_i_d,
      wadr => yt_rsc_3_12_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_3_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_3_0_i_clkr_en_d,
      d_d => yt_rsc_3_12_i_d_d,
      q_d => yt_rsc_3_12_i_q_d_1,
      radr_d => yt_rsc_3_12_i_radr_d,
      wadr_d => yt_rsc_3_12_i_wadr_d,
      we_d => yt_rsc_3_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_3_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_3_12_i_q <= yt_rsc_3_12_q;
  yt_rsc_3_12_radr <= yt_rsc_3_12_i_radr;
  yt_rsc_3_12_d <= yt_rsc_3_12_i_d;
  yt_rsc_3_12_wadr <= yt_rsc_3_12_i_wadr;
  yt_rsc_3_12_i_d_d <= yt_rsc_0_12_i_d_d_iff;
  yt_rsc_3_12_i_q_d <= yt_rsc_3_12_i_q_d_1;
  yt_rsc_3_12_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_3_12_i_wadr_d <= yt_rsc_0_3_i_wadr_d_iff;

  yt_rsc_3_13_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_116_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_3_13_clkr_en,
      clkw_en => yt_rsc_3_13_clkw_en,
      q => yt_rsc_3_13_i_q,
      radr => yt_rsc_3_13_i_radr,
      we => yt_rsc_3_13_we,
      d => yt_rsc_3_13_i_d,
      wadr => yt_rsc_3_13_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_3_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_3_0_i_clkr_en_d,
      d_d => yt_rsc_3_13_i_d_d,
      q_d => yt_rsc_3_13_i_q_d_1,
      radr_d => yt_rsc_3_13_i_radr_d,
      wadr_d => yt_rsc_3_13_i_wadr_d,
      we_d => yt_rsc_3_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_3_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_3_13_i_q <= yt_rsc_3_13_q;
  yt_rsc_3_13_radr <= yt_rsc_3_13_i_radr;
  yt_rsc_3_13_d <= yt_rsc_3_13_i_d;
  yt_rsc_3_13_wadr <= yt_rsc_3_13_i_wadr;
  yt_rsc_3_13_i_d_d <= yt_rsc_0_13_i_d_d_iff;
  yt_rsc_3_13_i_q_d <= yt_rsc_3_13_i_q_d_1;
  yt_rsc_3_13_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_3_13_i_wadr_d <= yt_rsc_0_4_i_wadr_d_iff;

  yt_rsc_3_14_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_117_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_3_14_clkr_en,
      clkw_en => yt_rsc_3_14_clkw_en,
      q => yt_rsc_3_14_i_q,
      radr => yt_rsc_3_14_i_radr,
      we => yt_rsc_3_14_we,
      d => yt_rsc_3_14_i_d,
      wadr => yt_rsc_3_14_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_3_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_3_0_i_clkr_en_d,
      d_d => yt_rsc_3_14_i_d_d,
      q_d => yt_rsc_3_14_i_q_d_1,
      radr_d => yt_rsc_3_14_i_radr_d,
      wadr_d => yt_rsc_3_14_i_wadr_d,
      we_d => yt_rsc_3_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_3_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_3_14_i_q <= yt_rsc_3_14_q;
  yt_rsc_3_14_radr <= yt_rsc_3_14_i_radr;
  yt_rsc_3_14_d <= yt_rsc_3_14_i_d;
  yt_rsc_3_14_wadr <= yt_rsc_3_14_i_wadr;
  yt_rsc_3_14_i_d_d <= yt_rsc_0_14_i_d_d_iff;
  yt_rsc_3_14_i_q_d <= yt_rsc_3_14_i_q_d_1;
  yt_rsc_3_14_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_3_14_i_wadr_d <= yt_rsc_0_5_i_wadr_d_iff;

  yt_rsc_3_15_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_118_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_3_15_clkr_en,
      clkw_en => yt_rsc_3_15_clkw_en,
      q => yt_rsc_3_15_i_q,
      radr => yt_rsc_3_15_i_radr,
      we => yt_rsc_3_15_we,
      d => yt_rsc_3_15_i_d,
      wadr => yt_rsc_3_15_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_3_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_3_0_i_clkr_en_d,
      d_d => yt_rsc_3_15_i_d_d,
      q_d => yt_rsc_3_15_i_q_d_1,
      radr_d => yt_rsc_3_15_i_radr_d,
      wadr_d => yt_rsc_3_15_i_wadr_d,
      we_d => yt_rsc_3_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_3_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_3_15_i_q <= yt_rsc_3_15_q;
  yt_rsc_3_15_radr <= yt_rsc_3_15_i_radr;
  yt_rsc_3_15_d <= yt_rsc_3_15_i_d;
  yt_rsc_3_15_wadr <= yt_rsc_3_15_i_wadr;
  yt_rsc_3_15_i_d_d <= yt_rsc_0_15_i_d_d_iff;
  yt_rsc_3_15_i_q_d <= yt_rsc_3_15_i_q_d_1;
  yt_rsc_3_15_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_3_15_i_wadr_d <= yt_rsc_0_6_i_wadr_d_iff;

  yt_rsc_3_16_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_119_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_3_16_clkr_en,
      clkw_en => yt_rsc_3_16_clkw_en,
      q => yt_rsc_3_16_i_q,
      radr => yt_rsc_3_16_i_radr,
      we => yt_rsc_3_16_we,
      d => yt_rsc_3_16_i_d,
      wadr => yt_rsc_3_16_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_3_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_3_16_i_clkr_en_d,
      d_d => yt_rsc_3_16_i_d_d,
      q_d => yt_rsc_3_16_i_q_d_1,
      radr_d => yt_rsc_3_16_i_radr_d,
      wadr_d => yt_rsc_3_16_i_wadr_d,
      we_d => yt_rsc_3_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_3_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_3_16_i_q <= yt_rsc_3_16_q;
  yt_rsc_3_16_radr <= yt_rsc_3_16_i_radr;
  yt_rsc_3_16_d <= yt_rsc_3_16_i_d;
  yt_rsc_3_16_wadr <= yt_rsc_3_16_i_wadr;
  yt_rsc_3_16_i_d_d <= yt_rsc_0_0_i_d_d_iff;
  yt_rsc_3_16_i_q_d <= yt_rsc_3_16_i_q_d_1;
  yt_rsc_3_16_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_3_16_i_wadr_d <= yt_rsc_0_0_i_wadr_d_iff;

  yt_rsc_3_17_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_120_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_3_17_clkr_en,
      clkw_en => yt_rsc_3_17_clkw_en,
      q => yt_rsc_3_17_i_q,
      radr => yt_rsc_3_17_i_radr,
      we => yt_rsc_3_17_we,
      d => yt_rsc_3_17_i_d,
      wadr => yt_rsc_3_17_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_3_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_3_16_i_clkr_en_d,
      d_d => yt_rsc_3_17_i_d_d,
      q_d => yt_rsc_3_17_i_q_d_1,
      radr_d => yt_rsc_3_17_i_radr_d,
      wadr_d => yt_rsc_3_17_i_wadr_d,
      we_d => yt_rsc_3_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_3_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_3_17_i_q <= yt_rsc_3_17_q;
  yt_rsc_3_17_radr <= yt_rsc_3_17_i_radr;
  yt_rsc_3_17_d <= yt_rsc_3_17_i_d;
  yt_rsc_3_17_wadr <= yt_rsc_3_17_i_wadr;
  yt_rsc_3_17_i_d_d <= yt_rsc_0_1_i_d_d_iff;
  yt_rsc_3_17_i_q_d <= yt_rsc_3_17_i_q_d_1;
  yt_rsc_3_17_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_3_17_i_wadr_d <= yt_rsc_0_1_i_wadr_d_iff;

  yt_rsc_3_18_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_121_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_3_18_clkr_en,
      clkw_en => yt_rsc_3_18_clkw_en,
      q => yt_rsc_3_18_i_q,
      radr => yt_rsc_3_18_i_radr,
      we => yt_rsc_3_18_we,
      d => yt_rsc_3_18_i_d,
      wadr => yt_rsc_3_18_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_3_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_3_16_i_clkr_en_d,
      d_d => yt_rsc_3_18_i_d_d,
      q_d => yt_rsc_3_18_i_q_d_1,
      radr_d => yt_rsc_3_18_i_radr_d,
      wadr_d => yt_rsc_3_18_i_wadr_d,
      we_d => yt_rsc_3_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_3_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_3_18_i_q <= yt_rsc_3_18_q;
  yt_rsc_3_18_radr <= yt_rsc_3_18_i_radr;
  yt_rsc_3_18_d <= yt_rsc_3_18_i_d;
  yt_rsc_3_18_wadr <= yt_rsc_3_18_i_wadr;
  yt_rsc_3_18_i_d_d <= yt_rsc_0_2_i_d_d_iff;
  yt_rsc_3_18_i_q_d <= yt_rsc_3_18_i_q_d_1;
  yt_rsc_3_18_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_3_18_i_wadr_d <= yt_rsc_0_2_i_wadr_d_iff;

  yt_rsc_3_19_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_122_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_3_19_clkr_en,
      clkw_en => yt_rsc_3_19_clkw_en,
      q => yt_rsc_3_19_i_q,
      radr => yt_rsc_3_19_i_radr,
      we => yt_rsc_3_19_we,
      d => yt_rsc_3_19_i_d,
      wadr => yt_rsc_3_19_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_3_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_3_16_i_clkr_en_d,
      d_d => yt_rsc_3_19_i_d_d,
      q_d => yt_rsc_3_19_i_q_d_1,
      radr_d => yt_rsc_3_19_i_radr_d,
      wadr_d => yt_rsc_3_19_i_wadr_d,
      we_d => yt_rsc_3_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_3_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_3_19_i_q <= yt_rsc_3_19_q;
  yt_rsc_3_19_radr <= yt_rsc_3_19_i_radr;
  yt_rsc_3_19_d <= yt_rsc_3_19_i_d;
  yt_rsc_3_19_wadr <= yt_rsc_3_19_i_wadr;
  yt_rsc_3_19_i_d_d <= yt_rsc_0_3_i_d_d_iff;
  yt_rsc_3_19_i_q_d <= yt_rsc_3_19_i_q_d_1;
  yt_rsc_3_19_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_3_19_i_wadr_d <= yt_rsc_0_3_i_wadr_d_iff;

  yt_rsc_3_20_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_123_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_3_20_clkr_en,
      clkw_en => yt_rsc_3_20_clkw_en,
      q => yt_rsc_3_20_i_q,
      radr => yt_rsc_3_20_i_radr,
      we => yt_rsc_3_20_we,
      d => yt_rsc_3_20_i_d,
      wadr => yt_rsc_3_20_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_3_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_3_16_i_clkr_en_d,
      d_d => yt_rsc_3_20_i_d_d,
      q_d => yt_rsc_3_20_i_q_d_1,
      radr_d => yt_rsc_3_20_i_radr_d,
      wadr_d => yt_rsc_3_20_i_wadr_d,
      we_d => yt_rsc_3_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_3_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_3_20_i_q <= yt_rsc_3_20_q;
  yt_rsc_3_20_radr <= yt_rsc_3_20_i_radr;
  yt_rsc_3_20_d <= yt_rsc_3_20_i_d;
  yt_rsc_3_20_wadr <= yt_rsc_3_20_i_wadr;
  yt_rsc_3_20_i_d_d <= yt_rsc_0_4_i_d_d_iff;
  yt_rsc_3_20_i_q_d <= yt_rsc_3_20_i_q_d_1;
  yt_rsc_3_20_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_3_20_i_wadr_d <= yt_rsc_0_4_i_wadr_d_iff;

  yt_rsc_3_21_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_124_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_3_21_clkr_en,
      clkw_en => yt_rsc_3_21_clkw_en,
      q => yt_rsc_3_21_i_q,
      radr => yt_rsc_3_21_i_radr,
      we => yt_rsc_3_21_we,
      d => yt_rsc_3_21_i_d,
      wadr => yt_rsc_3_21_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_3_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_3_16_i_clkr_en_d,
      d_d => yt_rsc_3_21_i_d_d,
      q_d => yt_rsc_3_21_i_q_d_1,
      radr_d => yt_rsc_3_21_i_radr_d,
      wadr_d => yt_rsc_3_21_i_wadr_d,
      we_d => yt_rsc_3_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_3_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_3_21_i_q <= yt_rsc_3_21_q;
  yt_rsc_3_21_radr <= yt_rsc_3_21_i_radr;
  yt_rsc_3_21_d <= yt_rsc_3_21_i_d;
  yt_rsc_3_21_wadr <= yt_rsc_3_21_i_wadr;
  yt_rsc_3_21_i_d_d <= yt_rsc_0_5_i_d_d_iff;
  yt_rsc_3_21_i_q_d <= yt_rsc_3_21_i_q_d_1;
  yt_rsc_3_21_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_3_21_i_wadr_d <= yt_rsc_0_5_i_wadr_d_iff;

  yt_rsc_3_22_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_125_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_3_22_clkr_en,
      clkw_en => yt_rsc_3_22_clkw_en,
      q => yt_rsc_3_22_i_q,
      radr => yt_rsc_3_22_i_radr,
      we => yt_rsc_3_22_we,
      d => yt_rsc_3_22_i_d,
      wadr => yt_rsc_3_22_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_3_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_3_16_i_clkr_en_d,
      d_d => yt_rsc_3_22_i_d_d,
      q_d => yt_rsc_3_22_i_q_d_1,
      radr_d => yt_rsc_3_22_i_radr_d,
      wadr_d => yt_rsc_3_22_i_wadr_d,
      we_d => yt_rsc_3_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_3_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_3_22_i_q <= yt_rsc_3_22_q;
  yt_rsc_3_22_radr <= yt_rsc_3_22_i_radr;
  yt_rsc_3_22_d <= yt_rsc_3_22_i_d;
  yt_rsc_3_22_wadr <= yt_rsc_3_22_i_wadr;
  yt_rsc_3_22_i_d_d <= yt_rsc_0_6_i_d_d_iff;
  yt_rsc_3_22_i_q_d <= yt_rsc_3_22_i_q_d_1;
  yt_rsc_3_22_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_3_22_i_wadr_d <= yt_rsc_0_6_i_wadr_d_iff;

  yt_rsc_3_23_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_126_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_3_23_clkr_en,
      clkw_en => yt_rsc_3_23_clkw_en,
      q => yt_rsc_3_23_i_q,
      radr => yt_rsc_3_23_i_radr,
      we => yt_rsc_3_23_we,
      d => yt_rsc_3_23_i_d,
      wadr => yt_rsc_3_23_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_3_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_3_16_i_clkr_en_d,
      d_d => yt_rsc_3_23_i_d_d,
      q_d => yt_rsc_3_23_i_q_d_1,
      radr_d => yt_rsc_3_23_i_radr_d,
      wadr_d => yt_rsc_3_23_i_wadr_d,
      we_d => yt_rsc_3_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_3_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_3_23_i_q <= yt_rsc_3_23_q;
  yt_rsc_3_23_radr <= yt_rsc_3_23_i_radr;
  yt_rsc_3_23_d <= yt_rsc_3_23_i_d;
  yt_rsc_3_23_wadr <= yt_rsc_3_23_i_wadr;
  yt_rsc_3_23_i_d_d <= yt_rsc_0_7_i_d_d_iff;
  yt_rsc_3_23_i_q_d <= yt_rsc_3_23_i_q_d_1;
  yt_rsc_3_23_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_3_23_i_wadr_d <= yt_rsc_0_0_i_wadr_d_iff;

  yt_rsc_3_24_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_127_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_3_24_clkr_en,
      clkw_en => yt_rsc_3_24_clkw_en,
      q => yt_rsc_3_24_i_q,
      radr => yt_rsc_3_24_i_radr,
      we => yt_rsc_3_24_we,
      d => yt_rsc_3_24_i_d,
      wadr => yt_rsc_3_24_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_3_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_3_16_i_clkr_en_d,
      d_d => yt_rsc_3_24_i_d_d,
      q_d => yt_rsc_3_24_i_q_d_1,
      radr_d => yt_rsc_3_24_i_radr_d,
      wadr_d => yt_rsc_3_24_i_wadr_d,
      we_d => yt_rsc_3_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_3_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_3_24_i_q <= yt_rsc_3_24_q;
  yt_rsc_3_24_radr <= yt_rsc_3_24_i_radr;
  yt_rsc_3_24_d <= yt_rsc_3_24_i_d;
  yt_rsc_3_24_wadr <= yt_rsc_3_24_i_wadr;
  yt_rsc_3_24_i_d_d <= yt_rsc_0_8_i_d_d_iff;
  yt_rsc_3_24_i_q_d <= yt_rsc_3_24_i_q_d_1;
  yt_rsc_3_24_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_3_24_i_wadr_d <= yt_rsc_0_1_i_wadr_d_iff;

  yt_rsc_3_25_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_128_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_3_25_clkr_en,
      clkw_en => yt_rsc_3_25_clkw_en,
      q => yt_rsc_3_25_i_q,
      radr => yt_rsc_3_25_i_radr,
      we => yt_rsc_3_25_we,
      d => yt_rsc_3_25_i_d,
      wadr => yt_rsc_3_25_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_3_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_3_16_i_clkr_en_d,
      d_d => yt_rsc_3_25_i_d_d,
      q_d => yt_rsc_3_25_i_q_d_1,
      radr_d => yt_rsc_3_25_i_radr_d,
      wadr_d => yt_rsc_3_25_i_wadr_d,
      we_d => yt_rsc_3_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_3_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_3_25_i_q <= yt_rsc_3_25_q;
  yt_rsc_3_25_radr <= yt_rsc_3_25_i_radr;
  yt_rsc_3_25_d <= yt_rsc_3_25_i_d;
  yt_rsc_3_25_wadr <= yt_rsc_3_25_i_wadr;
  yt_rsc_3_25_i_d_d <= yt_rsc_0_9_i_d_d_iff;
  yt_rsc_3_25_i_q_d <= yt_rsc_3_25_i_q_d_1;
  yt_rsc_3_25_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_3_25_i_wadr_d <= yt_rsc_0_2_i_wadr_d_iff;

  yt_rsc_3_26_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_129_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_3_26_clkr_en,
      clkw_en => yt_rsc_3_26_clkw_en,
      q => yt_rsc_3_26_i_q,
      radr => yt_rsc_3_26_i_radr,
      we => yt_rsc_3_26_we,
      d => yt_rsc_3_26_i_d,
      wadr => yt_rsc_3_26_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_3_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_3_16_i_clkr_en_d,
      d_d => yt_rsc_3_26_i_d_d,
      q_d => yt_rsc_3_26_i_q_d_1,
      radr_d => yt_rsc_3_26_i_radr_d,
      wadr_d => yt_rsc_3_26_i_wadr_d,
      we_d => yt_rsc_3_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_3_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_3_26_i_q <= yt_rsc_3_26_q;
  yt_rsc_3_26_radr <= yt_rsc_3_26_i_radr;
  yt_rsc_3_26_d <= yt_rsc_3_26_i_d;
  yt_rsc_3_26_wadr <= yt_rsc_3_26_i_wadr;
  yt_rsc_3_26_i_d_d <= yt_rsc_0_10_i_d_d_iff;
  yt_rsc_3_26_i_q_d <= yt_rsc_3_26_i_q_d_1;
  yt_rsc_3_26_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_3_26_i_wadr_d <= yt_rsc_0_10_i_wadr_d_iff;

  yt_rsc_3_27_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_130_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_3_27_clkr_en,
      clkw_en => yt_rsc_3_27_clkw_en,
      q => yt_rsc_3_27_i_q,
      radr => yt_rsc_3_27_i_radr,
      we => yt_rsc_3_27_we,
      d => yt_rsc_3_27_i_d,
      wadr => yt_rsc_3_27_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_3_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_3_16_i_clkr_en_d,
      d_d => yt_rsc_3_27_i_d_d,
      q_d => yt_rsc_3_27_i_q_d_1,
      radr_d => yt_rsc_3_27_i_radr_d,
      wadr_d => yt_rsc_3_27_i_wadr_d,
      we_d => yt_rsc_3_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_3_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_3_27_i_q <= yt_rsc_3_27_q;
  yt_rsc_3_27_radr <= yt_rsc_3_27_i_radr;
  yt_rsc_3_27_d <= yt_rsc_3_27_i_d;
  yt_rsc_3_27_wadr <= yt_rsc_3_27_i_wadr;
  yt_rsc_3_27_i_d_d <= yt_rsc_0_11_i_d_d_iff;
  yt_rsc_3_27_i_q_d <= yt_rsc_3_27_i_q_d_1;
  yt_rsc_3_27_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_3_27_i_wadr_d <= yt_rsc_0_11_i_wadr_d_iff;

  yt_rsc_3_28_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_131_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_3_28_clkr_en,
      clkw_en => yt_rsc_3_28_clkw_en,
      q => yt_rsc_3_28_i_q,
      radr => yt_rsc_3_28_i_radr,
      we => yt_rsc_3_28_we,
      d => yt_rsc_3_28_i_d,
      wadr => yt_rsc_3_28_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_3_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_3_16_i_clkr_en_d,
      d_d => yt_rsc_3_28_i_d_d,
      q_d => yt_rsc_3_28_i_q_d_1,
      radr_d => yt_rsc_3_28_i_radr_d,
      wadr_d => yt_rsc_3_28_i_wadr_d,
      we_d => yt_rsc_3_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_3_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_3_28_i_q <= yt_rsc_3_28_q;
  yt_rsc_3_28_radr <= yt_rsc_3_28_i_radr;
  yt_rsc_3_28_d <= yt_rsc_3_28_i_d;
  yt_rsc_3_28_wadr <= yt_rsc_3_28_i_wadr;
  yt_rsc_3_28_i_d_d <= yt_rsc_0_12_i_d_d_iff;
  yt_rsc_3_28_i_q_d <= yt_rsc_3_28_i_q_d_1;
  yt_rsc_3_28_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_3_28_i_wadr_d <= yt_rsc_0_3_i_wadr_d_iff;

  yt_rsc_3_29_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_132_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_3_29_clkr_en,
      clkw_en => yt_rsc_3_29_clkw_en,
      q => yt_rsc_3_29_i_q,
      radr => yt_rsc_3_29_i_radr,
      we => yt_rsc_3_29_we,
      d => yt_rsc_3_29_i_d,
      wadr => yt_rsc_3_29_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_3_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_3_16_i_clkr_en_d,
      d_d => yt_rsc_3_29_i_d_d,
      q_d => yt_rsc_3_29_i_q_d_1,
      radr_d => yt_rsc_3_29_i_radr_d,
      wadr_d => yt_rsc_3_29_i_wadr_d,
      we_d => yt_rsc_3_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_3_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_3_29_i_q <= yt_rsc_3_29_q;
  yt_rsc_3_29_radr <= yt_rsc_3_29_i_radr;
  yt_rsc_3_29_d <= yt_rsc_3_29_i_d;
  yt_rsc_3_29_wadr <= yt_rsc_3_29_i_wadr;
  yt_rsc_3_29_i_d_d <= yt_rsc_0_13_i_d_d_iff;
  yt_rsc_3_29_i_q_d <= yt_rsc_3_29_i_q_d_1;
  yt_rsc_3_29_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_3_29_i_wadr_d <= yt_rsc_0_4_i_wadr_d_iff;

  yt_rsc_3_30_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_133_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_3_30_clkr_en,
      clkw_en => yt_rsc_3_30_clkw_en,
      q => yt_rsc_3_30_i_q,
      radr => yt_rsc_3_30_i_radr,
      we => yt_rsc_3_30_we,
      d => yt_rsc_3_30_i_d,
      wadr => yt_rsc_3_30_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_3_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_3_16_i_clkr_en_d,
      d_d => yt_rsc_3_30_i_d_d,
      q_d => yt_rsc_3_30_i_q_d_1,
      radr_d => yt_rsc_3_30_i_radr_d,
      wadr_d => yt_rsc_3_30_i_wadr_d,
      we_d => yt_rsc_3_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_3_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_3_30_i_q <= yt_rsc_3_30_q;
  yt_rsc_3_30_radr <= yt_rsc_3_30_i_radr;
  yt_rsc_3_30_d <= yt_rsc_3_30_i_d;
  yt_rsc_3_30_wadr <= yt_rsc_3_30_i_wadr;
  yt_rsc_3_30_i_d_d <= yt_rsc_0_14_i_d_d_iff;
  yt_rsc_3_30_i_q_d <= yt_rsc_3_30_i_q_d_1;
  yt_rsc_3_30_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_3_30_i_wadr_d <= yt_rsc_0_5_i_wadr_d_iff;

  yt_rsc_3_31_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_134_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_3_31_clkr_en,
      clkw_en => yt_rsc_3_31_clkw_en,
      q => yt_rsc_3_31_i_q,
      radr => yt_rsc_3_31_i_radr,
      we => yt_rsc_3_31_we,
      d => yt_rsc_3_31_i_d,
      wadr => yt_rsc_3_31_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_3_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_3_16_i_clkr_en_d,
      d_d => yt_rsc_3_31_i_d_d,
      q_d => yt_rsc_3_31_i_q_d_1,
      radr_d => yt_rsc_3_31_i_radr_d,
      wadr_d => yt_rsc_3_31_i_wadr_d,
      we_d => yt_rsc_3_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_3_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_3_31_i_q <= yt_rsc_3_31_q;
  yt_rsc_3_31_radr <= yt_rsc_3_31_i_radr;
  yt_rsc_3_31_d <= yt_rsc_3_31_i_d;
  yt_rsc_3_31_wadr <= yt_rsc_3_31_i_wadr;
  yt_rsc_3_31_i_d_d <= yt_rsc_0_15_i_d_d_iff;
  yt_rsc_3_31_i_q_d <= yt_rsc_3_31_i_q_d_1;
  yt_rsc_3_31_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_3_31_i_wadr_d <= yt_rsc_0_6_i_wadr_d_iff;

  yt_rsc_4_0_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_135_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_4_0_clkr_en,
      clkw_en => yt_rsc_4_0_clkw_en,
      q => yt_rsc_4_0_i_q,
      radr => yt_rsc_4_0_i_radr,
      we => yt_rsc_4_0_we,
      d => yt_rsc_4_0_i_d,
      wadr => yt_rsc_4_0_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_4_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_4_0_i_clkr_en_d,
      d_d => yt_rsc_4_0_i_d_d,
      q_d => yt_rsc_4_0_i_q_d_1,
      radr_d => yt_rsc_4_0_i_radr_d,
      wadr_d => yt_rsc_4_0_i_wadr_d,
      we_d => yt_rsc_4_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_4_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_4_0_i_q <= yt_rsc_4_0_q;
  yt_rsc_4_0_radr <= yt_rsc_4_0_i_radr;
  yt_rsc_4_0_d <= yt_rsc_4_0_i_d;
  yt_rsc_4_0_wadr <= yt_rsc_4_0_i_wadr;
  yt_rsc_4_0_i_d_d <= yt_rsc_4_0_i_d_d_iff;
  yt_rsc_4_0_i_q_d <= yt_rsc_4_0_i_q_d_1;
  yt_rsc_4_0_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_4_0_i_wadr_d <= yt_rsc_4_0_i_wadr_d_iff;

  yt_rsc_4_1_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_136_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_4_1_clkr_en,
      clkw_en => yt_rsc_4_1_clkw_en,
      q => yt_rsc_4_1_i_q,
      radr => yt_rsc_4_1_i_radr,
      we => yt_rsc_4_1_we,
      d => yt_rsc_4_1_i_d,
      wadr => yt_rsc_4_1_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_4_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_4_0_i_clkr_en_d,
      d_d => yt_rsc_4_1_i_d_d,
      q_d => yt_rsc_4_1_i_q_d_1,
      radr_d => yt_rsc_4_1_i_radr_d,
      wadr_d => yt_rsc_4_1_i_wadr_d,
      we_d => yt_rsc_4_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_4_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_4_1_i_q <= yt_rsc_4_1_q;
  yt_rsc_4_1_radr <= yt_rsc_4_1_i_radr;
  yt_rsc_4_1_d <= yt_rsc_4_1_i_d;
  yt_rsc_4_1_wadr <= yt_rsc_4_1_i_wadr;
  yt_rsc_4_1_i_d_d <= yt_rsc_4_1_i_d_d_iff;
  yt_rsc_4_1_i_q_d <= yt_rsc_4_1_i_q_d_1;
  yt_rsc_4_1_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_4_1_i_wadr_d <= yt_rsc_4_1_i_wadr_d_iff;

  yt_rsc_4_2_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_137_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_4_2_clkr_en,
      clkw_en => yt_rsc_4_2_clkw_en,
      q => yt_rsc_4_2_i_q,
      radr => yt_rsc_4_2_i_radr,
      we => yt_rsc_4_2_we,
      d => yt_rsc_4_2_i_d,
      wadr => yt_rsc_4_2_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_4_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_4_0_i_clkr_en_d,
      d_d => yt_rsc_4_2_i_d_d,
      q_d => yt_rsc_4_2_i_q_d_1,
      radr_d => yt_rsc_4_2_i_radr_d,
      wadr_d => yt_rsc_4_2_i_wadr_d,
      we_d => yt_rsc_4_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_4_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_4_2_i_q <= yt_rsc_4_2_q;
  yt_rsc_4_2_radr <= yt_rsc_4_2_i_radr;
  yt_rsc_4_2_d <= yt_rsc_4_2_i_d;
  yt_rsc_4_2_wadr <= yt_rsc_4_2_i_wadr;
  yt_rsc_4_2_i_d_d <= yt_rsc_4_2_i_d_d_iff;
  yt_rsc_4_2_i_q_d <= yt_rsc_4_2_i_q_d_1;
  yt_rsc_4_2_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_4_2_i_wadr_d <= yt_rsc_4_2_i_wadr_d_iff;

  yt_rsc_4_3_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_138_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_4_3_clkr_en,
      clkw_en => yt_rsc_4_3_clkw_en,
      q => yt_rsc_4_3_i_q,
      radr => yt_rsc_4_3_i_radr,
      we => yt_rsc_4_3_we,
      d => yt_rsc_4_3_i_d,
      wadr => yt_rsc_4_3_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_4_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_4_0_i_clkr_en_d,
      d_d => yt_rsc_4_3_i_d_d,
      q_d => yt_rsc_4_3_i_q_d_1,
      radr_d => yt_rsc_4_3_i_radr_d,
      wadr_d => yt_rsc_4_3_i_wadr_d,
      we_d => yt_rsc_4_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_4_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_4_3_i_q <= yt_rsc_4_3_q;
  yt_rsc_4_3_radr <= yt_rsc_4_3_i_radr;
  yt_rsc_4_3_d <= yt_rsc_4_3_i_d;
  yt_rsc_4_3_wadr <= yt_rsc_4_3_i_wadr;
  yt_rsc_4_3_i_d_d <= yt_rsc_4_3_i_d_d_iff;
  yt_rsc_4_3_i_q_d <= yt_rsc_4_3_i_q_d_1;
  yt_rsc_4_3_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_4_3_i_wadr_d <= yt_rsc_4_3_i_wadr_d_iff;

  yt_rsc_4_4_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_139_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_4_4_clkr_en,
      clkw_en => yt_rsc_4_4_clkw_en,
      q => yt_rsc_4_4_i_q,
      radr => yt_rsc_4_4_i_radr,
      we => yt_rsc_4_4_we,
      d => yt_rsc_4_4_i_d,
      wadr => yt_rsc_4_4_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_4_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_4_0_i_clkr_en_d,
      d_d => yt_rsc_4_4_i_d_d,
      q_d => yt_rsc_4_4_i_q_d_1,
      radr_d => yt_rsc_4_4_i_radr_d,
      wadr_d => yt_rsc_4_4_i_wadr_d,
      we_d => yt_rsc_4_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_4_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_4_4_i_q <= yt_rsc_4_4_q;
  yt_rsc_4_4_radr <= yt_rsc_4_4_i_radr;
  yt_rsc_4_4_d <= yt_rsc_4_4_i_d;
  yt_rsc_4_4_wadr <= yt_rsc_4_4_i_wadr;
  yt_rsc_4_4_i_d_d <= yt_rsc_4_4_i_d_d_iff;
  yt_rsc_4_4_i_q_d <= yt_rsc_4_4_i_q_d_1;
  yt_rsc_4_4_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_4_4_i_wadr_d <= yt_rsc_4_4_i_wadr_d_iff;

  yt_rsc_4_5_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_140_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_4_5_clkr_en,
      clkw_en => yt_rsc_4_5_clkw_en,
      q => yt_rsc_4_5_i_q,
      radr => yt_rsc_4_5_i_radr,
      we => yt_rsc_4_5_we,
      d => yt_rsc_4_5_i_d,
      wadr => yt_rsc_4_5_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_4_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_4_0_i_clkr_en_d,
      d_d => yt_rsc_4_5_i_d_d,
      q_d => yt_rsc_4_5_i_q_d_1,
      radr_d => yt_rsc_4_5_i_radr_d,
      wadr_d => yt_rsc_4_5_i_wadr_d,
      we_d => yt_rsc_4_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_4_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_4_5_i_q <= yt_rsc_4_5_q;
  yt_rsc_4_5_radr <= yt_rsc_4_5_i_radr;
  yt_rsc_4_5_d <= yt_rsc_4_5_i_d;
  yt_rsc_4_5_wadr <= yt_rsc_4_5_i_wadr;
  yt_rsc_4_5_i_d_d <= yt_rsc_4_5_i_d_d_iff;
  yt_rsc_4_5_i_q_d <= yt_rsc_4_5_i_q_d_1;
  yt_rsc_4_5_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_4_5_i_wadr_d <= yt_rsc_4_5_i_wadr_d_iff;

  yt_rsc_4_6_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_141_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_4_6_clkr_en,
      clkw_en => yt_rsc_4_6_clkw_en,
      q => yt_rsc_4_6_i_q,
      radr => yt_rsc_4_6_i_radr,
      we => yt_rsc_4_6_we,
      d => yt_rsc_4_6_i_d,
      wadr => yt_rsc_4_6_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_4_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_4_0_i_clkr_en_d,
      d_d => yt_rsc_4_6_i_d_d,
      q_d => yt_rsc_4_6_i_q_d_1,
      radr_d => yt_rsc_4_6_i_radr_d,
      wadr_d => yt_rsc_4_6_i_wadr_d,
      we_d => yt_rsc_4_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_4_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_4_6_i_q <= yt_rsc_4_6_q;
  yt_rsc_4_6_radr <= yt_rsc_4_6_i_radr;
  yt_rsc_4_6_d <= yt_rsc_4_6_i_d;
  yt_rsc_4_6_wadr <= yt_rsc_4_6_i_wadr;
  yt_rsc_4_6_i_d_d <= yt_rsc_4_6_i_d_d_iff;
  yt_rsc_4_6_i_q_d <= yt_rsc_4_6_i_q_d_1;
  yt_rsc_4_6_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_4_6_i_wadr_d <= yt_rsc_4_6_i_wadr_d_iff;

  yt_rsc_4_7_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_142_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_4_7_clkr_en,
      clkw_en => yt_rsc_4_7_clkw_en,
      q => yt_rsc_4_7_i_q,
      radr => yt_rsc_4_7_i_radr,
      we => yt_rsc_4_7_we,
      d => yt_rsc_4_7_i_d,
      wadr => yt_rsc_4_7_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_4_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_4_0_i_clkr_en_d,
      d_d => yt_rsc_4_7_i_d_d,
      q_d => yt_rsc_4_7_i_q_d_1,
      radr_d => yt_rsc_4_7_i_radr_d,
      wadr_d => yt_rsc_4_7_i_wadr_d,
      we_d => yt_rsc_4_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_4_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_4_7_i_q <= yt_rsc_4_7_q;
  yt_rsc_4_7_radr <= yt_rsc_4_7_i_radr;
  yt_rsc_4_7_d <= yt_rsc_4_7_i_d;
  yt_rsc_4_7_wadr <= yt_rsc_4_7_i_wadr;
  yt_rsc_4_7_i_d_d <= yt_rsc_4_7_i_d_d_iff;
  yt_rsc_4_7_i_q_d <= yt_rsc_4_7_i_q_d_1;
  yt_rsc_4_7_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_4_7_i_wadr_d <= yt_rsc_4_0_i_wadr_d_iff;

  yt_rsc_4_8_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_143_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_4_8_clkr_en,
      clkw_en => yt_rsc_4_8_clkw_en,
      q => yt_rsc_4_8_i_q,
      radr => yt_rsc_4_8_i_radr,
      we => yt_rsc_4_8_we,
      d => yt_rsc_4_8_i_d,
      wadr => yt_rsc_4_8_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_4_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_4_0_i_clkr_en_d,
      d_d => yt_rsc_4_8_i_d_d,
      q_d => yt_rsc_4_8_i_q_d_1,
      radr_d => yt_rsc_4_8_i_radr_d,
      wadr_d => yt_rsc_4_8_i_wadr_d,
      we_d => yt_rsc_4_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_4_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_4_8_i_q <= yt_rsc_4_8_q;
  yt_rsc_4_8_radr <= yt_rsc_4_8_i_radr;
  yt_rsc_4_8_d <= yt_rsc_4_8_i_d;
  yt_rsc_4_8_wadr <= yt_rsc_4_8_i_wadr;
  yt_rsc_4_8_i_d_d <= yt_rsc_4_8_i_d_d_iff;
  yt_rsc_4_8_i_q_d <= yt_rsc_4_8_i_q_d_1;
  yt_rsc_4_8_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_4_8_i_wadr_d <= yt_rsc_4_1_i_wadr_d_iff;

  yt_rsc_4_9_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_144_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_4_9_clkr_en,
      clkw_en => yt_rsc_4_9_clkw_en,
      q => yt_rsc_4_9_i_q,
      radr => yt_rsc_4_9_i_radr,
      we => yt_rsc_4_9_we,
      d => yt_rsc_4_9_i_d,
      wadr => yt_rsc_4_9_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_4_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_4_0_i_clkr_en_d,
      d_d => yt_rsc_4_9_i_d_d,
      q_d => yt_rsc_4_9_i_q_d_1,
      radr_d => yt_rsc_4_9_i_radr_d,
      wadr_d => yt_rsc_4_9_i_wadr_d,
      we_d => yt_rsc_4_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_4_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_4_9_i_q <= yt_rsc_4_9_q;
  yt_rsc_4_9_radr <= yt_rsc_4_9_i_radr;
  yt_rsc_4_9_d <= yt_rsc_4_9_i_d;
  yt_rsc_4_9_wadr <= yt_rsc_4_9_i_wadr;
  yt_rsc_4_9_i_d_d <= yt_rsc_4_9_i_d_d_iff;
  yt_rsc_4_9_i_q_d <= yt_rsc_4_9_i_q_d_1;
  yt_rsc_4_9_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_4_9_i_wadr_d <= yt_rsc_4_9_i_wadr_d_iff;

  yt_rsc_4_10_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_145_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_4_10_clkr_en,
      clkw_en => yt_rsc_4_10_clkw_en,
      q => yt_rsc_4_10_i_q,
      radr => yt_rsc_4_10_i_radr,
      we => yt_rsc_4_10_we,
      d => yt_rsc_4_10_i_d,
      wadr => yt_rsc_4_10_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_4_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_4_0_i_clkr_en_d,
      d_d => yt_rsc_4_10_i_d_d,
      q_d => yt_rsc_4_10_i_q_d_1,
      radr_d => yt_rsc_4_10_i_radr_d,
      wadr_d => yt_rsc_4_10_i_wadr_d,
      we_d => yt_rsc_4_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_4_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_4_10_i_q <= yt_rsc_4_10_q;
  yt_rsc_4_10_radr <= yt_rsc_4_10_i_radr;
  yt_rsc_4_10_d <= yt_rsc_4_10_i_d;
  yt_rsc_4_10_wadr <= yt_rsc_4_10_i_wadr;
  yt_rsc_4_10_i_d_d <= yt_rsc_4_10_i_d_d_iff;
  yt_rsc_4_10_i_q_d <= yt_rsc_4_10_i_q_d_1;
  yt_rsc_4_10_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_4_10_i_wadr_d <= yt_rsc_4_10_i_wadr_d_iff;

  yt_rsc_4_11_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_146_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_4_11_clkr_en,
      clkw_en => yt_rsc_4_11_clkw_en,
      q => yt_rsc_4_11_i_q,
      radr => yt_rsc_4_11_i_radr,
      we => yt_rsc_4_11_we,
      d => yt_rsc_4_11_i_d,
      wadr => yt_rsc_4_11_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_4_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_4_0_i_clkr_en_d,
      d_d => yt_rsc_4_11_i_d_d,
      q_d => yt_rsc_4_11_i_q_d_1,
      radr_d => yt_rsc_4_11_i_radr_d,
      wadr_d => yt_rsc_4_11_i_wadr_d,
      we_d => yt_rsc_4_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_4_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_4_11_i_q <= yt_rsc_4_11_q;
  yt_rsc_4_11_radr <= yt_rsc_4_11_i_radr;
  yt_rsc_4_11_d <= yt_rsc_4_11_i_d;
  yt_rsc_4_11_wadr <= yt_rsc_4_11_i_wadr;
  yt_rsc_4_11_i_d_d <= yt_rsc_4_11_i_d_d_iff;
  yt_rsc_4_11_i_q_d <= yt_rsc_4_11_i_q_d_1;
  yt_rsc_4_11_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_4_11_i_wadr_d <= yt_rsc_4_11_i_wadr_d_iff;

  yt_rsc_4_12_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_147_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_4_12_clkr_en,
      clkw_en => yt_rsc_4_12_clkw_en,
      q => yt_rsc_4_12_i_q,
      radr => yt_rsc_4_12_i_radr,
      we => yt_rsc_4_12_we,
      d => yt_rsc_4_12_i_d,
      wadr => yt_rsc_4_12_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_4_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_4_0_i_clkr_en_d,
      d_d => yt_rsc_4_12_i_d_d,
      q_d => yt_rsc_4_12_i_q_d_1,
      radr_d => yt_rsc_4_12_i_radr_d,
      wadr_d => yt_rsc_4_12_i_wadr_d,
      we_d => yt_rsc_4_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_4_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_4_12_i_q <= yt_rsc_4_12_q;
  yt_rsc_4_12_radr <= yt_rsc_4_12_i_radr;
  yt_rsc_4_12_d <= yt_rsc_4_12_i_d;
  yt_rsc_4_12_wadr <= yt_rsc_4_12_i_wadr;
  yt_rsc_4_12_i_d_d <= yt_rsc_4_12_i_d_d_iff;
  yt_rsc_4_12_i_q_d <= yt_rsc_4_12_i_q_d_1;
  yt_rsc_4_12_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_4_12_i_wadr_d <= yt_rsc_4_3_i_wadr_d_iff;

  yt_rsc_4_13_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_148_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_4_13_clkr_en,
      clkw_en => yt_rsc_4_13_clkw_en,
      q => yt_rsc_4_13_i_q,
      radr => yt_rsc_4_13_i_radr,
      we => yt_rsc_4_13_we,
      d => yt_rsc_4_13_i_d,
      wadr => yt_rsc_4_13_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_4_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_4_0_i_clkr_en_d,
      d_d => yt_rsc_4_13_i_d_d,
      q_d => yt_rsc_4_13_i_q_d_1,
      radr_d => yt_rsc_4_13_i_radr_d,
      wadr_d => yt_rsc_4_13_i_wadr_d,
      we_d => yt_rsc_4_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_4_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_4_13_i_q <= yt_rsc_4_13_q;
  yt_rsc_4_13_radr <= yt_rsc_4_13_i_radr;
  yt_rsc_4_13_d <= yt_rsc_4_13_i_d;
  yt_rsc_4_13_wadr <= yt_rsc_4_13_i_wadr;
  yt_rsc_4_13_i_d_d <= yt_rsc_4_13_i_d_d_iff;
  yt_rsc_4_13_i_q_d <= yt_rsc_4_13_i_q_d_1;
  yt_rsc_4_13_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_4_13_i_wadr_d <= yt_rsc_4_4_i_wadr_d_iff;

  yt_rsc_4_14_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_149_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_4_14_clkr_en,
      clkw_en => yt_rsc_4_14_clkw_en,
      q => yt_rsc_4_14_i_q,
      radr => yt_rsc_4_14_i_radr,
      we => yt_rsc_4_14_we,
      d => yt_rsc_4_14_i_d,
      wadr => yt_rsc_4_14_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_4_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_4_0_i_clkr_en_d,
      d_d => yt_rsc_4_14_i_d_d,
      q_d => yt_rsc_4_14_i_q_d_1,
      radr_d => yt_rsc_4_14_i_radr_d,
      wadr_d => yt_rsc_4_14_i_wadr_d,
      we_d => yt_rsc_4_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_4_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_4_14_i_q <= yt_rsc_4_14_q;
  yt_rsc_4_14_radr <= yt_rsc_4_14_i_radr;
  yt_rsc_4_14_d <= yt_rsc_4_14_i_d;
  yt_rsc_4_14_wadr <= yt_rsc_4_14_i_wadr;
  yt_rsc_4_14_i_d_d <= yt_rsc_4_14_i_d_d_iff;
  yt_rsc_4_14_i_q_d <= yt_rsc_4_14_i_q_d_1;
  yt_rsc_4_14_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_4_14_i_wadr_d <= yt_rsc_4_5_i_wadr_d_iff;

  yt_rsc_4_15_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_150_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_4_15_clkr_en,
      clkw_en => yt_rsc_4_15_clkw_en,
      q => yt_rsc_4_15_i_q,
      radr => yt_rsc_4_15_i_radr,
      we => yt_rsc_4_15_we,
      d => yt_rsc_4_15_i_d,
      wadr => yt_rsc_4_15_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_4_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_4_0_i_clkr_en_d,
      d_d => yt_rsc_4_15_i_d_d,
      q_d => yt_rsc_4_15_i_q_d_1,
      radr_d => yt_rsc_4_15_i_radr_d,
      wadr_d => yt_rsc_4_15_i_wadr_d,
      we_d => yt_rsc_4_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_4_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_4_15_i_q <= yt_rsc_4_15_q;
  yt_rsc_4_15_radr <= yt_rsc_4_15_i_radr;
  yt_rsc_4_15_d <= yt_rsc_4_15_i_d;
  yt_rsc_4_15_wadr <= yt_rsc_4_15_i_wadr;
  yt_rsc_4_15_i_d_d <= yt_rsc_4_15_i_d_d_iff;
  yt_rsc_4_15_i_q_d <= yt_rsc_4_15_i_q_d_1;
  yt_rsc_4_15_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_4_15_i_wadr_d <= yt_rsc_4_6_i_wadr_d_iff;

  yt_rsc_4_16_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_151_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_4_16_clkr_en,
      clkw_en => yt_rsc_4_16_clkw_en,
      q => yt_rsc_4_16_i_q,
      radr => yt_rsc_4_16_i_radr,
      we => yt_rsc_4_16_we,
      d => yt_rsc_4_16_i_d,
      wadr => yt_rsc_4_16_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_4_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_4_16_i_clkr_en_d,
      d_d => yt_rsc_4_16_i_d_d,
      q_d => yt_rsc_4_16_i_q_d_1,
      radr_d => yt_rsc_4_16_i_radr_d,
      wadr_d => yt_rsc_4_16_i_wadr_d,
      we_d => yt_rsc_4_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_4_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_4_16_i_q <= yt_rsc_4_16_q;
  yt_rsc_4_16_radr <= yt_rsc_4_16_i_radr;
  yt_rsc_4_16_d <= yt_rsc_4_16_i_d;
  yt_rsc_4_16_wadr <= yt_rsc_4_16_i_wadr;
  yt_rsc_4_16_i_d_d <= yt_rsc_4_0_i_d_d_iff;
  yt_rsc_4_16_i_q_d <= yt_rsc_4_16_i_q_d_1;
  yt_rsc_4_16_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_4_16_i_wadr_d <= yt_rsc_4_0_i_wadr_d_iff;

  yt_rsc_4_17_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_152_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_4_17_clkr_en,
      clkw_en => yt_rsc_4_17_clkw_en,
      q => yt_rsc_4_17_i_q,
      radr => yt_rsc_4_17_i_radr,
      we => yt_rsc_4_17_we,
      d => yt_rsc_4_17_i_d,
      wadr => yt_rsc_4_17_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_4_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_4_16_i_clkr_en_d,
      d_d => yt_rsc_4_17_i_d_d,
      q_d => yt_rsc_4_17_i_q_d_1,
      radr_d => yt_rsc_4_17_i_radr_d,
      wadr_d => yt_rsc_4_17_i_wadr_d,
      we_d => yt_rsc_4_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_4_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_4_17_i_q <= yt_rsc_4_17_q;
  yt_rsc_4_17_radr <= yt_rsc_4_17_i_radr;
  yt_rsc_4_17_d <= yt_rsc_4_17_i_d;
  yt_rsc_4_17_wadr <= yt_rsc_4_17_i_wadr;
  yt_rsc_4_17_i_d_d <= yt_rsc_4_1_i_d_d_iff;
  yt_rsc_4_17_i_q_d <= yt_rsc_4_17_i_q_d_1;
  yt_rsc_4_17_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_4_17_i_wadr_d <= yt_rsc_4_1_i_wadr_d_iff;

  yt_rsc_4_18_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_153_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_4_18_clkr_en,
      clkw_en => yt_rsc_4_18_clkw_en,
      q => yt_rsc_4_18_i_q,
      radr => yt_rsc_4_18_i_radr,
      we => yt_rsc_4_18_we,
      d => yt_rsc_4_18_i_d,
      wadr => yt_rsc_4_18_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_4_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_4_16_i_clkr_en_d,
      d_d => yt_rsc_4_18_i_d_d,
      q_d => yt_rsc_4_18_i_q_d_1,
      radr_d => yt_rsc_4_18_i_radr_d,
      wadr_d => yt_rsc_4_18_i_wadr_d,
      we_d => yt_rsc_4_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_4_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_4_18_i_q <= yt_rsc_4_18_q;
  yt_rsc_4_18_radr <= yt_rsc_4_18_i_radr;
  yt_rsc_4_18_d <= yt_rsc_4_18_i_d;
  yt_rsc_4_18_wadr <= yt_rsc_4_18_i_wadr;
  yt_rsc_4_18_i_d_d <= yt_rsc_4_2_i_d_d_iff;
  yt_rsc_4_18_i_q_d <= yt_rsc_4_18_i_q_d_1;
  yt_rsc_4_18_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_4_18_i_wadr_d <= yt_rsc_4_2_i_wadr_d_iff;

  yt_rsc_4_19_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_154_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_4_19_clkr_en,
      clkw_en => yt_rsc_4_19_clkw_en,
      q => yt_rsc_4_19_i_q,
      radr => yt_rsc_4_19_i_radr,
      we => yt_rsc_4_19_we,
      d => yt_rsc_4_19_i_d,
      wadr => yt_rsc_4_19_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_4_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_4_16_i_clkr_en_d,
      d_d => yt_rsc_4_19_i_d_d,
      q_d => yt_rsc_4_19_i_q_d_1,
      radr_d => yt_rsc_4_19_i_radr_d,
      wadr_d => yt_rsc_4_19_i_wadr_d,
      we_d => yt_rsc_4_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_4_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_4_19_i_q <= yt_rsc_4_19_q;
  yt_rsc_4_19_radr <= yt_rsc_4_19_i_radr;
  yt_rsc_4_19_d <= yt_rsc_4_19_i_d;
  yt_rsc_4_19_wadr <= yt_rsc_4_19_i_wadr;
  yt_rsc_4_19_i_d_d <= yt_rsc_4_3_i_d_d_iff;
  yt_rsc_4_19_i_q_d <= yt_rsc_4_19_i_q_d_1;
  yt_rsc_4_19_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_4_19_i_wadr_d <= yt_rsc_4_3_i_wadr_d_iff;

  yt_rsc_4_20_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_155_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_4_20_clkr_en,
      clkw_en => yt_rsc_4_20_clkw_en,
      q => yt_rsc_4_20_i_q,
      radr => yt_rsc_4_20_i_radr,
      we => yt_rsc_4_20_we,
      d => yt_rsc_4_20_i_d,
      wadr => yt_rsc_4_20_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_4_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_4_16_i_clkr_en_d,
      d_d => yt_rsc_4_20_i_d_d,
      q_d => yt_rsc_4_20_i_q_d_1,
      radr_d => yt_rsc_4_20_i_radr_d,
      wadr_d => yt_rsc_4_20_i_wadr_d,
      we_d => yt_rsc_4_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_4_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_4_20_i_q <= yt_rsc_4_20_q;
  yt_rsc_4_20_radr <= yt_rsc_4_20_i_radr;
  yt_rsc_4_20_d <= yt_rsc_4_20_i_d;
  yt_rsc_4_20_wadr <= yt_rsc_4_20_i_wadr;
  yt_rsc_4_20_i_d_d <= yt_rsc_4_4_i_d_d_iff;
  yt_rsc_4_20_i_q_d <= yt_rsc_4_20_i_q_d_1;
  yt_rsc_4_20_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_4_20_i_wadr_d <= yt_rsc_4_4_i_wadr_d_iff;

  yt_rsc_4_21_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_156_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_4_21_clkr_en,
      clkw_en => yt_rsc_4_21_clkw_en,
      q => yt_rsc_4_21_i_q,
      radr => yt_rsc_4_21_i_radr,
      we => yt_rsc_4_21_we,
      d => yt_rsc_4_21_i_d,
      wadr => yt_rsc_4_21_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_4_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_4_16_i_clkr_en_d,
      d_d => yt_rsc_4_21_i_d_d,
      q_d => yt_rsc_4_21_i_q_d_1,
      radr_d => yt_rsc_4_21_i_radr_d,
      wadr_d => yt_rsc_4_21_i_wadr_d,
      we_d => yt_rsc_4_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_4_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_4_21_i_q <= yt_rsc_4_21_q;
  yt_rsc_4_21_radr <= yt_rsc_4_21_i_radr;
  yt_rsc_4_21_d <= yt_rsc_4_21_i_d;
  yt_rsc_4_21_wadr <= yt_rsc_4_21_i_wadr;
  yt_rsc_4_21_i_d_d <= yt_rsc_4_5_i_d_d_iff;
  yt_rsc_4_21_i_q_d <= yt_rsc_4_21_i_q_d_1;
  yt_rsc_4_21_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_4_21_i_wadr_d <= yt_rsc_4_5_i_wadr_d_iff;

  yt_rsc_4_22_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_157_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_4_22_clkr_en,
      clkw_en => yt_rsc_4_22_clkw_en,
      q => yt_rsc_4_22_i_q,
      radr => yt_rsc_4_22_i_radr,
      we => yt_rsc_4_22_we,
      d => yt_rsc_4_22_i_d,
      wadr => yt_rsc_4_22_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_4_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_4_16_i_clkr_en_d,
      d_d => yt_rsc_4_22_i_d_d,
      q_d => yt_rsc_4_22_i_q_d_1,
      radr_d => yt_rsc_4_22_i_radr_d,
      wadr_d => yt_rsc_4_22_i_wadr_d,
      we_d => yt_rsc_4_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_4_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_4_22_i_q <= yt_rsc_4_22_q;
  yt_rsc_4_22_radr <= yt_rsc_4_22_i_radr;
  yt_rsc_4_22_d <= yt_rsc_4_22_i_d;
  yt_rsc_4_22_wadr <= yt_rsc_4_22_i_wadr;
  yt_rsc_4_22_i_d_d <= yt_rsc_4_6_i_d_d_iff;
  yt_rsc_4_22_i_q_d <= yt_rsc_4_22_i_q_d_1;
  yt_rsc_4_22_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_4_22_i_wadr_d <= yt_rsc_4_6_i_wadr_d_iff;

  yt_rsc_4_23_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_158_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_4_23_clkr_en,
      clkw_en => yt_rsc_4_23_clkw_en,
      q => yt_rsc_4_23_i_q,
      radr => yt_rsc_4_23_i_radr,
      we => yt_rsc_4_23_we,
      d => yt_rsc_4_23_i_d,
      wadr => yt_rsc_4_23_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_4_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_4_16_i_clkr_en_d,
      d_d => yt_rsc_4_23_i_d_d,
      q_d => yt_rsc_4_23_i_q_d_1,
      radr_d => yt_rsc_4_23_i_radr_d,
      wadr_d => yt_rsc_4_23_i_wadr_d,
      we_d => yt_rsc_4_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_4_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_4_23_i_q <= yt_rsc_4_23_q;
  yt_rsc_4_23_radr <= yt_rsc_4_23_i_radr;
  yt_rsc_4_23_d <= yt_rsc_4_23_i_d;
  yt_rsc_4_23_wadr <= yt_rsc_4_23_i_wadr;
  yt_rsc_4_23_i_d_d <= yt_rsc_4_7_i_d_d_iff;
  yt_rsc_4_23_i_q_d <= yt_rsc_4_23_i_q_d_1;
  yt_rsc_4_23_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_4_23_i_wadr_d <= yt_rsc_4_0_i_wadr_d_iff;

  yt_rsc_4_24_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_159_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_4_24_clkr_en,
      clkw_en => yt_rsc_4_24_clkw_en,
      q => yt_rsc_4_24_i_q,
      radr => yt_rsc_4_24_i_radr,
      we => yt_rsc_4_24_we,
      d => yt_rsc_4_24_i_d,
      wadr => yt_rsc_4_24_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_4_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_4_16_i_clkr_en_d,
      d_d => yt_rsc_4_24_i_d_d,
      q_d => yt_rsc_4_24_i_q_d_1,
      radr_d => yt_rsc_4_24_i_radr_d,
      wadr_d => yt_rsc_4_24_i_wadr_d,
      we_d => yt_rsc_4_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_4_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_4_24_i_q <= yt_rsc_4_24_q;
  yt_rsc_4_24_radr <= yt_rsc_4_24_i_radr;
  yt_rsc_4_24_d <= yt_rsc_4_24_i_d;
  yt_rsc_4_24_wadr <= yt_rsc_4_24_i_wadr;
  yt_rsc_4_24_i_d_d <= yt_rsc_4_8_i_d_d_iff;
  yt_rsc_4_24_i_q_d <= yt_rsc_4_24_i_q_d_1;
  yt_rsc_4_24_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_4_24_i_wadr_d <= yt_rsc_4_1_i_wadr_d_iff;

  yt_rsc_4_25_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_160_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_4_25_clkr_en,
      clkw_en => yt_rsc_4_25_clkw_en,
      q => yt_rsc_4_25_i_q,
      radr => yt_rsc_4_25_i_radr,
      we => yt_rsc_4_25_we,
      d => yt_rsc_4_25_i_d,
      wadr => yt_rsc_4_25_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_4_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_4_16_i_clkr_en_d,
      d_d => yt_rsc_4_25_i_d_d,
      q_d => yt_rsc_4_25_i_q_d_1,
      radr_d => yt_rsc_4_25_i_radr_d,
      wadr_d => yt_rsc_4_25_i_wadr_d,
      we_d => yt_rsc_4_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_4_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_4_25_i_q <= yt_rsc_4_25_q;
  yt_rsc_4_25_radr <= yt_rsc_4_25_i_radr;
  yt_rsc_4_25_d <= yt_rsc_4_25_i_d;
  yt_rsc_4_25_wadr <= yt_rsc_4_25_i_wadr;
  yt_rsc_4_25_i_d_d <= yt_rsc_4_9_i_d_d_iff;
  yt_rsc_4_25_i_q_d <= yt_rsc_4_25_i_q_d_1;
  yt_rsc_4_25_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_4_25_i_wadr_d <= yt_rsc_4_9_i_wadr_d_iff;

  yt_rsc_4_26_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_161_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_4_26_clkr_en,
      clkw_en => yt_rsc_4_26_clkw_en,
      q => yt_rsc_4_26_i_q,
      radr => yt_rsc_4_26_i_radr,
      we => yt_rsc_4_26_we,
      d => yt_rsc_4_26_i_d,
      wadr => yt_rsc_4_26_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_4_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_4_16_i_clkr_en_d,
      d_d => yt_rsc_4_26_i_d_d,
      q_d => yt_rsc_4_26_i_q_d_1,
      radr_d => yt_rsc_4_26_i_radr_d,
      wadr_d => yt_rsc_4_26_i_wadr_d,
      we_d => yt_rsc_4_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_4_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_4_26_i_q <= yt_rsc_4_26_q;
  yt_rsc_4_26_radr <= yt_rsc_4_26_i_radr;
  yt_rsc_4_26_d <= yt_rsc_4_26_i_d;
  yt_rsc_4_26_wadr <= yt_rsc_4_26_i_wadr;
  yt_rsc_4_26_i_d_d <= yt_rsc_4_10_i_d_d_iff;
  yt_rsc_4_26_i_q_d <= yt_rsc_4_26_i_q_d_1;
  yt_rsc_4_26_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_4_26_i_wadr_d <= yt_rsc_4_10_i_wadr_d_iff;

  yt_rsc_4_27_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_162_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_4_27_clkr_en,
      clkw_en => yt_rsc_4_27_clkw_en,
      q => yt_rsc_4_27_i_q,
      radr => yt_rsc_4_27_i_radr,
      we => yt_rsc_4_27_we,
      d => yt_rsc_4_27_i_d,
      wadr => yt_rsc_4_27_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_4_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_4_16_i_clkr_en_d,
      d_d => yt_rsc_4_27_i_d_d,
      q_d => yt_rsc_4_27_i_q_d_1,
      radr_d => yt_rsc_4_27_i_radr_d,
      wadr_d => yt_rsc_4_27_i_wadr_d,
      we_d => yt_rsc_4_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_4_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_4_27_i_q <= yt_rsc_4_27_q;
  yt_rsc_4_27_radr <= yt_rsc_4_27_i_radr;
  yt_rsc_4_27_d <= yt_rsc_4_27_i_d;
  yt_rsc_4_27_wadr <= yt_rsc_4_27_i_wadr;
  yt_rsc_4_27_i_d_d <= yt_rsc_4_11_i_d_d_iff;
  yt_rsc_4_27_i_q_d <= yt_rsc_4_27_i_q_d_1;
  yt_rsc_4_27_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_4_27_i_wadr_d <= yt_rsc_4_11_i_wadr_d_iff;

  yt_rsc_4_28_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_163_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_4_28_clkr_en,
      clkw_en => yt_rsc_4_28_clkw_en,
      q => yt_rsc_4_28_i_q,
      radr => yt_rsc_4_28_i_radr,
      we => yt_rsc_4_28_we,
      d => yt_rsc_4_28_i_d,
      wadr => yt_rsc_4_28_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_4_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_4_16_i_clkr_en_d,
      d_d => yt_rsc_4_28_i_d_d,
      q_d => yt_rsc_4_28_i_q_d_1,
      radr_d => yt_rsc_4_28_i_radr_d,
      wadr_d => yt_rsc_4_28_i_wadr_d,
      we_d => yt_rsc_4_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_4_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_4_28_i_q <= yt_rsc_4_28_q;
  yt_rsc_4_28_radr <= yt_rsc_4_28_i_radr;
  yt_rsc_4_28_d <= yt_rsc_4_28_i_d;
  yt_rsc_4_28_wadr <= yt_rsc_4_28_i_wadr;
  yt_rsc_4_28_i_d_d <= yt_rsc_4_12_i_d_d_iff;
  yt_rsc_4_28_i_q_d <= yt_rsc_4_28_i_q_d_1;
  yt_rsc_4_28_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_4_28_i_wadr_d <= yt_rsc_4_3_i_wadr_d_iff;

  yt_rsc_4_29_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_164_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_4_29_clkr_en,
      clkw_en => yt_rsc_4_29_clkw_en,
      q => yt_rsc_4_29_i_q,
      radr => yt_rsc_4_29_i_radr,
      we => yt_rsc_4_29_we,
      d => yt_rsc_4_29_i_d,
      wadr => yt_rsc_4_29_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_4_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_4_16_i_clkr_en_d,
      d_d => yt_rsc_4_29_i_d_d,
      q_d => yt_rsc_4_29_i_q_d_1,
      radr_d => yt_rsc_4_29_i_radr_d,
      wadr_d => yt_rsc_4_29_i_wadr_d,
      we_d => yt_rsc_4_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_4_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_4_29_i_q <= yt_rsc_4_29_q;
  yt_rsc_4_29_radr <= yt_rsc_4_29_i_radr;
  yt_rsc_4_29_d <= yt_rsc_4_29_i_d;
  yt_rsc_4_29_wadr <= yt_rsc_4_29_i_wadr;
  yt_rsc_4_29_i_d_d <= yt_rsc_4_13_i_d_d_iff;
  yt_rsc_4_29_i_q_d <= yt_rsc_4_29_i_q_d_1;
  yt_rsc_4_29_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_4_29_i_wadr_d <= yt_rsc_4_4_i_wadr_d_iff;

  yt_rsc_4_30_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_165_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_4_30_clkr_en,
      clkw_en => yt_rsc_4_30_clkw_en,
      q => yt_rsc_4_30_i_q,
      radr => yt_rsc_4_30_i_radr,
      we => yt_rsc_4_30_we,
      d => yt_rsc_4_30_i_d,
      wadr => yt_rsc_4_30_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_4_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_4_16_i_clkr_en_d,
      d_d => yt_rsc_4_30_i_d_d,
      q_d => yt_rsc_4_30_i_q_d_1,
      radr_d => yt_rsc_4_30_i_radr_d,
      wadr_d => yt_rsc_4_30_i_wadr_d,
      we_d => yt_rsc_4_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_4_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_4_30_i_q <= yt_rsc_4_30_q;
  yt_rsc_4_30_radr <= yt_rsc_4_30_i_radr;
  yt_rsc_4_30_d <= yt_rsc_4_30_i_d;
  yt_rsc_4_30_wadr <= yt_rsc_4_30_i_wadr;
  yt_rsc_4_30_i_d_d <= yt_rsc_4_14_i_d_d_iff;
  yt_rsc_4_30_i_q_d <= yt_rsc_4_30_i_q_d_1;
  yt_rsc_4_30_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_4_30_i_wadr_d <= yt_rsc_4_5_i_wadr_d_iff;

  yt_rsc_4_31_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_166_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_4_31_clkr_en,
      clkw_en => yt_rsc_4_31_clkw_en,
      q => yt_rsc_4_31_i_q,
      radr => yt_rsc_4_31_i_radr,
      we => yt_rsc_4_31_we,
      d => yt_rsc_4_31_i_d,
      wadr => yt_rsc_4_31_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_4_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_4_16_i_clkr_en_d,
      d_d => yt_rsc_4_31_i_d_d,
      q_d => yt_rsc_4_31_i_q_d_1,
      radr_d => yt_rsc_4_31_i_radr_d,
      wadr_d => yt_rsc_4_31_i_wadr_d,
      we_d => yt_rsc_4_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_4_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_4_31_i_q <= yt_rsc_4_31_q;
  yt_rsc_4_31_radr <= yt_rsc_4_31_i_radr;
  yt_rsc_4_31_d <= yt_rsc_4_31_i_d;
  yt_rsc_4_31_wadr <= yt_rsc_4_31_i_wadr;
  yt_rsc_4_31_i_d_d <= yt_rsc_4_15_i_d_d_iff;
  yt_rsc_4_31_i_q_d <= yt_rsc_4_31_i_q_d_1;
  yt_rsc_4_31_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_4_31_i_wadr_d <= yt_rsc_4_6_i_wadr_d_iff;

  yt_rsc_5_0_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_167_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_5_0_clkr_en,
      clkw_en => yt_rsc_5_0_clkw_en,
      q => yt_rsc_5_0_i_q,
      radr => yt_rsc_5_0_i_radr,
      we => yt_rsc_5_0_we,
      d => yt_rsc_5_0_i_d,
      wadr => yt_rsc_5_0_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_5_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_5_0_i_clkr_en_d,
      d_d => yt_rsc_5_0_i_d_d,
      q_d => yt_rsc_5_0_i_q_d_1,
      radr_d => yt_rsc_5_0_i_radr_d,
      wadr_d => yt_rsc_5_0_i_wadr_d,
      we_d => yt_rsc_5_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_5_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_5_0_i_q <= yt_rsc_5_0_q;
  yt_rsc_5_0_radr <= yt_rsc_5_0_i_radr;
  yt_rsc_5_0_d <= yt_rsc_5_0_i_d;
  yt_rsc_5_0_wadr <= yt_rsc_5_0_i_wadr;
  yt_rsc_5_0_i_d_d <= yt_rsc_4_0_i_d_d_iff;
  yt_rsc_5_0_i_q_d <= yt_rsc_5_0_i_q_d_1;
  yt_rsc_5_0_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_5_0_i_wadr_d <= yt_rsc_4_0_i_wadr_d_iff;

  yt_rsc_5_1_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_168_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_5_1_clkr_en,
      clkw_en => yt_rsc_5_1_clkw_en,
      q => yt_rsc_5_1_i_q,
      radr => yt_rsc_5_1_i_radr,
      we => yt_rsc_5_1_we,
      d => yt_rsc_5_1_i_d,
      wadr => yt_rsc_5_1_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_5_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_5_0_i_clkr_en_d,
      d_d => yt_rsc_5_1_i_d_d,
      q_d => yt_rsc_5_1_i_q_d_1,
      radr_d => yt_rsc_5_1_i_radr_d,
      wadr_d => yt_rsc_5_1_i_wadr_d,
      we_d => yt_rsc_5_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_5_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_5_1_i_q <= yt_rsc_5_1_q;
  yt_rsc_5_1_radr <= yt_rsc_5_1_i_radr;
  yt_rsc_5_1_d <= yt_rsc_5_1_i_d;
  yt_rsc_5_1_wadr <= yt_rsc_5_1_i_wadr;
  yt_rsc_5_1_i_d_d <= yt_rsc_4_1_i_d_d_iff;
  yt_rsc_5_1_i_q_d <= yt_rsc_5_1_i_q_d_1;
  yt_rsc_5_1_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_5_1_i_wadr_d <= yt_rsc_4_1_i_wadr_d_iff;

  yt_rsc_5_2_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_169_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_5_2_clkr_en,
      clkw_en => yt_rsc_5_2_clkw_en,
      q => yt_rsc_5_2_i_q,
      radr => yt_rsc_5_2_i_radr,
      we => yt_rsc_5_2_we,
      d => yt_rsc_5_2_i_d,
      wadr => yt_rsc_5_2_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_5_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_5_0_i_clkr_en_d,
      d_d => yt_rsc_5_2_i_d_d,
      q_d => yt_rsc_5_2_i_q_d_1,
      radr_d => yt_rsc_5_2_i_radr_d,
      wadr_d => yt_rsc_5_2_i_wadr_d,
      we_d => yt_rsc_5_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_5_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_5_2_i_q <= yt_rsc_5_2_q;
  yt_rsc_5_2_radr <= yt_rsc_5_2_i_radr;
  yt_rsc_5_2_d <= yt_rsc_5_2_i_d;
  yt_rsc_5_2_wadr <= yt_rsc_5_2_i_wadr;
  yt_rsc_5_2_i_d_d <= yt_rsc_4_2_i_d_d_iff;
  yt_rsc_5_2_i_q_d <= yt_rsc_5_2_i_q_d_1;
  yt_rsc_5_2_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_5_2_i_wadr_d <= yt_rsc_4_2_i_wadr_d_iff;

  yt_rsc_5_3_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_170_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_5_3_clkr_en,
      clkw_en => yt_rsc_5_3_clkw_en,
      q => yt_rsc_5_3_i_q,
      radr => yt_rsc_5_3_i_radr,
      we => yt_rsc_5_3_we,
      d => yt_rsc_5_3_i_d,
      wadr => yt_rsc_5_3_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_5_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_5_0_i_clkr_en_d,
      d_d => yt_rsc_5_3_i_d_d,
      q_d => yt_rsc_5_3_i_q_d_1,
      radr_d => yt_rsc_5_3_i_radr_d,
      wadr_d => yt_rsc_5_3_i_wadr_d,
      we_d => yt_rsc_5_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_5_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_5_3_i_q <= yt_rsc_5_3_q;
  yt_rsc_5_3_radr <= yt_rsc_5_3_i_radr;
  yt_rsc_5_3_d <= yt_rsc_5_3_i_d;
  yt_rsc_5_3_wadr <= yt_rsc_5_3_i_wadr;
  yt_rsc_5_3_i_d_d <= yt_rsc_4_3_i_d_d_iff;
  yt_rsc_5_3_i_q_d <= yt_rsc_5_3_i_q_d_1;
  yt_rsc_5_3_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_5_3_i_wadr_d <= yt_rsc_4_3_i_wadr_d_iff;

  yt_rsc_5_4_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_171_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_5_4_clkr_en,
      clkw_en => yt_rsc_5_4_clkw_en,
      q => yt_rsc_5_4_i_q,
      radr => yt_rsc_5_4_i_radr,
      we => yt_rsc_5_4_we,
      d => yt_rsc_5_4_i_d,
      wadr => yt_rsc_5_4_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_5_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_5_0_i_clkr_en_d,
      d_d => yt_rsc_5_4_i_d_d,
      q_d => yt_rsc_5_4_i_q_d_1,
      radr_d => yt_rsc_5_4_i_radr_d,
      wadr_d => yt_rsc_5_4_i_wadr_d,
      we_d => yt_rsc_5_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_5_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_5_4_i_q <= yt_rsc_5_4_q;
  yt_rsc_5_4_radr <= yt_rsc_5_4_i_radr;
  yt_rsc_5_4_d <= yt_rsc_5_4_i_d;
  yt_rsc_5_4_wadr <= yt_rsc_5_4_i_wadr;
  yt_rsc_5_4_i_d_d <= yt_rsc_4_4_i_d_d_iff;
  yt_rsc_5_4_i_q_d <= yt_rsc_5_4_i_q_d_1;
  yt_rsc_5_4_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_5_4_i_wadr_d <= yt_rsc_4_4_i_wadr_d_iff;

  yt_rsc_5_5_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_172_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_5_5_clkr_en,
      clkw_en => yt_rsc_5_5_clkw_en,
      q => yt_rsc_5_5_i_q,
      radr => yt_rsc_5_5_i_radr,
      we => yt_rsc_5_5_we,
      d => yt_rsc_5_5_i_d,
      wadr => yt_rsc_5_5_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_5_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_5_0_i_clkr_en_d,
      d_d => yt_rsc_5_5_i_d_d,
      q_d => yt_rsc_5_5_i_q_d_1,
      radr_d => yt_rsc_5_5_i_radr_d,
      wadr_d => yt_rsc_5_5_i_wadr_d,
      we_d => yt_rsc_5_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_5_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_5_5_i_q <= yt_rsc_5_5_q;
  yt_rsc_5_5_radr <= yt_rsc_5_5_i_radr;
  yt_rsc_5_5_d <= yt_rsc_5_5_i_d;
  yt_rsc_5_5_wadr <= yt_rsc_5_5_i_wadr;
  yt_rsc_5_5_i_d_d <= yt_rsc_4_5_i_d_d_iff;
  yt_rsc_5_5_i_q_d <= yt_rsc_5_5_i_q_d_1;
  yt_rsc_5_5_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_5_5_i_wadr_d <= yt_rsc_4_5_i_wadr_d_iff;

  yt_rsc_5_6_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_173_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_5_6_clkr_en,
      clkw_en => yt_rsc_5_6_clkw_en,
      q => yt_rsc_5_6_i_q,
      radr => yt_rsc_5_6_i_radr,
      we => yt_rsc_5_6_we,
      d => yt_rsc_5_6_i_d,
      wadr => yt_rsc_5_6_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_5_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_5_0_i_clkr_en_d,
      d_d => yt_rsc_5_6_i_d_d,
      q_d => yt_rsc_5_6_i_q_d_1,
      radr_d => yt_rsc_5_6_i_radr_d,
      wadr_d => yt_rsc_5_6_i_wadr_d,
      we_d => yt_rsc_5_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_5_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_5_6_i_q <= yt_rsc_5_6_q;
  yt_rsc_5_6_radr <= yt_rsc_5_6_i_radr;
  yt_rsc_5_6_d <= yt_rsc_5_6_i_d;
  yt_rsc_5_6_wadr <= yt_rsc_5_6_i_wadr;
  yt_rsc_5_6_i_d_d <= yt_rsc_4_6_i_d_d_iff;
  yt_rsc_5_6_i_q_d <= yt_rsc_5_6_i_q_d_1;
  yt_rsc_5_6_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_5_6_i_wadr_d <= yt_rsc_4_6_i_wadr_d_iff;

  yt_rsc_5_7_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_174_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_5_7_clkr_en,
      clkw_en => yt_rsc_5_7_clkw_en,
      q => yt_rsc_5_7_i_q,
      radr => yt_rsc_5_7_i_radr,
      we => yt_rsc_5_7_we,
      d => yt_rsc_5_7_i_d,
      wadr => yt_rsc_5_7_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_5_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_5_0_i_clkr_en_d,
      d_d => yt_rsc_5_7_i_d_d,
      q_d => yt_rsc_5_7_i_q_d_1,
      radr_d => yt_rsc_5_7_i_radr_d,
      wadr_d => yt_rsc_5_7_i_wadr_d,
      we_d => yt_rsc_5_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_5_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_5_7_i_q <= yt_rsc_5_7_q;
  yt_rsc_5_7_radr <= yt_rsc_5_7_i_radr;
  yt_rsc_5_7_d <= yt_rsc_5_7_i_d;
  yt_rsc_5_7_wadr <= yt_rsc_5_7_i_wadr;
  yt_rsc_5_7_i_d_d <= yt_rsc_4_7_i_d_d_iff;
  yt_rsc_5_7_i_q_d <= yt_rsc_5_7_i_q_d_1;
  yt_rsc_5_7_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_5_7_i_wadr_d <= yt_rsc_4_0_i_wadr_d_iff;

  yt_rsc_5_8_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_175_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_5_8_clkr_en,
      clkw_en => yt_rsc_5_8_clkw_en,
      q => yt_rsc_5_8_i_q,
      radr => yt_rsc_5_8_i_radr,
      we => yt_rsc_5_8_we,
      d => yt_rsc_5_8_i_d,
      wadr => yt_rsc_5_8_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_5_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_5_0_i_clkr_en_d,
      d_d => yt_rsc_5_8_i_d_d,
      q_d => yt_rsc_5_8_i_q_d_1,
      radr_d => yt_rsc_5_8_i_radr_d,
      wadr_d => yt_rsc_5_8_i_wadr_d,
      we_d => yt_rsc_5_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_5_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_5_8_i_q <= yt_rsc_5_8_q;
  yt_rsc_5_8_radr <= yt_rsc_5_8_i_radr;
  yt_rsc_5_8_d <= yt_rsc_5_8_i_d;
  yt_rsc_5_8_wadr <= yt_rsc_5_8_i_wadr;
  yt_rsc_5_8_i_d_d <= yt_rsc_4_8_i_d_d_iff;
  yt_rsc_5_8_i_q_d <= yt_rsc_5_8_i_q_d_1;
  yt_rsc_5_8_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_5_8_i_wadr_d <= yt_rsc_4_1_i_wadr_d_iff;

  yt_rsc_5_9_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_176_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_5_9_clkr_en,
      clkw_en => yt_rsc_5_9_clkw_en,
      q => yt_rsc_5_9_i_q,
      radr => yt_rsc_5_9_i_radr,
      we => yt_rsc_5_9_we,
      d => yt_rsc_5_9_i_d,
      wadr => yt_rsc_5_9_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_5_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_5_0_i_clkr_en_d,
      d_d => yt_rsc_5_9_i_d_d,
      q_d => yt_rsc_5_9_i_q_d_1,
      radr_d => yt_rsc_5_9_i_radr_d,
      wadr_d => yt_rsc_5_9_i_wadr_d,
      we_d => yt_rsc_5_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_5_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_5_9_i_q <= yt_rsc_5_9_q;
  yt_rsc_5_9_radr <= yt_rsc_5_9_i_radr;
  yt_rsc_5_9_d <= yt_rsc_5_9_i_d;
  yt_rsc_5_9_wadr <= yt_rsc_5_9_i_wadr;
  yt_rsc_5_9_i_d_d <= yt_rsc_4_9_i_d_d_iff;
  yt_rsc_5_9_i_q_d <= yt_rsc_5_9_i_q_d_1;
  yt_rsc_5_9_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_5_9_i_wadr_d <= yt_rsc_4_9_i_wadr_d_iff;

  yt_rsc_5_10_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_177_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_5_10_clkr_en,
      clkw_en => yt_rsc_5_10_clkw_en,
      q => yt_rsc_5_10_i_q,
      radr => yt_rsc_5_10_i_radr,
      we => yt_rsc_5_10_we,
      d => yt_rsc_5_10_i_d,
      wadr => yt_rsc_5_10_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_5_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_5_0_i_clkr_en_d,
      d_d => yt_rsc_5_10_i_d_d,
      q_d => yt_rsc_5_10_i_q_d_1,
      radr_d => yt_rsc_5_10_i_radr_d,
      wadr_d => yt_rsc_5_10_i_wadr_d,
      we_d => yt_rsc_5_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_5_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_5_10_i_q <= yt_rsc_5_10_q;
  yt_rsc_5_10_radr <= yt_rsc_5_10_i_radr;
  yt_rsc_5_10_d <= yt_rsc_5_10_i_d;
  yt_rsc_5_10_wadr <= yt_rsc_5_10_i_wadr;
  yt_rsc_5_10_i_d_d <= yt_rsc_4_10_i_d_d_iff;
  yt_rsc_5_10_i_q_d <= yt_rsc_5_10_i_q_d_1;
  yt_rsc_5_10_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_5_10_i_wadr_d <= yt_rsc_4_10_i_wadr_d_iff;

  yt_rsc_5_11_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_178_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_5_11_clkr_en,
      clkw_en => yt_rsc_5_11_clkw_en,
      q => yt_rsc_5_11_i_q,
      radr => yt_rsc_5_11_i_radr,
      we => yt_rsc_5_11_we,
      d => yt_rsc_5_11_i_d,
      wadr => yt_rsc_5_11_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_5_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_5_0_i_clkr_en_d,
      d_d => yt_rsc_5_11_i_d_d,
      q_d => yt_rsc_5_11_i_q_d_1,
      radr_d => yt_rsc_5_11_i_radr_d,
      wadr_d => yt_rsc_5_11_i_wadr_d,
      we_d => yt_rsc_5_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_5_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_5_11_i_q <= yt_rsc_5_11_q;
  yt_rsc_5_11_radr <= yt_rsc_5_11_i_radr;
  yt_rsc_5_11_d <= yt_rsc_5_11_i_d;
  yt_rsc_5_11_wadr <= yt_rsc_5_11_i_wadr;
  yt_rsc_5_11_i_d_d <= yt_rsc_4_11_i_d_d_iff;
  yt_rsc_5_11_i_q_d <= yt_rsc_5_11_i_q_d_1;
  yt_rsc_5_11_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_5_11_i_wadr_d <= yt_rsc_4_11_i_wadr_d_iff;

  yt_rsc_5_12_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_179_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_5_12_clkr_en,
      clkw_en => yt_rsc_5_12_clkw_en,
      q => yt_rsc_5_12_i_q,
      radr => yt_rsc_5_12_i_radr,
      we => yt_rsc_5_12_we,
      d => yt_rsc_5_12_i_d,
      wadr => yt_rsc_5_12_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_5_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_5_0_i_clkr_en_d,
      d_d => yt_rsc_5_12_i_d_d,
      q_d => yt_rsc_5_12_i_q_d_1,
      radr_d => yt_rsc_5_12_i_radr_d,
      wadr_d => yt_rsc_5_12_i_wadr_d,
      we_d => yt_rsc_5_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_5_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_5_12_i_q <= yt_rsc_5_12_q;
  yt_rsc_5_12_radr <= yt_rsc_5_12_i_radr;
  yt_rsc_5_12_d <= yt_rsc_5_12_i_d;
  yt_rsc_5_12_wadr <= yt_rsc_5_12_i_wadr;
  yt_rsc_5_12_i_d_d <= yt_rsc_4_12_i_d_d_iff;
  yt_rsc_5_12_i_q_d <= yt_rsc_5_12_i_q_d_1;
  yt_rsc_5_12_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_5_12_i_wadr_d <= yt_rsc_4_3_i_wadr_d_iff;

  yt_rsc_5_13_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_180_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_5_13_clkr_en,
      clkw_en => yt_rsc_5_13_clkw_en,
      q => yt_rsc_5_13_i_q,
      radr => yt_rsc_5_13_i_radr,
      we => yt_rsc_5_13_we,
      d => yt_rsc_5_13_i_d,
      wadr => yt_rsc_5_13_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_5_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_5_0_i_clkr_en_d,
      d_d => yt_rsc_5_13_i_d_d,
      q_d => yt_rsc_5_13_i_q_d_1,
      radr_d => yt_rsc_5_13_i_radr_d,
      wadr_d => yt_rsc_5_13_i_wadr_d,
      we_d => yt_rsc_5_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_5_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_5_13_i_q <= yt_rsc_5_13_q;
  yt_rsc_5_13_radr <= yt_rsc_5_13_i_radr;
  yt_rsc_5_13_d <= yt_rsc_5_13_i_d;
  yt_rsc_5_13_wadr <= yt_rsc_5_13_i_wadr;
  yt_rsc_5_13_i_d_d <= yt_rsc_4_13_i_d_d_iff;
  yt_rsc_5_13_i_q_d <= yt_rsc_5_13_i_q_d_1;
  yt_rsc_5_13_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_5_13_i_wadr_d <= yt_rsc_4_4_i_wadr_d_iff;

  yt_rsc_5_14_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_181_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_5_14_clkr_en,
      clkw_en => yt_rsc_5_14_clkw_en,
      q => yt_rsc_5_14_i_q,
      radr => yt_rsc_5_14_i_radr,
      we => yt_rsc_5_14_we,
      d => yt_rsc_5_14_i_d,
      wadr => yt_rsc_5_14_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_5_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_5_0_i_clkr_en_d,
      d_d => yt_rsc_5_14_i_d_d,
      q_d => yt_rsc_5_14_i_q_d_1,
      radr_d => yt_rsc_5_14_i_radr_d,
      wadr_d => yt_rsc_5_14_i_wadr_d,
      we_d => yt_rsc_5_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_5_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_5_14_i_q <= yt_rsc_5_14_q;
  yt_rsc_5_14_radr <= yt_rsc_5_14_i_radr;
  yt_rsc_5_14_d <= yt_rsc_5_14_i_d;
  yt_rsc_5_14_wadr <= yt_rsc_5_14_i_wadr;
  yt_rsc_5_14_i_d_d <= yt_rsc_4_14_i_d_d_iff;
  yt_rsc_5_14_i_q_d <= yt_rsc_5_14_i_q_d_1;
  yt_rsc_5_14_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_5_14_i_wadr_d <= yt_rsc_4_5_i_wadr_d_iff;

  yt_rsc_5_15_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_182_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_5_15_clkr_en,
      clkw_en => yt_rsc_5_15_clkw_en,
      q => yt_rsc_5_15_i_q,
      radr => yt_rsc_5_15_i_radr,
      we => yt_rsc_5_15_we,
      d => yt_rsc_5_15_i_d,
      wadr => yt_rsc_5_15_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_5_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_5_0_i_clkr_en_d,
      d_d => yt_rsc_5_15_i_d_d,
      q_d => yt_rsc_5_15_i_q_d_1,
      radr_d => yt_rsc_5_15_i_radr_d,
      wadr_d => yt_rsc_5_15_i_wadr_d,
      we_d => yt_rsc_5_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_5_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_5_15_i_q <= yt_rsc_5_15_q;
  yt_rsc_5_15_radr <= yt_rsc_5_15_i_radr;
  yt_rsc_5_15_d <= yt_rsc_5_15_i_d;
  yt_rsc_5_15_wadr <= yt_rsc_5_15_i_wadr;
  yt_rsc_5_15_i_d_d <= yt_rsc_4_15_i_d_d_iff;
  yt_rsc_5_15_i_q_d <= yt_rsc_5_15_i_q_d_1;
  yt_rsc_5_15_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_5_15_i_wadr_d <= yt_rsc_4_6_i_wadr_d_iff;

  yt_rsc_5_16_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_183_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_5_16_clkr_en,
      clkw_en => yt_rsc_5_16_clkw_en,
      q => yt_rsc_5_16_i_q,
      radr => yt_rsc_5_16_i_radr,
      we => yt_rsc_5_16_we,
      d => yt_rsc_5_16_i_d,
      wadr => yt_rsc_5_16_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_5_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_5_16_i_clkr_en_d,
      d_d => yt_rsc_5_16_i_d_d,
      q_d => yt_rsc_5_16_i_q_d_1,
      radr_d => yt_rsc_5_16_i_radr_d,
      wadr_d => yt_rsc_5_16_i_wadr_d,
      we_d => yt_rsc_5_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_5_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_5_16_i_q <= yt_rsc_5_16_q;
  yt_rsc_5_16_radr <= yt_rsc_5_16_i_radr;
  yt_rsc_5_16_d <= yt_rsc_5_16_i_d;
  yt_rsc_5_16_wadr <= yt_rsc_5_16_i_wadr;
  yt_rsc_5_16_i_d_d <= yt_rsc_4_0_i_d_d_iff;
  yt_rsc_5_16_i_q_d <= yt_rsc_5_16_i_q_d_1;
  yt_rsc_5_16_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_5_16_i_wadr_d <= yt_rsc_4_0_i_wadr_d_iff;

  yt_rsc_5_17_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_184_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_5_17_clkr_en,
      clkw_en => yt_rsc_5_17_clkw_en,
      q => yt_rsc_5_17_i_q,
      radr => yt_rsc_5_17_i_radr,
      we => yt_rsc_5_17_we,
      d => yt_rsc_5_17_i_d,
      wadr => yt_rsc_5_17_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_5_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_5_16_i_clkr_en_d,
      d_d => yt_rsc_5_17_i_d_d,
      q_d => yt_rsc_5_17_i_q_d_1,
      radr_d => yt_rsc_5_17_i_radr_d,
      wadr_d => yt_rsc_5_17_i_wadr_d,
      we_d => yt_rsc_5_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_5_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_5_17_i_q <= yt_rsc_5_17_q;
  yt_rsc_5_17_radr <= yt_rsc_5_17_i_radr;
  yt_rsc_5_17_d <= yt_rsc_5_17_i_d;
  yt_rsc_5_17_wadr <= yt_rsc_5_17_i_wadr;
  yt_rsc_5_17_i_d_d <= yt_rsc_4_1_i_d_d_iff;
  yt_rsc_5_17_i_q_d <= yt_rsc_5_17_i_q_d_1;
  yt_rsc_5_17_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_5_17_i_wadr_d <= yt_rsc_4_1_i_wadr_d_iff;

  yt_rsc_5_18_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_185_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_5_18_clkr_en,
      clkw_en => yt_rsc_5_18_clkw_en,
      q => yt_rsc_5_18_i_q,
      radr => yt_rsc_5_18_i_radr,
      we => yt_rsc_5_18_we,
      d => yt_rsc_5_18_i_d,
      wadr => yt_rsc_5_18_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_5_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_5_16_i_clkr_en_d,
      d_d => yt_rsc_5_18_i_d_d,
      q_d => yt_rsc_5_18_i_q_d_1,
      radr_d => yt_rsc_5_18_i_radr_d,
      wadr_d => yt_rsc_5_18_i_wadr_d,
      we_d => yt_rsc_5_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_5_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_5_18_i_q <= yt_rsc_5_18_q;
  yt_rsc_5_18_radr <= yt_rsc_5_18_i_radr;
  yt_rsc_5_18_d <= yt_rsc_5_18_i_d;
  yt_rsc_5_18_wadr <= yt_rsc_5_18_i_wadr;
  yt_rsc_5_18_i_d_d <= yt_rsc_4_2_i_d_d_iff;
  yt_rsc_5_18_i_q_d <= yt_rsc_5_18_i_q_d_1;
  yt_rsc_5_18_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_5_18_i_wadr_d <= yt_rsc_4_2_i_wadr_d_iff;

  yt_rsc_5_19_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_186_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_5_19_clkr_en,
      clkw_en => yt_rsc_5_19_clkw_en,
      q => yt_rsc_5_19_i_q,
      radr => yt_rsc_5_19_i_radr,
      we => yt_rsc_5_19_we,
      d => yt_rsc_5_19_i_d,
      wadr => yt_rsc_5_19_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_5_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_5_16_i_clkr_en_d,
      d_d => yt_rsc_5_19_i_d_d,
      q_d => yt_rsc_5_19_i_q_d_1,
      radr_d => yt_rsc_5_19_i_radr_d,
      wadr_d => yt_rsc_5_19_i_wadr_d,
      we_d => yt_rsc_5_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_5_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_5_19_i_q <= yt_rsc_5_19_q;
  yt_rsc_5_19_radr <= yt_rsc_5_19_i_radr;
  yt_rsc_5_19_d <= yt_rsc_5_19_i_d;
  yt_rsc_5_19_wadr <= yt_rsc_5_19_i_wadr;
  yt_rsc_5_19_i_d_d <= yt_rsc_4_3_i_d_d_iff;
  yt_rsc_5_19_i_q_d <= yt_rsc_5_19_i_q_d_1;
  yt_rsc_5_19_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_5_19_i_wadr_d <= yt_rsc_4_3_i_wadr_d_iff;

  yt_rsc_5_20_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_187_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_5_20_clkr_en,
      clkw_en => yt_rsc_5_20_clkw_en,
      q => yt_rsc_5_20_i_q,
      radr => yt_rsc_5_20_i_radr,
      we => yt_rsc_5_20_we,
      d => yt_rsc_5_20_i_d,
      wadr => yt_rsc_5_20_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_5_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_5_16_i_clkr_en_d,
      d_d => yt_rsc_5_20_i_d_d,
      q_d => yt_rsc_5_20_i_q_d_1,
      radr_d => yt_rsc_5_20_i_radr_d,
      wadr_d => yt_rsc_5_20_i_wadr_d,
      we_d => yt_rsc_5_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_5_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_5_20_i_q <= yt_rsc_5_20_q;
  yt_rsc_5_20_radr <= yt_rsc_5_20_i_radr;
  yt_rsc_5_20_d <= yt_rsc_5_20_i_d;
  yt_rsc_5_20_wadr <= yt_rsc_5_20_i_wadr;
  yt_rsc_5_20_i_d_d <= yt_rsc_4_4_i_d_d_iff;
  yt_rsc_5_20_i_q_d <= yt_rsc_5_20_i_q_d_1;
  yt_rsc_5_20_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_5_20_i_wadr_d <= yt_rsc_4_4_i_wadr_d_iff;

  yt_rsc_5_21_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_188_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_5_21_clkr_en,
      clkw_en => yt_rsc_5_21_clkw_en,
      q => yt_rsc_5_21_i_q,
      radr => yt_rsc_5_21_i_radr,
      we => yt_rsc_5_21_we,
      d => yt_rsc_5_21_i_d,
      wadr => yt_rsc_5_21_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_5_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_5_16_i_clkr_en_d,
      d_d => yt_rsc_5_21_i_d_d,
      q_d => yt_rsc_5_21_i_q_d_1,
      radr_d => yt_rsc_5_21_i_radr_d,
      wadr_d => yt_rsc_5_21_i_wadr_d,
      we_d => yt_rsc_5_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_5_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_5_21_i_q <= yt_rsc_5_21_q;
  yt_rsc_5_21_radr <= yt_rsc_5_21_i_radr;
  yt_rsc_5_21_d <= yt_rsc_5_21_i_d;
  yt_rsc_5_21_wadr <= yt_rsc_5_21_i_wadr;
  yt_rsc_5_21_i_d_d <= yt_rsc_4_5_i_d_d_iff;
  yt_rsc_5_21_i_q_d <= yt_rsc_5_21_i_q_d_1;
  yt_rsc_5_21_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_5_21_i_wadr_d <= yt_rsc_4_5_i_wadr_d_iff;

  yt_rsc_5_22_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_189_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_5_22_clkr_en,
      clkw_en => yt_rsc_5_22_clkw_en,
      q => yt_rsc_5_22_i_q,
      radr => yt_rsc_5_22_i_radr,
      we => yt_rsc_5_22_we,
      d => yt_rsc_5_22_i_d,
      wadr => yt_rsc_5_22_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_5_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_5_16_i_clkr_en_d,
      d_d => yt_rsc_5_22_i_d_d,
      q_d => yt_rsc_5_22_i_q_d_1,
      radr_d => yt_rsc_5_22_i_radr_d,
      wadr_d => yt_rsc_5_22_i_wadr_d,
      we_d => yt_rsc_5_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_5_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_5_22_i_q <= yt_rsc_5_22_q;
  yt_rsc_5_22_radr <= yt_rsc_5_22_i_radr;
  yt_rsc_5_22_d <= yt_rsc_5_22_i_d;
  yt_rsc_5_22_wadr <= yt_rsc_5_22_i_wadr;
  yt_rsc_5_22_i_d_d <= yt_rsc_4_6_i_d_d_iff;
  yt_rsc_5_22_i_q_d <= yt_rsc_5_22_i_q_d_1;
  yt_rsc_5_22_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_5_22_i_wadr_d <= yt_rsc_4_6_i_wadr_d_iff;

  yt_rsc_5_23_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_190_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_5_23_clkr_en,
      clkw_en => yt_rsc_5_23_clkw_en,
      q => yt_rsc_5_23_i_q,
      radr => yt_rsc_5_23_i_radr,
      we => yt_rsc_5_23_we,
      d => yt_rsc_5_23_i_d,
      wadr => yt_rsc_5_23_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_5_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_5_16_i_clkr_en_d,
      d_d => yt_rsc_5_23_i_d_d,
      q_d => yt_rsc_5_23_i_q_d_1,
      radr_d => yt_rsc_5_23_i_radr_d,
      wadr_d => yt_rsc_5_23_i_wadr_d,
      we_d => yt_rsc_5_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_5_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_5_23_i_q <= yt_rsc_5_23_q;
  yt_rsc_5_23_radr <= yt_rsc_5_23_i_radr;
  yt_rsc_5_23_d <= yt_rsc_5_23_i_d;
  yt_rsc_5_23_wadr <= yt_rsc_5_23_i_wadr;
  yt_rsc_5_23_i_d_d <= yt_rsc_4_7_i_d_d_iff;
  yt_rsc_5_23_i_q_d <= yt_rsc_5_23_i_q_d_1;
  yt_rsc_5_23_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_5_23_i_wadr_d <= yt_rsc_4_0_i_wadr_d_iff;

  yt_rsc_5_24_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_191_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_5_24_clkr_en,
      clkw_en => yt_rsc_5_24_clkw_en,
      q => yt_rsc_5_24_i_q,
      radr => yt_rsc_5_24_i_radr,
      we => yt_rsc_5_24_we,
      d => yt_rsc_5_24_i_d,
      wadr => yt_rsc_5_24_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_5_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_5_16_i_clkr_en_d,
      d_d => yt_rsc_5_24_i_d_d,
      q_d => yt_rsc_5_24_i_q_d_1,
      radr_d => yt_rsc_5_24_i_radr_d,
      wadr_d => yt_rsc_5_24_i_wadr_d,
      we_d => yt_rsc_5_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_5_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_5_24_i_q <= yt_rsc_5_24_q;
  yt_rsc_5_24_radr <= yt_rsc_5_24_i_radr;
  yt_rsc_5_24_d <= yt_rsc_5_24_i_d;
  yt_rsc_5_24_wadr <= yt_rsc_5_24_i_wadr;
  yt_rsc_5_24_i_d_d <= yt_rsc_4_8_i_d_d_iff;
  yt_rsc_5_24_i_q_d <= yt_rsc_5_24_i_q_d_1;
  yt_rsc_5_24_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_5_24_i_wadr_d <= yt_rsc_4_1_i_wadr_d_iff;

  yt_rsc_5_25_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_192_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_5_25_clkr_en,
      clkw_en => yt_rsc_5_25_clkw_en,
      q => yt_rsc_5_25_i_q,
      radr => yt_rsc_5_25_i_radr,
      we => yt_rsc_5_25_we,
      d => yt_rsc_5_25_i_d,
      wadr => yt_rsc_5_25_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_5_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_5_16_i_clkr_en_d,
      d_d => yt_rsc_5_25_i_d_d,
      q_d => yt_rsc_5_25_i_q_d_1,
      radr_d => yt_rsc_5_25_i_radr_d,
      wadr_d => yt_rsc_5_25_i_wadr_d,
      we_d => yt_rsc_5_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_5_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_5_25_i_q <= yt_rsc_5_25_q;
  yt_rsc_5_25_radr <= yt_rsc_5_25_i_radr;
  yt_rsc_5_25_d <= yt_rsc_5_25_i_d;
  yt_rsc_5_25_wadr <= yt_rsc_5_25_i_wadr;
  yt_rsc_5_25_i_d_d <= yt_rsc_4_9_i_d_d_iff;
  yt_rsc_5_25_i_q_d <= yt_rsc_5_25_i_q_d_1;
  yt_rsc_5_25_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_5_25_i_wadr_d <= yt_rsc_4_9_i_wadr_d_iff;

  yt_rsc_5_26_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_193_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_5_26_clkr_en,
      clkw_en => yt_rsc_5_26_clkw_en,
      q => yt_rsc_5_26_i_q,
      radr => yt_rsc_5_26_i_radr,
      we => yt_rsc_5_26_we,
      d => yt_rsc_5_26_i_d,
      wadr => yt_rsc_5_26_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_5_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_5_16_i_clkr_en_d,
      d_d => yt_rsc_5_26_i_d_d,
      q_d => yt_rsc_5_26_i_q_d_1,
      radr_d => yt_rsc_5_26_i_radr_d,
      wadr_d => yt_rsc_5_26_i_wadr_d,
      we_d => yt_rsc_5_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_5_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_5_26_i_q <= yt_rsc_5_26_q;
  yt_rsc_5_26_radr <= yt_rsc_5_26_i_radr;
  yt_rsc_5_26_d <= yt_rsc_5_26_i_d;
  yt_rsc_5_26_wadr <= yt_rsc_5_26_i_wadr;
  yt_rsc_5_26_i_d_d <= yt_rsc_4_10_i_d_d_iff;
  yt_rsc_5_26_i_q_d <= yt_rsc_5_26_i_q_d_1;
  yt_rsc_5_26_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_5_26_i_wadr_d <= yt_rsc_4_10_i_wadr_d_iff;

  yt_rsc_5_27_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_194_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_5_27_clkr_en,
      clkw_en => yt_rsc_5_27_clkw_en,
      q => yt_rsc_5_27_i_q,
      radr => yt_rsc_5_27_i_radr,
      we => yt_rsc_5_27_we,
      d => yt_rsc_5_27_i_d,
      wadr => yt_rsc_5_27_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_5_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_5_16_i_clkr_en_d,
      d_d => yt_rsc_5_27_i_d_d,
      q_d => yt_rsc_5_27_i_q_d_1,
      radr_d => yt_rsc_5_27_i_radr_d,
      wadr_d => yt_rsc_5_27_i_wadr_d,
      we_d => yt_rsc_5_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_5_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_5_27_i_q <= yt_rsc_5_27_q;
  yt_rsc_5_27_radr <= yt_rsc_5_27_i_radr;
  yt_rsc_5_27_d <= yt_rsc_5_27_i_d;
  yt_rsc_5_27_wadr <= yt_rsc_5_27_i_wadr;
  yt_rsc_5_27_i_d_d <= yt_rsc_4_11_i_d_d_iff;
  yt_rsc_5_27_i_q_d <= yt_rsc_5_27_i_q_d_1;
  yt_rsc_5_27_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_5_27_i_wadr_d <= yt_rsc_4_11_i_wadr_d_iff;

  yt_rsc_5_28_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_195_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_5_28_clkr_en,
      clkw_en => yt_rsc_5_28_clkw_en,
      q => yt_rsc_5_28_i_q,
      radr => yt_rsc_5_28_i_radr,
      we => yt_rsc_5_28_we,
      d => yt_rsc_5_28_i_d,
      wadr => yt_rsc_5_28_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_5_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_5_16_i_clkr_en_d,
      d_d => yt_rsc_5_28_i_d_d,
      q_d => yt_rsc_5_28_i_q_d_1,
      radr_d => yt_rsc_5_28_i_radr_d,
      wadr_d => yt_rsc_5_28_i_wadr_d,
      we_d => yt_rsc_5_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_5_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_5_28_i_q <= yt_rsc_5_28_q;
  yt_rsc_5_28_radr <= yt_rsc_5_28_i_radr;
  yt_rsc_5_28_d <= yt_rsc_5_28_i_d;
  yt_rsc_5_28_wadr <= yt_rsc_5_28_i_wadr;
  yt_rsc_5_28_i_d_d <= yt_rsc_4_12_i_d_d_iff;
  yt_rsc_5_28_i_q_d <= yt_rsc_5_28_i_q_d_1;
  yt_rsc_5_28_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_5_28_i_wadr_d <= yt_rsc_4_3_i_wadr_d_iff;

  yt_rsc_5_29_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_196_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_5_29_clkr_en,
      clkw_en => yt_rsc_5_29_clkw_en,
      q => yt_rsc_5_29_i_q,
      radr => yt_rsc_5_29_i_radr,
      we => yt_rsc_5_29_we,
      d => yt_rsc_5_29_i_d,
      wadr => yt_rsc_5_29_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_5_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_5_16_i_clkr_en_d,
      d_d => yt_rsc_5_29_i_d_d,
      q_d => yt_rsc_5_29_i_q_d_1,
      radr_d => yt_rsc_5_29_i_radr_d,
      wadr_d => yt_rsc_5_29_i_wadr_d,
      we_d => yt_rsc_5_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_5_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_5_29_i_q <= yt_rsc_5_29_q;
  yt_rsc_5_29_radr <= yt_rsc_5_29_i_radr;
  yt_rsc_5_29_d <= yt_rsc_5_29_i_d;
  yt_rsc_5_29_wadr <= yt_rsc_5_29_i_wadr;
  yt_rsc_5_29_i_d_d <= yt_rsc_4_13_i_d_d_iff;
  yt_rsc_5_29_i_q_d <= yt_rsc_5_29_i_q_d_1;
  yt_rsc_5_29_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_5_29_i_wadr_d <= yt_rsc_4_4_i_wadr_d_iff;

  yt_rsc_5_30_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_197_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_5_30_clkr_en,
      clkw_en => yt_rsc_5_30_clkw_en,
      q => yt_rsc_5_30_i_q,
      radr => yt_rsc_5_30_i_radr,
      we => yt_rsc_5_30_we,
      d => yt_rsc_5_30_i_d,
      wadr => yt_rsc_5_30_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_5_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_5_16_i_clkr_en_d,
      d_d => yt_rsc_5_30_i_d_d,
      q_d => yt_rsc_5_30_i_q_d_1,
      radr_d => yt_rsc_5_30_i_radr_d,
      wadr_d => yt_rsc_5_30_i_wadr_d,
      we_d => yt_rsc_5_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_5_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_5_30_i_q <= yt_rsc_5_30_q;
  yt_rsc_5_30_radr <= yt_rsc_5_30_i_radr;
  yt_rsc_5_30_d <= yt_rsc_5_30_i_d;
  yt_rsc_5_30_wadr <= yt_rsc_5_30_i_wadr;
  yt_rsc_5_30_i_d_d <= yt_rsc_4_14_i_d_d_iff;
  yt_rsc_5_30_i_q_d <= yt_rsc_5_30_i_q_d_1;
  yt_rsc_5_30_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_5_30_i_wadr_d <= yt_rsc_4_5_i_wadr_d_iff;

  yt_rsc_5_31_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_198_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_5_31_clkr_en,
      clkw_en => yt_rsc_5_31_clkw_en,
      q => yt_rsc_5_31_i_q,
      radr => yt_rsc_5_31_i_radr,
      we => yt_rsc_5_31_we,
      d => yt_rsc_5_31_i_d,
      wadr => yt_rsc_5_31_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_5_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_5_16_i_clkr_en_d,
      d_d => yt_rsc_5_31_i_d_d,
      q_d => yt_rsc_5_31_i_q_d_1,
      radr_d => yt_rsc_5_31_i_radr_d,
      wadr_d => yt_rsc_5_31_i_wadr_d,
      we_d => yt_rsc_5_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_5_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_5_31_i_q <= yt_rsc_5_31_q;
  yt_rsc_5_31_radr <= yt_rsc_5_31_i_radr;
  yt_rsc_5_31_d <= yt_rsc_5_31_i_d;
  yt_rsc_5_31_wadr <= yt_rsc_5_31_i_wadr;
  yt_rsc_5_31_i_d_d <= yt_rsc_4_15_i_d_d_iff;
  yt_rsc_5_31_i_q_d <= yt_rsc_5_31_i_q_d_1;
  yt_rsc_5_31_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_5_31_i_wadr_d <= yt_rsc_4_6_i_wadr_d_iff;

  yt_rsc_6_0_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_199_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_6_0_clkr_en,
      clkw_en => yt_rsc_6_0_clkw_en,
      q => yt_rsc_6_0_i_q,
      radr => yt_rsc_6_0_i_radr,
      we => yt_rsc_6_0_we,
      d => yt_rsc_6_0_i_d,
      wadr => yt_rsc_6_0_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_6_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_6_0_i_clkr_en_d,
      d_d => yt_rsc_6_0_i_d_d,
      q_d => yt_rsc_6_0_i_q_d_1,
      radr_d => yt_rsc_6_0_i_radr_d,
      wadr_d => yt_rsc_6_0_i_wadr_d,
      we_d => yt_rsc_6_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_6_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_6_0_i_q <= yt_rsc_6_0_q;
  yt_rsc_6_0_radr <= yt_rsc_6_0_i_radr;
  yt_rsc_6_0_d <= yt_rsc_6_0_i_d;
  yt_rsc_6_0_wadr <= yt_rsc_6_0_i_wadr;
  yt_rsc_6_0_i_d_d <= yt_rsc_4_0_i_d_d_iff;
  yt_rsc_6_0_i_q_d <= yt_rsc_6_0_i_q_d_1;
  yt_rsc_6_0_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_6_0_i_wadr_d <= yt_rsc_4_0_i_wadr_d_iff;

  yt_rsc_6_1_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_200_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_6_1_clkr_en,
      clkw_en => yt_rsc_6_1_clkw_en,
      q => yt_rsc_6_1_i_q,
      radr => yt_rsc_6_1_i_radr,
      we => yt_rsc_6_1_we,
      d => yt_rsc_6_1_i_d,
      wadr => yt_rsc_6_1_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_6_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_6_0_i_clkr_en_d,
      d_d => yt_rsc_6_1_i_d_d,
      q_d => yt_rsc_6_1_i_q_d_1,
      radr_d => yt_rsc_6_1_i_radr_d,
      wadr_d => yt_rsc_6_1_i_wadr_d,
      we_d => yt_rsc_6_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_6_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_6_1_i_q <= yt_rsc_6_1_q;
  yt_rsc_6_1_radr <= yt_rsc_6_1_i_radr;
  yt_rsc_6_1_d <= yt_rsc_6_1_i_d;
  yt_rsc_6_1_wadr <= yt_rsc_6_1_i_wadr;
  yt_rsc_6_1_i_d_d <= yt_rsc_4_1_i_d_d_iff;
  yt_rsc_6_1_i_q_d <= yt_rsc_6_1_i_q_d_1;
  yt_rsc_6_1_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_6_1_i_wadr_d <= yt_rsc_4_1_i_wadr_d_iff;

  yt_rsc_6_2_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_201_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_6_2_clkr_en,
      clkw_en => yt_rsc_6_2_clkw_en,
      q => yt_rsc_6_2_i_q,
      radr => yt_rsc_6_2_i_radr,
      we => yt_rsc_6_2_we,
      d => yt_rsc_6_2_i_d,
      wadr => yt_rsc_6_2_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_6_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_6_0_i_clkr_en_d,
      d_d => yt_rsc_6_2_i_d_d,
      q_d => yt_rsc_6_2_i_q_d_1,
      radr_d => yt_rsc_6_2_i_radr_d,
      wadr_d => yt_rsc_6_2_i_wadr_d,
      we_d => yt_rsc_6_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_6_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_6_2_i_q <= yt_rsc_6_2_q;
  yt_rsc_6_2_radr <= yt_rsc_6_2_i_radr;
  yt_rsc_6_2_d <= yt_rsc_6_2_i_d;
  yt_rsc_6_2_wadr <= yt_rsc_6_2_i_wadr;
  yt_rsc_6_2_i_d_d <= yt_rsc_4_2_i_d_d_iff;
  yt_rsc_6_2_i_q_d <= yt_rsc_6_2_i_q_d_1;
  yt_rsc_6_2_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_6_2_i_wadr_d <= yt_rsc_4_2_i_wadr_d_iff;

  yt_rsc_6_3_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_202_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_6_3_clkr_en,
      clkw_en => yt_rsc_6_3_clkw_en,
      q => yt_rsc_6_3_i_q,
      radr => yt_rsc_6_3_i_radr,
      we => yt_rsc_6_3_we,
      d => yt_rsc_6_3_i_d,
      wadr => yt_rsc_6_3_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_6_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_6_0_i_clkr_en_d,
      d_d => yt_rsc_6_3_i_d_d,
      q_d => yt_rsc_6_3_i_q_d_1,
      radr_d => yt_rsc_6_3_i_radr_d,
      wadr_d => yt_rsc_6_3_i_wadr_d,
      we_d => yt_rsc_6_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_6_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_6_3_i_q <= yt_rsc_6_3_q;
  yt_rsc_6_3_radr <= yt_rsc_6_3_i_radr;
  yt_rsc_6_3_d <= yt_rsc_6_3_i_d;
  yt_rsc_6_3_wadr <= yt_rsc_6_3_i_wadr;
  yt_rsc_6_3_i_d_d <= yt_rsc_4_3_i_d_d_iff;
  yt_rsc_6_3_i_q_d <= yt_rsc_6_3_i_q_d_1;
  yt_rsc_6_3_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_6_3_i_wadr_d <= yt_rsc_4_3_i_wadr_d_iff;

  yt_rsc_6_4_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_203_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_6_4_clkr_en,
      clkw_en => yt_rsc_6_4_clkw_en,
      q => yt_rsc_6_4_i_q,
      radr => yt_rsc_6_4_i_radr,
      we => yt_rsc_6_4_we,
      d => yt_rsc_6_4_i_d,
      wadr => yt_rsc_6_4_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_6_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_6_0_i_clkr_en_d,
      d_d => yt_rsc_6_4_i_d_d,
      q_d => yt_rsc_6_4_i_q_d_1,
      radr_d => yt_rsc_6_4_i_radr_d,
      wadr_d => yt_rsc_6_4_i_wadr_d,
      we_d => yt_rsc_6_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_6_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_6_4_i_q <= yt_rsc_6_4_q;
  yt_rsc_6_4_radr <= yt_rsc_6_4_i_radr;
  yt_rsc_6_4_d <= yt_rsc_6_4_i_d;
  yt_rsc_6_4_wadr <= yt_rsc_6_4_i_wadr;
  yt_rsc_6_4_i_d_d <= yt_rsc_4_4_i_d_d_iff;
  yt_rsc_6_4_i_q_d <= yt_rsc_6_4_i_q_d_1;
  yt_rsc_6_4_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_6_4_i_wadr_d <= yt_rsc_4_4_i_wadr_d_iff;

  yt_rsc_6_5_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_204_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_6_5_clkr_en,
      clkw_en => yt_rsc_6_5_clkw_en,
      q => yt_rsc_6_5_i_q,
      radr => yt_rsc_6_5_i_radr,
      we => yt_rsc_6_5_we,
      d => yt_rsc_6_5_i_d,
      wadr => yt_rsc_6_5_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_6_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_6_0_i_clkr_en_d,
      d_d => yt_rsc_6_5_i_d_d,
      q_d => yt_rsc_6_5_i_q_d_1,
      radr_d => yt_rsc_6_5_i_radr_d,
      wadr_d => yt_rsc_6_5_i_wadr_d,
      we_d => yt_rsc_6_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_6_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_6_5_i_q <= yt_rsc_6_5_q;
  yt_rsc_6_5_radr <= yt_rsc_6_5_i_radr;
  yt_rsc_6_5_d <= yt_rsc_6_5_i_d;
  yt_rsc_6_5_wadr <= yt_rsc_6_5_i_wadr;
  yt_rsc_6_5_i_d_d <= yt_rsc_4_5_i_d_d_iff;
  yt_rsc_6_5_i_q_d <= yt_rsc_6_5_i_q_d_1;
  yt_rsc_6_5_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_6_5_i_wadr_d <= yt_rsc_4_5_i_wadr_d_iff;

  yt_rsc_6_6_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_205_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_6_6_clkr_en,
      clkw_en => yt_rsc_6_6_clkw_en,
      q => yt_rsc_6_6_i_q,
      radr => yt_rsc_6_6_i_radr,
      we => yt_rsc_6_6_we,
      d => yt_rsc_6_6_i_d,
      wadr => yt_rsc_6_6_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_6_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_6_0_i_clkr_en_d,
      d_d => yt_rsc_6_6_i_d_d,
      q_d => yt_rsc_6_6_i_q_d_1,
      radr_d => yt_rsc_6_6_i_radr_d,
      wadr_d => yt_rsc_6_6_i_wadr_d,
      we_d => yt_rsc_6_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_6_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_6_6_i_q <= yt_rsc_6_6_q;
  yt_rsc_6_6_radr <= yt_rsc_6_6_i_radr;
  yt_rsc_6_6_d <= yt_rsc_6_6_i_d;
  yt_rsc_6_6_wadr <= yt_rsc_6_6_i_wadr;
  yt_rsc_6_6_i_d_d <= yt_rsc_4_6_i_d_d_iff;
  yt_rsc_6_6_i_q_d <= yt_rsc_6_6_i_q_d_1;
  yt_rsc_6_6_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_6_6_i_wadr_d <= yt_rsc_4_6_i_wadr_d_iff;

  yt_rsc_6_7_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_206_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_6_7_clkr_en,
      clkw_en => yt_rsc_6_7_clkw_en,
      q => yt_rsc_6_7_i_q,
      radr => yt_rsc_6_7_i_radr,
      we => yt_rsc_6_7_we,
      d => yt_rsc_6_7_i_d,
      wadr => yt_rsc_6_7_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_6_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_6_0_i_clkr_en_d,
      d_d => yt_rsc_6_7_i_d_d,
      q_d => yt_rsc_6_7_i_q_d_1,
      radr_d => yt_rsc_6_7_i_radr_d,
      wadr_d => yt_rsc_6_7_i_wadr_d,
      we_d => yt_rsc_6_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_6_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_6_7_i_q <= yt_rsc_6_7_q;
  yt_rsc_6_7_radr <= yt_rsc_6_7_i_radr;
  yt_rsc_6_7_d <= yt_rsc_6_7_i_d;
  yt_rsc_6_7_wadr <= yt_rsc_6_7_i_wadr;
  yt_rsc_6_7_i_d_d <= yt_rsc_4_7_i_d_d_iff;
  yt_rsc_6_7_i_q_d <= yt_rsc_6_7_i_q_d_1;
  yt_rsc_6_7_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_6_7_i_wadr_d <= yt_rsc_4_0_i_wadr_d_iff;

  yt_rsc_6_8_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_207_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_6_8_clkr_en,
      clkw_en => yt_rsc_6_8_clkw_en,
      q => yt_rsc_6_8_i_q,
      radr => yt_rsc_6_8_i_radr,
      we => yt_rsc_6_8_we,
      d => yt_rsc_6_8_i_d,
      wadr => yt_rsc_6_8_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_6_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_6_0_i_clkr_en_d,
      d_d => yt_rsc_6_8_i_d_d,
      q_d => yt_rsc_6_8_i_q_d_1,
      radr_d => yt_rsc_6_8_i_radr_d,
      wadr_d => yt_rsc_6_8_i_wadr_d,
      we_d => yt_rsc_6_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_6_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_6_8_i_q <= yt_rsc_6_8_q;
  yt_rsc_6_8_radr <= yt_rsc_6_8_i_radr;
  yt_rsc_6_8_d <= yt_rsc_6_8_i_d;
  yt_rsc_6_8_wadr <= yt_rsc_6_8_i_wadr;
  yt_rsc_6_8_i_d_d <= yt_rsc_4_8_i_d_d_iff;
  yt_rsc_6_8_i_q_d <= yt_rsc_6_8_i_q_d_1;
  yt_rsc_6_8_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_6_8_i_wadr_d <= yt_rsc_4_1_i_wadr_d_iff;

  yt_rsc_6_9_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_208_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_6_9_clkr_en,
      clkw_en => yt_rsc_6_9_clkw_en,
      q => yt_rsc_6_9_i_q,
      radr => yt_rsc_6_9_i_radr,
      we => yt_rsc_6_9_we,
      d => yt_rsc_6_9_i_d,
      wadr => yt_rsc_6_9_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_6_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_6_0_i_clkr_en_d,
      d_d => yt_rsc_6_9_i_d_d,
      q_d => yt_rsc_6_9_i_q_d_1,
      radr_d => yt_rsc_6_9_i_radr_d,
      wadr_d => yt_rsc_6_9_i_wadr_d,
      we_d => yt_rsc_6_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_6_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_6_9_i_q <= yt_rsc_6_9_q;
  yt_rsc_6_9_radr <= yt_rsc_6_9_i_radr;
  yt_rsc_6_9_d <= yt_rsc_6_9_i_d;
  yt_rsc_6_9_wadr <= yt_rsc_6_9_i_wadr;
  yt_rsc_6_9_i_d_d <= yt_rsc_4_9_i_d_d_iff;
  yt_rsc_6_9_i_q_d <= yt_rsc_6_9_i_q_d_1;
  yt_rsc_6_9_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_6_9_i_wadr_d <= yt_rsc_4_9_i_wadr_d_iff;

  yt_rsc_6_10_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_209_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_6_10_clkr_en,
      clkw_en => yt_rsc_6_10_clkw_en,
      q => yt_rsc_6_10_i_q,
      radr => yt_rsc_6_10_i_radr,
      we => yt_rsc_6_10_we,
      d => yt_rsc_6_10_i_d,
      wadr => yt_rsc_6_10_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_6_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_6_0_i_clkr_en_d,
      d_d => yt_rsc_6_10_i_d_d,
      q_d => yt_rsc_6_10_i_q_d_1,
      radr_d => yt_rsc_6_10_i_radr_d,
      wadr_d => yt_rsc_6_10_i_wadr_d,
      we_d => yt_rsc_6_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_6_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_6_10_i_q <= yt_rsc_6_10_q;
  yt_rsc_6_10_radr <= yt_rsc_6_10_i_radr;
  yt_rsc_6_10_d <= yt_rsc_6_10_i_d;
  yt_rsc_6_10_wadr <= yt_rsc_6_10_i_wadr;
  yt_rsc_6_10_i_d_d <= yt_rsc_4_10_i_d_d_iff;
  yt_rsc_6_10_i_q_d <= yt_rsc_6_10_i_q_d_1;
  yt_rsc_6_10_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_6_10_i_wadr_d <= yt_rsc_4_10_i_wadr_d_iff;

  yt_rsc_6_11_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_210_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_6_11_clkr_en,
      clkw_en => yt_rsc_6_11_clkw_en,
      q => yt_rsc_6_11_i_q,
      radr => yt_rsc_6_11_i_radr,
      we => yt_rsc_6_11_we,
      d => yt_rsc_6_11_i_d,
      wadr => yt_rsc_6_11_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_6_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_6_0_i_clkr_en_d,
      d_d => yt_rsc_6_11_i_d_d,
      q_d => yt_rsc_6_11_i_q_d_1,
      radr_d => yt_rsc_6_11_i_radr_d,
      wadr_d => yt_rsc_6_11_i_wadr_d,
      we_d => yt_rsc_6_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_6_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_6_11_i_q <= yt_rsc_6_11_q;
  yt_rsc_6_11_radr <= yt_rsc_6_11_i_radr;
  yt_rsc_6_11_d <= yt_rsc_6_11_i_d;
  yt_rsc_6_11_wadr <= yt_rsc_6_11_i_wadr;
  yt_rsc_6_11_i_d_d <= yt_rsc_4_11_i_d_d_iff;
  yt_rsc_6_11_i_q_d <= yt_rsc_6_11_i_q_d_1;
  yt_rsc_6_11_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_6_11_i_wadr_d <= yt_rsc_4_11_i_wadr_d_iff;

  yt_rsc_6_12_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_211_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_6_12_clkr_en,
      clkw_en => yt_rsc_6_12_clkw_en,
      q => yt_rsc_6_12_i_q,
      radr => yt_rsc_6_12_i_radr,
      we => yt_rsc_6_12_we,
      d => yt_rsc_6_12_i_d,
      wadr => yt_rsc_6_12_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_6_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_6_0_i_clkr_en_d,
      d_d => yt_rsc_6_12_i_d_d,
      q_d => yt_rsc_6_12_i_q_d_1,
      radr_d => yt_rsc_6_12_i_radr_d,
      wadr_d => yt_rsc_6_12_i_wadr_d,
      we_d => yt_rsc_6_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_6_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_6_12_i_q <= yt_rsc_6_12_q;
  yt_rsc_6_12_radr <= yt_rsc_6_12_i_radr;
  yt_rsc_6_12_d <= yt_rsc_6_12_i_d;
  yt_rsc_6_12_wadr <= yt_rsc_6_12_i_wadr;
  yt_rsc_6_12_i_d_d <= yt_rsc_4_12_i_d_d_iff;
  yt_rsc_6_12_i_q_d <= yt_rsc_6_12_i_q_d_1;
  yt_rsc_6_12_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_6_12_i_wadr_d <= yt_rsc_4_3_i_wadr_d_iff;

  yt_rsc_6_13_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_212_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_6_13_clkr_en,
      clkw_en => yt_rsc_6_13_clkw_en,
      q => yt_rsc_6_13_i_q,
      radr => yt_rsc_6_13_i_radr,
      we => yt_rsc_6_13_we,
      d => yt_rsc_6_13_i_d,
      wadr => yt_rsc_6_13_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_6_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_6_0_i_clkr_en_d,
      d_d => yt_rsc_6_13_i_d_d,
      q_d => yt_rsc_6_13_i_q_d_1,
      radr_d => yt_rsc_6_13_i_radr_d,
      wadr_d => yt_rsc_6_13_i_wadr_d,
      we_d => yt_rsc_6_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_6_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_6_13_i_q <= yt_rsc_6_13_q;
  yt_rsc_6_13_radr <= yt_rsc_6_13_i_radr;
  yt_rsc_6_13_d <= yt_rsc_6_13_i_d;
  yt_rsc_6_13_wadr <= yt_rsc_6_13_i_wadr;
  yt_rsc_6_13_i_d_d <= yt_rsc_4_13_i_d_d_iff;
  yt_rsc_6_13_i_q_d <= yt_rsc_6_13_i_q_d_1;
  yt_rsc_6_13_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_6_13_i_wadr_d <= yt_rsc_4_4_i_wadr_d_iff;

  yt_rsc_6_14_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_213_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_6_14_clkr_en,
      clkw_en => yt_rsc_6_14_clkw_en,
      q => yt_rsc_6_14_i_q,
      radr => yt_rsc_6_14_i_radr,
      we => yt_rsc_6_14_we,
      d => yt_rsc_6_14_i_d,
      wadr => yt_rsc_6_14_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_6_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_6_0_i_clkr_en_d,
      d_d => yt_rsc_6_14_i_d_d,
      q_d => yt_rsc_6_14_i_q_d_1,
      radr_d => yt_rsc_6_14_i_radr_d,
      wadr_d => yt_rsc_6_14_i_wadr_d,
      we_d => yt_rsc_6_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_6_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_6_14_i_q <= yt_rsc_6_14_q;
  yt_rsc_6_14_radr <= yt_rsc_6_14_i_radr;
  yt_rsc_6_14_d <= yt_rsc_6_14_i_d;
  yt_rsc_6_14_wadr <= yt_rsc_6_14_i_wadr;
  yt_rsc_6_14_i_d_d <= yt_rsc_4_14_i_d_d_iff;
  yt_rsc_6_14_i_q_d <= yt_rsc_6_14_i_q_d_1;
  yt_rsc_6_14_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_6_14_i_wadr_d <= yt_rsc_4_5_i_wadr_d_iff;

  yt_rsc_6_15_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_214_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_6_15_clkr_en,
      clkw_en => yt_rsc_6_15_clkw_en,
      q => yt_rsc_6_15_i_q,
      radr => yt_rsc_6_15_i_radr,
      we => yt_rsc_6_15_we,
      d => yt_rsc_6_15_i_d,
      wadr => yt_rsc_6_15_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_6_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_6_0_i_clkr_en_d,
      d_d => yt_rsc_6_15_i_d_d,
      q_d => yt_rsc_6_15_i_q_d_1,
      radr_d => yt_rsc_6_15_i_radr_d,
      wadr_d => yt_rsc_6_15_i_wadr_d,
      we_d => yt_rsc_6_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_6_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_6_15_i_q <= yt_rsc_6_15_q;
  yt_rsc_6_15_radr <= yt_rsc_6_15_i_radr;
  yt_rsc_6_15_d <= yt_rsc_6_15_i_d;
  yt_rsc_6_15_wadr <= yt_rsc_6_15_i_wadr;
  yt_rsc_6_15_i_d_d <= yt_rsc_4_15_i_d_d_iff;
  yt_rsc_6_15_i_q_d <= yt_rsc_6_15_i_q_d_1;
  yt_rsc_6_15_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_6_15_i_wadr_d <= yt_rsc_4_6_i_wadr_d_iff;

  yt_rsc_6_16_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_215_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_6_16_clkr_en,
      clkw_en => yt_rsc_6_16_clkw_en,
      q => yt_rsc_6_16_i_q,
      radr => yt_rsc_6_16_i_radr,
      we => yt_rsc_6_16_we,
      d => yt_rsc_6_16_i_d,
      wadr => yt_rsc_6_16_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_6_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_6_16_i_clkr_en_d,
      d_d => yt_rsc_6_16_i_d_d,
      q_d => yt_rsc_6_16_i_q_d_1,
      radr_d => yt_rsc_6_16_i_radr_d,
      wadr_d => yt_rsc_6_16_i_wadr_d,
      we_d => yt_rsc_6_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_6_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_6_16_i_q <= yt_rsc_6_16_q;
  yt_rsc_6_16_radr <= yt_rsc_6_16_i_radr;
  yt_rsc_6_16_d <= yt_rsc_6_16_i_d;
  yt_rsc_6_16_wadr <= yt_rsc_6_16_i_wadr;
  yt_rsc_6_16_i_d_d <= yt_rsc_4_0_i_d_d_iff;
  yt_rsc_6_16_i_q_d <= yt_rsc_6_16_i_q_d_1;
  yt_rsc_6_16_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_6_16_i_wadr_d <= yt_rsc_4_0_i_wadr_d_iff;

  yt_rsc_6_17_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_216_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_6_17_clkr_en,
      clkw_en => yt_rsc_6_17_clkw_en,
      q => yt_rsc_6_17_i_q,
      radr => yt_rsc_6_17_i_radr,
      we => yt_rsc_6_17_we,
      d => yt_rsc_6_17_i_d,
      wadr => yt_rsc_6_17_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_6_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_6_16_i_clkr_en_d,
      d_d => yt_rsc_6_17_i_d_d,
      q_d => yt_rsc_6_17_i_q_d_1,
      radr_d => yt_rsc_6_17_i_radr_d,
      wadr_d => yt_rsc_6_17_i_wadr_d,
      we_d => yt_rsc_6_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_6_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_6_17_i_q <= yt_rsc_6_17_q;
  yt_rsc_6_17_radr <= yt_rsc_6_17_i_radr;
  yt_rsc_6_17_d <= yt_rsc_6_17_i_d;
  yt_rsc_6_17_wadr <= yt_rsc_6_17_i_wadr;
  yt_rsc_6_17_i_d_d <= yt_rsc_4_1_i_d_d_iff;
  yt_rsc_6_17_i_q_d <= yt_rsc_6_17_i_q_d_1;
  yt_rsc_6_17_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_6_17_i_wadr_d <= yt_rsc_4_1_i_wadr_d_iff;

  yt_rsc_6_18_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_217_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_6_18_clkr_en,
      clkw_en => yt_rsc_6_18_clkw_en,
      q => yt_rsc_6_18_i_q,
      radr => yt_rsc_6_18_i_radr,
      we => yt_rsc_6_18_we,
      d => yt_rsc_6_18_i_d,
      wadr => yt_rsc_6_18_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_6_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_6_16_i_clkr_en_d,
      d_d => yt_rsc_6_18_i_d_d,
      q_d => yt_rsc_6_18_i_q_d_1,
      radr_d => yt_rsc_6_18_i_radr_d,
      wadr_d => yt_rsc_6_18_i_wadr_d,
      we_d => yt_rsc_6_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_6_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_6_18_i_q <= yt_rsc_6_18_q;
  yt_rsc_6_18_radr <= yt_rsc_6_18_i_radr;
  yt_rsc_6_18_d <= yt_rsc_6_18_i_d;
  yt_rsc_6_18_wadr <= yt_rsc_6_18_i_wadr;
  yt_rsc_6_18_i_d_d <= yt_rsc_4_2_i_d_d_iff;
  yt_rsc_6_18_i_q_d <= yt_rsc_6_18_i_q_d_1;
  yt_rsc_6_18_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_6_18_i_wadr_d <= yt_rsc_4_2_i_wadr_d_iff;

  yt_rsc_6_19_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_218_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_6_19_clkr_en,
      clkw_en => yt_rsc_6_19_clkw_en,
      q => yt_rsc_6_19_i_q,
      radr => yt_rsc_6_19_i_radr,
      we => yt_rsc_6_19_we,
      d => yt_rsc_6_19_i_d,
      wadr => yt_rsc_6_19_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_6_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_6_16_i_clkr_en_d,
      d_d => yt_rsc_6_19_i_d_d,
      q_d => yt_rsc_6_19_i_q_d_1,
      radr_d => yt_rsc_6_19_i_radr_d,
      wadr_d => yt_rsc_6_19_i_wadr_d,
      we_d => yt_rsc_6_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_6_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_6_19_i_q <= yt_rsc_6_19_q;
  yt_rsc_6_19_radr <= yt_rsc_6_19_i_radr;
  yt_rsc_6_19_d <= yt_rsc_6_19_i_d;
  yt_rsc_6_19_wadr <= yt_rsc_6_19_i_wadr;
  yt_rsc_6_19_i_d_d <= yt_rsc_4_3_i_d_d_iff;
  yt_rsc_6_19_i_q_d <= yt_rsc_6_19_i_q_d_1;
  yt_rsc_6_19_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_6_19_i_wadr_d <= yt_rsc_4_3_i_wadr_d_iff;

  yt_rsc_6_20_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_219_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_6_20_clkr_en,
      clkw_en => yt_rsc_6_20_clkw_en,
      q => yt_rsc_6_20_i_q,
      radr => yt_rsc_6_20_i_radr,
      we => yt_rsc_6_20_we,
      d => yt_rsc_6_20_i_d,
      wadr => yt_rsc_6_20_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_6_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_6_16_i_clkr_en_d,
      d_d => yt_rsc_6_20_i_d_d,
      q_d => yt_rsc_6_20_i_q_d_1,
      radr_d => yt_rsc_6_20_i_radr_d,
      wadr_d => yt_rsc_6_20_i_wadr_d,
      we_d => yt_rsc_6_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_6_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_6_20_i_q <= yt_rsc_6_20_q;
  yt_rsc_6_20_radr <= yt_rsc_6_20_i_radr;
  yt_rsc_6_20_d <= yt_rsc_6_20_i_d;
  yt_rsc_6_20_wadr <= yt_rsc_6_20_i_wadr;
  yt_rsc_6_20_i_d_d <= yt_rsc_4_4_i_d_d_iff;
  yt_rsc_6_20_i_q_d <= yt_rsc_6_20_i_q_d_1;
  yt_rsc_6_20_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_6_20_i_wadr_d <= yt_rsc_4_4_i_wadr_d_iff;

  yt_rsc_6_21_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_220_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_6_21_clkr_en,
      clkw_en => yt_rsc_6_21_clkw_en,
      q => yt_rsc_6_21_i_q,
      radr => yt_rsc_6_21_i_radr,
      we => yt_rsc_6_21_we,
      d => yt_rsc_6_21_i_d,
      wadr => yt_rsc_6_21_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_6_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_6_16_i_clkr_en_d,
      d_d => yt_rsc_6_21_i_d_d,
      q_d => yt_rsc_6_21_i_q_d_1,
      radr_d => yt_rsc_6_21_i_radr_d,
      wadr_d => yt_rsc_6_21_i_wadr_d,
      we_d => yt_rsc_6_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_6_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_6_21_i_q <= yt_rsc_6_21_q;
  yt_rsc_6_21_radr <= yt_rsc_6_21_i_radr;
  yt_rsc_6_21_d <= yt_rsc_6_21_i_d;
  yt_rsc_6_21_wadr <= yt_rsc_6_21_i_wadr;
  yt_rsc_6_21_i_d_d <= yt_rsc_4_5_i_d_d_iff;
  yt_rsc_6_21_i_q_d <= yt_rsc_6_21_i_q_d_1;
  yt_rsc_6_21_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_6_21_i_wadr_d <= yt_rsc_4_5_i_wadr_d_iff;

  yt_rsc_6_22_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_221_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_6_22_clkr_en,
      clkw_en => yt_rsc_6_22_clkw_en,
      q => yt_rsc_6_22_i_q,
      radr => yt_rsc_6_22_i_radr,
      we => yt_rsc_6_22_we,
      d => yt_rsc_6_22_i_d,
      wadr => yt_rsc_6_22_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_6_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_6_16_i_clkr_en_d,
      d_d => yt_rsc_6_22_i_d_d,
      q_d => yt_rsc_6_22_i_q_d_1,
      radr_d => yt_rsc_6_22_i_radr_d,
      wadr_d => yt_rsc_6_22_i_wadr_d,
      we_d => yt_rsc_6_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_6_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_6_22_i_q <= yt_rsc_6_22_q;
  yt_rsc_6_22_radr <= yt_rsc_6_22_i_radr;
  yt_rsc_6_22_d <= yt_rsc_6_22_i_d;
  yt_rsc_6_22_wadr <= yt_rsc_6_22_i_wadr;
  yt_rsc_6_22_i_d_d <= yt_rsc_4_6_i_d_d_iff;
  yt_rsc_6_22_i_q_d <= yt_rsc_6_22_i_q_d_1;
  yt_rsc_6_22_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_6_22_i_wadr_d <= yt_rsc_4_6_i_wadr_d_iff;

  yt_rsc_6_23_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_222_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_6_23_clkr_en,
      clkw_en => yt_rsc_6_23_clkw_en,
      q => yt_rsc_6_23_i_q,
      radr => yt_rsc_6_23_i_radr,
      we => yt_rsc_6_23_we,
      d => yt_rsc_6_23_i_d,
      wadr => yt_rsc_6_23_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_6_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_6_16_i_clkr_en_d,
      d_d => yt_rsc_6_23_i_d_d,
      q_d => yt_rsc_6_23_i_q_d_1,
      radr_d => yt_rsc_6_23_i_radr_d,
      wadr_d => yt_rsc_6_23_i_wadr_d,
      we_d => yt_rsc_6_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_6_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_6_23_i_q <= yt_rsc_6_23_q;
  yt_rsc_6_23_radr <= yt_rsc_6_23_i_radr;
  yt_rsc_6_23_d <= yt_rsc_6_23_i_d;
  yt_rsc_6_23_wadr <= yt_rsc_6_23_i_wadr;
  yt_rsc_6_23_i_d_d <= yt_rsc_4_7_i_d_d_iff;
  yt_rsc_6_23_i_q_d <= yt_rsc_6_23_i_q_d_1;
  yt_rsc_6_23_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_6_23_i_wadr_d <= yt_rsc_4_0_i_wadr_d_iff;

  yt_rsc_6_24_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_223_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_6_24_clkr_en,
      clkw_en => yt_rsc_6_24_clkw_en,
      q => yt_rsc_6_24_i_q,
      radr => yt_rsc_6_24_i_radr,
      we => yt_rsc_6_24_we,
      d => yt_rsc_6_24_i_d,
      wadr => yt_rsc_6_24_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_6_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_6_16_i_clkr_en_d,
      d_d => yt_rsc_6_24_i_d_d,
      q_d => yt_rsc_6_24_i_q_d_1,
      radr_d => yt_rsc_6_24_i_radr_d,
      wadr_d => yt_rsc_6_24_i_wadr_d,
      we_d => yt_rsc_6_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_6_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_6_24_i_q <= yt_rsc_6_24_q;
  yt_rsc_6_24_radr <= yt_rsc_6_24_i_radr;
  yt_rsc_6_24_d <= yt_rsc_6_24_i_d;
  yt_rsc_6_24_wadr <= yt_rsc_6_24_i_wadr;
  yt_rsc_6_24_i_d_d <= yt_rsc_4_8_i_d_d_iff;
  yt_rsc_6_24_i_q_d <= yt_rsc_6_24_i_q_d_1;
  yt_rsc_6_24_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_6_24_i_wadr_d <= yt_rsc_4_1_i_wadr_d_iff;

  yt_rsc_6_25_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_224_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_6_25_clkr_en,
      clkw_en => yt_rsc_6_25_clkw_en,
      q => yt_rsc_6_25_i_q,
      radr => yt_rsc_6_25_i_radr,
      we => yt_rsc_6_25_we,
      d => yt_rsc_6_25_i_d,
      wadr => yt_rsc_6_25_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_6_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_6_16_i_clkr_en_d,
      d_d => yt_rsc_6_25_i_d_d,
      q_d => yt_rsc_6_25_i_q_d_1,
      radr_d => yt_rsc_6_25_i_radr_d,
      wadr_d => yt_rsc_6_25_i_wadr_d,
      we_d => yt_rsc_6_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_6_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_6_25_i_q <= yt_rsc_6_25_q;
  yt_rsc_6_25_radr <= yt_rsc_6_25_i_radr;
  yt_rsc_6_25_d <= yt_rsc_6_25_i_d;
  yt_rsc_6_25_wadr <= yt_rsc_6_25_i_wadr;
  yt_rsc_6_25_i_d_d <= yt_rsc_4_9_i_d_d_iff;
  yt_rsc_6_25_i_q_d <= yt_rsc_6_25_i_q_d_1;
  yt_rsc_6_25_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_6_25_i_wadr_d <= yt_rsc_4_9_i_wadr_d_iff;

  yt_rsc_6_26_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_225_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_6_26_clkr_en,
      clkw_en => yt_rsc_6_26_clkw_en,
      q => yt_rsc_6_26_i_q,
      radr => yt_rsc_6_26_i_radr,
      we => yt_rsc_6_26_we,
      d => yt_rsc_6_26_i_d,
      wadr => yt_rsc_6_26_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_6_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_6_16_i_clkr_en_d,
      d_d => yt_rsc_6_26_i_d_d,
      q_d => yt_rsc_6_26_i_q_d_1,
      radr_d => yt_rsc_6_26_i_radr_d,
      wadr_d => yt_rsc_6_26_i_wadr_d,
      we_d => yt_rsc_6_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_6_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_6_26_i_q <= yt_rsc_6_26_q;
  yt_rsc_6_26_radr <= yt_rsc_6_26_i_radr;
  yt_rsc_6_26_d <= yt_rsc_6_26_i_d;
  yt_rsc_6_26_wadr <= yt_rsc_6_26_i_wadr;
  yt_rsc_6_26_i_d_d <= yt_rsc_4_10_i_d_d_iff;
  yt_rsc_6_26_i_q_d <= yt_rsc_6_26_i_q_d_1;
  yt_rsc_6_26_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_6_26_i_wadr_d <= yt_rsc_4_10_i_wadr_d_iff;

  yt_rsc_6_27_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_226_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_6_27_clkr_en,
      clkw_en => yt_rsc_6_27_clkw_en,
      q => yt_rsc_6_27_i_q,
      radr => yt_rsc_6_27_i_radr,
      we => yt_rsc_6_27_we,
      d => yt_rsc_6_27_i_d,
      wadr => yt_rsc_6_27_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_6_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_6_16_i_clkr_en_d,
      d_d => yt_rsc_6_27_i_d_d,
      q_d => yt_rsc_6_27_i_q_d_1,
      radr_d => yt_rsc_6_27_i_radr_d,
      wadr_d => yt_rsc_6_27_i_wadr_d,
      we_d => yt_rsc_6_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_6_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_6_27_i_q <= yt_rsc_6_27_q;
  yt_rsc_6_27_radr <= yt_rsc_6_27_i_radr;
  yt_rsc_6_27_d <= yt_rsc_6_27_i_d;
  yt_rsc_6_27_wadr <= yt_rsc_6_27_i_wadr;
  yt_rsc_6_27_i_d_d <= yt_rsc_4_11_i_d_d_iff;
  yt_rsc_6_27_i_q_d <= yt_rsc_6_27_i_q_d_1;
  yt_rsc_6_27_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_6_27_i_wadr_d <= yt_rsc_4_11_i_wadr_d_iff;

  yt_rsc_6_28_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_227_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_6_28_clkr_en,
      clkw_en => yt_rsc_6_28_clkw_en,
      q => yt_rsc_6_28_i_q,
      radr => yt_rsc_6_28_i_radr,
      we => yt_rsc_6_28_we,
      d => yt_rsc_6_28_i_d,
      wadr => yt_rsc_6_28_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_6_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_6_16_i_clkr_en_d,
      d_d => yt_rsc_6_28_i_d_d,
      q_d => yt_rsc_6_28_i_q_d_1,
      radr_d => yt_rsc_6_28_i_radr_d,
      wadr_d => yt_rsc_6_28_i_wadr_d,
      we_d => yt_rsc_6_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_6_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_6_28_i_q <= yt_rsc_6_28_q;
  yt_rsc_6_28_radr <= yt_rsc_6_28_i_radr;
  yt_rsc_6_28_d <= yt_rsc_6_28_i_d;
  yt_rsc_6_28_wadr <= yt_rsc_6_28_i_wadr;
  yt_rsc_6_28_i_d_d <= yt_rsc_4_12_i_d_d_iff;
  yt_rsc_6_28_i_q_d <= yt_rsc_6_28_i_q_d_1;
  yt_rsc_6_28_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_6_28_i_wadr_d <= yt_rsc_4_3_i_wadr_d_iff;

  yt_rsc_6_29_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_228_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_6_29_clkr_en,
      clkw_en => yt_rsc_6_29_clkw_en,
      q => yt_rsc_6_29_i_q,
      radr => yt_rsc_6_29_i_radr,
      we => yt_rsc_6_29_we,
      d => yt_rsc_6_29_i_d,
      wadr => yt_rsc_6_29_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_6_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_6_16_i_clkr_en_d,
      d_d => yt_rsc_6_29_i_d_d,
      q_d => yt_rsc_6_29_i_q_d_1,
      radr_d => yt_rsc_6_29_i_radr_d,
      wadr_d => yt_rsc_6_29_i_wadr_d,
      we_d => yt_rsc_6_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_6_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_6_29_i_q <= yt_rsc_6_29_q;
  yt_rsc_6_29_radr <= yt_rsc_6_29_i_radr;
  yt_rsc_6_29_d <= yt_rsc_6_29_i_d;
  yt_rsc_6_29_wadr <= yt_rsc_6_29_i_wadr;
  yt_rsc_6_29_i_d_d <= yt_rsc_4_13_i_d_d_iff;
  yt_rsc_6_29_i_q_d <= yt_rsc_6_29_i_q_d_1;
  yt_rsc_6_29_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_6_29_i_wadr_d <= yt_rsc_4_4_i_wadr_d_iff;

  yt_rsc_6_30_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_229_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_6_30_clkr_en,
      clkw_en => yt_rsc_6_30_clkw_en,
      q => yt_rsc_6_30_i_q,
      radr => yt_rsc_6_30_i_radr,
      we => yt_rsc_6_30_we,
      d => yt_rsc_6_30_i_d,
      wadr => yt_rsc_6_30_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_6_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_6_16_i_clkr_en_d,
      d_d => yt_rsc_6_30_i_d_d,
      q_d => yt_rsc_6_30_i_q_d_1,
      radr_d => yt_rsc_6_30_i_radr_d,
      wadr_d => yt_rsc_6_30_i_wadr_d,
      we_d => yt_rsc_6_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_6_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_6_30_i_q <= yt_rsc_6_30_q;
  yt_rsc_6_30_radr <= yt_rsc_6_30_i_radr;
  yt_rsc_6_30_d <= yt_rsc_6_30_i_d;
  yt_rsc_6_30_wadr <= yt_rsc_6_30_i_wadr;
  yt_rsc_6_30_i_d_d <= yt_rsc_4_14_i_d_d_iff;
  yt_rsc_6_30_i_q_d <= yt_rsc_6_30_i_q_d_1;
  yt_rsc_6_30_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_6_30_i_wadr_d <= yt_rsc_4_5_i_wadr_d_iff;

  yt_rsc_6_31_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_230_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_6_31_clkr_en,
      clkw_en => yt_rsc_6_31_clkw_en,
      q => yt_rsc_6_31_i_q,
      radr => yt_rsc_6_31_i_radr,
      we => yt_rsc_6_31_we,
      d => yt_rsc_6_31_i_d,
      wadr => yt_rsc_6_31_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_6_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_6_16_i_clkr_en_d,
      d_d => yt_rsc_6_31_i_d_d,
      q_d => yt_rsc_6_31_i_q_d_1,
      radr_d => yt_rsc_6_31_i_radr_d,
      wadr_d => yt_rsc_6_31_i_wadr_d,
      we_d => yt_rsc_6_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_6_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_6_31_i_q <= yt_rsc_6_31_q;
  yt_rsc_6_31_radr <= yt_rsc_6_31_i_radr;
  yt_rsc_6_31_d <= yt_rsc_6_31_i_d;
  yt_rsc_6_31_wadr <= yt_rsc_6_31_i_wadr;
  yt_rsc_6_31_i_d_d <= yt_rsc_4_15_i_d_d_iff;
  yt_rsc_6_31_i_q_d <= yt_rsc_6_31_i_q_d_1;
  yt_rsc_6_31_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_6_31_i_wadr_d <= yt_rsc_4_6_i_wadr_d_iff;

  yt_rsc_7_0_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_231_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_7_0_clkr_en,
      clkw_en => yt_rsc_7_0_clkw_en,
      q => yt_rsc_7_0_i_q,
      radr => yt_rsc_7_0_i_radr,
      we => yt_rsc_7_0_we,
      d => yt_rsc_7_0_i_d,
      wadr => yt_rsc_7_0_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_7_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_7_0_i_clkr_en_d,
      d_d => yt_rsc_7_0_i_d_d,
      q_d => yt_rsc_7_0_i_q_d_1,
      radr_d => yt_rsc_7_0_i_radr_d,
      wadr_d => yt_rsc_7_0_i_wadr_d,
      we_d => yt_rsc_7_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_7_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_7_0_i_q <= yt_rsc_7_0_q;
  yt_rsc_7_0_radr <= yt_rsc_7_0_i_radr;
  yt_rsc_7_0_d <= yt_rsc_7_0_i_d;
  yt_rsc_7_0_wadr <= yt_rsc_7_0_i_wadr;
  yt_rsc_7_0_i_d_d <= yt_rsc_4_0_i_d_d_iff;
  yt_rsc_7_0_i_q_d <= yt_rsc_7_0_i_q_d_1;
  yt_rsc_7_0_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_7_0_i_wadr_d <= yt_rsc_4_0_i_wadr_d_iff;

  yt_rsc_7_1_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_232_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_7_1_clkr_en,
      clkw_en => yt_rsc_7_1_clkw_en,
      q => yt_rsc_7_1_i_q,
      radr => yt_rsc_7_1_i_radr,
      we => yt_rsc_7_1_we,
      d => yt_rsc_7_1_i_d,
      wadr => yt_rsc_7_1_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_7_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_7_0_i_clkr_en_d,
      d_d => yt_rsc_7_1_i_d_d,
      q_d => yt_rsc_7_1_i_q_d_1,
      radr_d => yt_rsc_7_1_i_radr_d,
      wadr_d => yt_rsc_7_1_i_wadr_d,
      we_d => yt_rsc_7_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_7_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_7_1_i_q <= yt_rsc_7_1_q;
  yt_rsc_7_1_radr <= yt_rsc_7_1_i_radr;
  yt_rsc_7_1_d <= yt_rsc_7_1_i_d;
  yt_rsc_7_1_wadr <= yt_rsc_7_1_i_wadr;
  yt_rsc_7_1_i_d_d <= yt_rsc_4_1_i_d_d_iff;
  yt_rsc_7_1_i_q_d <= yt_rsc_7_1_i_q_d_1;
  yt_rsc_7_1_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_7_1_i_wadr_d <= yt_rsc_4_1_i_wadr_d_iff;

  yt_rsc_7_2_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_233_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_7_2_clkr_en,
      clkw_en => yt_rsc_7_2_clkw_en,
      q => yt_rsc_7_2_i_q,
      radr => yt_rsc_7_2_i_radr,
      we => yt_rsc_7_2_we,
      d => yt_rsc_7_2_i_d,
      wadr => yt_rsc_7_2_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_7_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_7_0_i_clkr_en_d,
      d_d => yt_rsc_7_2_i_d_d,
      q_d => yt_rsc_7_2_i_q_d_1,
      radr_d => yt_rsc_7_2_i_radr_d,
      wadr_d => yt_rsc_7_2_i_wadr_d,
      we_d => yt_rsc_7_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_7_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_7_2_i_q <= yt_rsc_7_2_q;
  yt_rsc_7_2_radr <= yt_rsc_7_2_i_radr;
  yt_rsc_7_2_d <= yt_rsc_7_2_i_d;
  yt_rsc_7_2_wadr <= yt_rsc_7_2_i_wadr;
  yt_rsc_7_2_i_d_d <= yt_rsc_4_2_i_d_d_iff;
  yt_rsc_7_2_i_q_d <= yt_rsc_7_2_i_q_d_1;
  yt_rsc_7_2_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_7_2_i_wadr_d <= yt_rsc_4_2_i_wadr_d_iff;

  yt_rsc_7_3_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_234_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_7_3_clkr_en,
      clkw_en => yt_rsc_7_3_clkw_en,
      q => yt_rsc_7_3_i_q,
      radr => yt_rsc_7_3_i_radr,
      we => yt_rsc_7_3_we,
      d => yt_rsc_7_3_i_d,
      wadr => yt_rsc_7_3_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_7_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_7_0_i_clkr_en_d,
      d_d => yt_rsc_7_3_i_d_d,
      q_d => yt_rsc_7_3_i_q_d_1,
      radr_d => yt_rsc_7_3_i_radr_d,
      wadr_d => yt_rsc_7_3_i_wadr_d,
      we_d => yt_rsc_7_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_7_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_7_3_i_q <= yt_rsc_7_3_q;
  yt_rsc_7_3_radr <= yt_rsc_7_3_i_radr;
  yt_rsc_7_3_d <= yt_rsc_7_3_i_d;
  yt_rsc_7_3_wadr <= yt_rsc_7_3_i_wadr;
  yt_rsc_7_3_i_d_d <= yt_rsc_4_3_i_d_d_iff;
  yt_rsc_7_3_i_q_d <= yt_rsc_7_3_i_q_d_1;
  yt_rsc_7_3_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_7_3_i_wadr_d <= yt_rsc_4_3_i_wadr_d_iff;

  yt_rsc_7_4_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_235_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_7_4_clkr_en,
      clkw_en => yt_rsc_7_4_clkw_en,
      q => yt_rsc_7_4_i_q,
      radr => yt_rsc_7_4_i_radr,
      we => yt_rsc_7_4_we,
      d => yt_rsc_7_4_i_d,
      wadr => yt_rsc_7_4_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_7_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_7_0_i_clkr_en_d,
      d_d => yt_rsc_7_4_i_d_d,
      q_d => yt_rsc_7_4_i_q_d_1,
      radr_d => yt_rsc_7_4_i_radr_d,
      wadr_d => yt_rsc_7_4_i_wadr_d,
      we_d => yt_rsc_7_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_7_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_7_4_i_q <= yt_rsc_7_4_q;
  yt_rsc_7_4_radr <= yt_rsc_7_4_i_radr;
  yt_rsc_7_4_d <= yt_rsc_7_4_i_d;
  yt_rsc_7_4_wadr <= yt_rsc_7_4_i_wadr;
  yt_rsc_7_4_i_d_d <= yt_rsc_4_4_i_d_d_iff;
  yt_rsc_7_4_i_q_d <= yt_rsc_7_4_i_q_d_1;
  yt_rsc_7_4_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_7_4_i_wadr_d <= yt_rsc_4_4_i_wadr_d_iff;

  yt_rsc_7_5_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_236_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_7_5_clkr_en,
      clkw_en => yt_rsc_7_5_clkw_en,
      q => yt_rsc_7_5_i_q,
      radr => yt_rsc_7_5_i_radr,
      we => yt_rsc_7_5_we,
      d => yt_rsc_7_5_i_d,
      wadr => yt_rsc_7_5_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_7_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_7_0_i_clkr_en_d,
      d_d => yt_rsc_7_5_i_d_d,
      q_d => yt_rsc_7_5_i_q_d_1,
      radr_d => yt_rsc_7_5_i_radr_d,
      wadr_d => yt_rsc_7_5_i_wadr_d,
      we_d => yt_rsc_7_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_7_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_7_5_i_q <= yt_rsc_7_5_q;
  yt_rsc_7_5_radr <= yt_rsc_7_5_i_radr;
  yt_rsc_7_5_d <= yt_rsc_7_5_i_d;
  yt_rsc_7_5_wadr <= yt_rsc_7_5_i_wadr;
  yt_rsc_7_5_i_d_d <= yt_rsc_4_5_i_d_d_iff;
  yt_rsc_7_5_i_q_d <= yt_rsc_7_5_i_q_d_1;
  yt_rsc_7_5_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_7_5_i_wadr_d <= yt_rsc_4_5_i_wadr_d_iff;

  yt_rsc_7_6_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_237_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_7_6_clkr_en,
      clkw_en => yt_rsc_7_6_clkw_en,
      q => yt_rsc_7_6_i_q,
      radr => yt_rsc_7_6_i_radr,
      we => yt_rsc_7_6_we,
      d => yt_rsc_7_6_i_d,
      wadr => yt_rsc_7_6_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_7_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_7_0_i_clkr_en_d,
      d_d => yt_rsc_7_6_i_d_d,
      q_d => yt_rsc_7_6_i_q_d_1,
      radr_d => yt_rsc_7_6_i_radr_d,
      wadr_d => yt_rsc_7_6_i_wadr_d,
      we_d => yt_rsc_7_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_7_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_7_6_i_q <= yt_rsc_7_6_q;
  yt_rsc_7_6_radr <= yt_rsc_7_6_i_radr;
  yt_rsc_7_6_d <= yt_rsc_7_6_i_d;
  yt_rsc_7_6_wadr <= yt_rsc_7_6_i_wadr;
  yt_rsc_7_6_i_d_d <= yt_rsc_4_6_i_d_d_iff;
  yt_rsc_7_6_i_q_d <= yt_rsc_7_6_i_q_d_1;
  yt_rsc_7_6_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_7_6_i_wadr_d <= yt_rsc_4_6_i_wadr_d_iff;

  yt_rsc_7_7_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_238_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_7_7_clkr_en,
      clkw_en => yt_rsc_7_7_clkw_en,
      q => yt_rsc_7_7_i_q,
      radr => yt_rsc_7_7_i_radr,
      we => yt_rsc_7_7_we,
      d => yt_rsc_7_7_i_d,
      wadr => yt_rsc_7_7_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_7_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_7_0_i_clkr_en_d,
      d_d => yt_rsc_7_7_i_d_d,
      q_d => yt_rsc_7_7_i_q_d_1,
      radr_d => yt_rsc_7_7_i_radr_d,
      wadr_d => yt_rsc_7_7_i_wadr_d,
      we_d => yt_rsc_7_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_7_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_7_7_i_q <= yt_rsc_7_7_q;
  yt_rsc_7_7_radr <= yt_rsc_7_7_i_radr;
  yt_rsc_7_7_d <= yt_rsc_7_7_i_d;
  yt_rsc_7_7_wadr <= yt_rsc_7_7_i_wadr;
  yt_rsc_7_7_i_d_d <= yt_rsc_4_7_i_d_d_iff;
  yt_rsc_7_7_i_q_d <= yt_rsc_7_7_i_q_d_1;
  yt_rsc_7_7_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_7_7_i_wadr_d <= yt_rsc_4_0_i_wadr_d_iff;

  yt_rsc_7_8_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_239_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_7_8_clkr_en,
      clkw_en => yt_rsc_7_8_clkw_en,
      q => yt_rsc_7_8_i_q,
      radr => yt_rsc_7_8_i_radr,
      we => yt_rsc_7_8_we,
      d => yt_rsc_7_8_i_d,
      wadr => yt_rsc_7_8_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_7_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_7_0_i_clkr_en_d,
      d_d => yt_rsc_7_8_i_d_d,
      q_d => yt_rsc_7_8_i_q_d_1,
      radr_d => yt_rsc_7_8_i_radr_d,
      wadr_d => yt_rsc_7_8_i_wadr_d,
      we_d => yt_rsc_7_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_7_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_7_8_i_q <= yt_rsc_7_8_q;
  yt_rsc_7_8_radr <= yt_rsc_7_8_i_radr;
  yt_rsc_7_8_d <= yt_rsc_7_8_i_d;
  yt_rsc_7_8_wadr <= yt_rsc_7_8_i_wadr;
  yt_rsc_7_8_i_d_d <= yt_rsc_4_8_i_d_d_iff;
  yt_rsc_7_8_i_q_d <= yt_rsc_7_8_i_q_d_1;
  yt_rsc_7_8_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_7_8_i_wadr_d <= yt_rsc_4_1_i_wadr_d_iff;

  yt_rsc_7_9_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_240_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_7_9_clkr_en,
      clkw_en => yt_rsc_7_9_clkw_en,
      q => yt_rsc_7_9_i_q,
      radr => yt_rsc_7_9_i_radr,
      we => yt_rsc_7_9_we,
      d => yt_rsc_7_9_i_d,
      wadr => yt_rsc_7_9_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_7_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_7_0_i_clkr_en_d,
      d_d => yt_rsc_7_9_i_d_d,
      q_d => yt_rsc_7_9_i_q_d_1,
      radr_d => yt_rsc_7_9_i_radr_d,
      wadr_d => yt_rsc_7_9_i_wadr_d,
      we_d => yt_rsc_7_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_7_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_7_9_i_q <= yt_rsc_7_9_q;
  yt_rsc_7_9_radr <= yt_rsc_7_9_i_radr;
  yt_rsc_7_9_d <= yt_rsc_7_9_i_d;
  yt_rsc_7_9_wadr <= yt_rsc_7_9_i_wadr;
  yt_rsc_7_9_i_d_d <= yt_rsc_4_9_i_d_d_iff;
  yt_rsc_7_9_i_q_d <= yt_rsc_7_9_i_q_d_1;
  yt_rsc_7_9_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_7_9_i_wadr_d <= yt_rsc_4_9_i_wadr_d_iff;

  yt_rsc_7_10_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_241_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_7_10_clkr_en,
      clkw_en => yt_rsc_7_10_clkw_en,
      q => yt_rsc_7_10_i_q,
      radr => yt_rsc_7_10_i_radr,
      we => yt_rsc_7_10_we,
      d => yt_rsc_7_10_i_d,
      wadr => yt_rsc_7_10_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_7_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_7_0_i_clkr_en_d,
      d_d => yt_rsc_7_10_i_d_d,
      q_d => yt_rsc_7_10_i_q_d_1,
      radr_d => yt_rsc_7_10_i_radr_d,
      wadr_d => yt_rsc_7_10_i_wadr_d,
      we_d => yt_rsc_7_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_7_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_7_10_i_q <= yt_rsc_7_10_q;
  yt_rsc_7_10_radr <= yt_rsc_7_10_i_radr;
  yt_rsc_7_10_d <= yt_rsc_7_10_i_d;
  yt_rsc_7_10_wadr <= yt_rsc_7_10_i_wadr;
  yt_rsc_7_10_i_d_d <= yt_rsc_4_10_i_d_d_iff;
  yt_rsc_7_10_i_q_d <= yt_rsc_7_10_i_q_d_1;
  yt_rsc_7_10_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_7_10_i_wadr_d <= yt_rsc_4_10_i_wadr_d_iff;

  yt_rsc_7_11_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_242_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_7_11_clkr_en,
      clkw_en => yt_rsc_7_11_clkw_en,
      q => yt_rsc_7_11_i_q,
      radr => yt_rsc_7_11_i_radr,
      we => yt_rsc_7_11_we,
      d => yt_rsc_7_11_i_d,
      wadr => yt_rsc_7_11_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_7_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_7_0_i_clkr_en_d,
      d_d => yt_rsc_7_11_i_d_d,
      q_d => yt_rsc_7_11_i_q_d_1,
      radr_d => yt_rsc_7_11_i_radr_d,
      wadr_d => yt_rsc_7_11_i_wadr_d,
      we_d => yt_rsc_7_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_7_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_7_11_i_q <= yt_rsc_7_11_q;
  yt_rsc_7_11_radr <= yt_rsc_7_11_i_radr;
  yt_rsc_7_11_d <= yt_rsc_7_11_i_d;
  yt_rsc_7_11_wadr <= yt_rsc_7_11_i_wadr;
  yt_rsc_7_11_i_d_d <= yt_rsc_4_11_i_d_d_iff;
  yt_rsc_7_11_i_q_d <= yt_rsc_7_11_i_q_d_1;
  yt_rsc_7_11_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_7_11_i_wadr_d <= yt_rsc_4_11_i_wadr_d_iff;

  yt_rsc_7_12_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_243_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_7_12_clkr_en,
      clkw_en => yt_rsc_7_12_clkw_en,
      q => yt_rsc_7_12_i_q,
      radr => yt_rsc_7_12_i_radr,
      we => yt_rsc_7_12_we,
      d => yt_rsc_7_12_i_d,
      wadr => yt_rsc_7_12_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_7_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_7_0_i_clkr_en_d,
      d_d => yt_rsc_7_12_i_d_d,
      q_d => yt_rsc_7_12_i_q_d_1,
      radr_d => yt_rsc_7_12_i_radr_d,
      wadr_d => yt_rsc_7_12_i_wadr_d,
      we_d => yt_rsc_7_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_7_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_7_12_i_q <= yt_rsc_7_12_q;
  yt_rsc_7_12_radr <= yt_rsc_7_12_i_radr;
  yt_rsc_7_12_d <= yt_rsc_7_12_i_d;
  yt_rsc_7_12_wadr <= yt_rsc_7_12_i_wadr;
  yt_rsc_7_12_i_d_d <= yt_rsc_4_12_i_d_d_iff;
  yt_rsc_7_12_i_q_d <= yt_rsc_7_12_i_q_d_1;
  yt_rsc_7_12_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_7_12_i_wadr_d <= yt_rsc_4_3_i_wadr_d_iff;

  yt_rsc_7_13_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_244_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_7_13_clkr_en,
      clkw_en => yt_rsc_7_13_clkw_en,
      q => yt_rsc_7_13_i_q,
      radr => yt_rsc_7_13_i_radr,
      we => yt_rsc_7_13_we,
      d => yt_rsc_7_13_i_d,
      wadr => yt_rsc_7_13_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_7_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_7_0_i_clkr_en_d,
      d_d => yt_rsc_7_13_i_d_d,
      q_d => yt_rsc_7_13_i_q_d_1,
      radr_d => yt_rsc_7_13_i_radr_d,
      wadr_d => yt_rsc_7_13_i_wadr_d,
      we_d => yt_rsc_7_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_7_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_7_13_i_q <= yt_rsc_7_13_q;
  yt_rsc_7_13_radr <= yt_rsc_7_13_i_radr;
  yt_rsc_7_13_d <= yt_rsc_7_13_i_d;
  yt_rsc_7_13_wadr <= yt_rsc_7_13_i_wadr;
  yt_rsc_7_13_i_d_d <= yt_rsc_4_13_i_d_d_iff;
  yt_rsc_7_13_i_q_d <= yt_rsc_7_13_i_q_d_1;
  yt_rsc_7_13_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_7_13_i_wadr_d <= yt_rsc_4_4_i_wadr_d_iff;

  yt_rsc_7_14_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_245_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_7_14_clkr_en,
      clkw_en => yt_rsc_7_14_clkw_en,
      q => yt_rsc_7_14_i_q,
      radr => yt_rsc_7_14_i_radr,
      we => yt_rsc_7_14_we,
      d => yt_rsc_7_14_i_d,
      wadr => yt_rsc_7_14_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_7_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_7_0_i_clkr_en_d,
      d_d => yt_rsc_7_14_i_d_d,
      q_d => yt_rsc_7_14_i_q_d_1,
      radr_d => yt_rsc_7_14_i_radr_d,
      wadr_d => yt_rsc_7_14_i_wadr_d,
      we_d => yt_rsc_7_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_7_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_7_14_i_q <= yt_rsc_7_14_q;
  yt_rsc_7_14_radr <= yt_rsc_7_14_i_radr;
  yt_rsc_7_14_d <= yt_rsc_7_14_i_d;
  yt_rsc_7_14_wadr <= yt_rsc_7_14_i_wadr;
  yt_rsc_7_14_i_d_d <= yt_rsc_4_14_i_d_d_iff;
  yt_rsc_7_14_i_q_d <= yt_rsc_7_14_i_q_d_1;
  yt_rsc_7_14_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_7_14_i_wadr_d <= yt_rsc_4_5_i_wadr_d_iff;

  yt_rsc_7_15_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_246_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_7_15_clkr_en,
      clkw_en => yt_rsc_7_15_clkw_en,
      q => yt_rsc_7_15_i_q,
      radr => yt_rsc_7_15_i_radr,
      we => yt_rsc_7_15_we,
      d => yt_rsc_7_15_i_d,
      wadr => yt_rsc_7_15_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_7_0_i_clkr_en_d,
      clkw_en_d => yt_rsc_7_0_i_clkr_en_d,
      d_d => yt_rsc_7_15_i_d_d,
      q_d => yt_rsc_7_15_i_q_d_1,
      radr_d => yt_rsc_7_15_i_radr_d,
      wadr_d => yt_rsc_7_15_i_wadr_d,
      we_d => yt_rsc_7_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_7_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_7_15_i_q <= yt_rsc_7_15_q;
  yt_rsc_7_15_radr <= yt_rsc_7_15_i_radr;
  yt_rsc_7_15_d <= yt_rsc_7_15_i_d;
  yt_rsc_7_15_wadr <= yt_rsc_7_15_i_wadr;
  yt_rsc_7_15_i_d_d <= yt_rsc_4_15_i_d_d_iff;
  yt_rsc_7_15_i_q_d <= yt_rsc_7_15_i_q_d_1;
  yt_rsc_7_15_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_7_15_i_wadr_d <= yt_rsc_4_6_i_wadr_d_iff;

  yt_rsc_7_16_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_247_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_7_16_clkr_en,
      clkw_en => yt_rsc_7_16_clkw_en,
      q => yt_rsc_7_16_i_q,
      radr => yt_rsc_7_16_i_radr,
      we => yt_rsc_7_16_we,
      d => yt_rsc_7_16_i_d,
      wadr => yt_rsc_7_16_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_7_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_7_16_i_clkr_en_d,
      d_d => yt_rsc_7_16_i_d_d,
      q_d => yt_rsc_7_16_i_q_d_1,
      radr_d => yt_rsc_7_16_i_radr_d,
      wadr_d => yt_rsc_7_16_i_wadr_d,
      we_d => yt_rsc_7_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_7_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_7_16_i_q <= yt_rsc_7_16_q;
  yt_rsc_7_16_radr <= yt_rsc_7_16_i_radr;
  yt_rsc_7_16_d <= yt_rsc_7_16_i_d;
  yt_rsc_7_16_wadr <= yt_rsc_7_16_i_wadr;
  yt_rsc_7_16_i_d_d <= yt_rsc_4_0_i_d_d_iff;
  yt_rsc_7_16_i_q_d <= yt_rsc_7_16_i_q_d_1;
  yt_rsc_7_16_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_7_16_i_wadr_d <= yt_rsc_4_0_i_wadr_d_iff;

  yt_rsc_7_17_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_248_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_7_17_clkr_en,
      clkw_en => yt_rsc_7_17_clkw_en,
      q => yt_rsc_7_17_i_q,
      radr => yt_rsc_7_17_i_radr,
      we => yt_rsc_7_17_we,
      d => yt_rsc_7_17_i_d,
      wadr => yt_rsc_7_17_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_7_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_7_16_i_clkr_en_d,
      d_d => yt_rsc_7_17_i_d_d,
      q_d => yt_rsc_7_17_i_q_d_1,
      radr_d => yt_rsc_7_17_i_radr_d,
      wadr_d => yt_rsc_7_17_i_wadr_d,
      we_d => yt_rsc_7_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_7_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_7_17_i_q <= yt_rsc_7_17_q;
  yt_rsc_7_17_radr <= yt_rsc_7_17_i_radr;
  yt_rsc_7_17_d <= yt_rsc_7_17_i_d;
  yt_rsc_7_17_wadr <= yt_rsc_7_17_i_wadr;
  yt_rsc_7_17_i_d_d <= yt_rsc_4_1_i_d_d_iff;
  yt_rsc_7_17_i_q_d <= yt_rsc_7_17_i_q_d_1;
  yt_rsc_7_17_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_7_17_i_wadr_d <= yt_rsc_4_1_i_wadr_d_iff;

  yt_rsc_7_18_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_249_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_7_18_clkr_en,
      clkw_en => yt_rsc_7_18_clkw_en,
      q => yt_rsc_7_18_i_q,
      radr => yt_rsc_7_18_i_radr,
      we => yt_rsc_7_18_we,
      d => yt_rsc_7_18_i_d,
      wadr => yt_rsc_7_18_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_7_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_7_16_i_clkr_en_d,
      d_d => yt_rsc_7_18_i_d_d,
      q_d => yt_rsc_7_18_i_q_d_1,
      radr_d => yt_rsc_7_18_i_radr_d,
      wadr_d => yt_rsc_7_18_i_wadr_d,
      we_d => yt_rsc_7_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_7_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_7_18_i_q <= yt_rsc_7_18_q;
  yt_rsc_7_18_radr <= yt_rsc_7_18_i_radr;
  yt_rsc_7_18_d <= yt_rsc_7_18_i_d;
  yt_rsc_7_18_wadr <= yt_rsc_7_18_i_wadr;
  yt_rsc_7_18_i_d_d <= yt_rsc_4_2_i_d_d_iff;
  yt_rsc_7_18_i_q_d <= yt_rsc_7_18_i_q_d_1;
  yt_rsc_7_18_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_7_18_i_wadr_d <= yt_rsc_4_2_i_wadr_d_iff;

  yt_rsc_7_19_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_250_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_7_19_clkr_en,
      clkw_en => yt_rsc_7_19_clkw_en,
      q => yt_rsc_7_19_i_q,
      radr => yt_rsc_7_19_i_radr,
      we => yt_rsc_7_19_we,
      d => yt_rsc_7_19_i_d,
      wadr => yt_rsc_7_19_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_7_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_7_16_i_clkr_en_d,
      d_d => yt_rsc_7_19_i_d_d,
      q_d => yt_rsc_7_19_i_q_d_1,
      radr_d => yt_rsc_7_19_i_radr_d,
      wadr_d => yt_rsc_7_19_i_wadr_d,
      we_d => yt_rsc_7_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_7_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_7_19_i_q <= yt_rsc_7_19_q;
  yt_rsc_7_19_radr <= yt_rsc_7_19_i_radr;
  yt_rsc_7_19_d <= yt_rsc_7_19_i_d;
  yt_rsc_7_19_wadr <= yt_rsc_7_19_i_wadr;
  yt_rsc_7_19_i_d_d <= yt_rsc_4_3_i_d_d_iff;
  yt_rsc_7_19_i_q_d <= yt_rsc_7_19_i_q_d_1;
  yt_rsc_7_19_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_7_19_i_wadr_d <= yt_rsc_4_3_i_wadr_d_iff;

  yt_rsc_7_20_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_251_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_7_20_clkr_en,
      clkw_en => yt_rsc_7_20_clkw_en,
      q => yt_rsc_7_20_i_q,
      radr => yt_rsc_7_20_i_radr,
      we => yt_rsc_7_20_we,
      d => yt_rsc_7_20_i_d,
      wadr => yt_rsc_7_20_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_7_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_7_16_i_clkr_en_d,
      d_d => yt_rsc_7_20_i_d_d,
      q_d => yt_rsc_7_20_i_q_d_1,
      radr_d => yt_rsc_7_20_i_radr_d,
      wadr_d => yt_rsc_7_20_i_wadr_d,
      we_d => yt_rsc_7_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_7_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_7_20_i_q <= yt_rsc_7_20_q;
  yt_rsc_7_20_radr <= yt_rsc_7_20_i_radr;
  yt_rsc_7_20_d <= yt_rsc_7_20_i_d;
  yt_rsc_7_20_wadr <= yt_rsc_7_20_i_wadr;
  yt_rsc_7_20_i_d_d <= yt_rsc_4_4_i_d_d_iff;
  yt_rsc_7_20_i_q_d <= yt_rsc_7_20_i_q_d_1;
  yt_rsc_7_20_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_7_20_i_wadr_d <= yt_rsc_4_4_i_wadr_d_iff;

  yt_rsc_7_21_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_252_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_7_21_clkr_en,
      clkw_en => yt_rsc_7_21_clkw_en,
      q => yt_rsc_7_21_i_q,
      radr => yt_rsc_7_21_i_radr,
      we => yt_rsc_7_21_we,
      d => yt_rsc_7_21_i_d,
      wadr => yt_rsc_7_21_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_7_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_7_16_i_clkr_en_d,
      d_d => yt_rsc_7_21_i_d_d,
      q_d => yt_rsc_7_21_i_q_d_1,
      radr_d => yt_rsc_7_21_i_radr_d,
      wadr_d => yt_rsc_7_21_i_wadr_d,
      we_d => yt_rsc_7_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_7_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_7_21_i_q <= yt_rsc_7_21_q;
  yt_rsc_7_21_radr <= yt_rsc_7_21_i_radr;
  yt_rsc_7_21_d <= yt_rsc_7_21_i_d;
  yt_rsc_7_21_wadr <= yt_rsc_7_21_i_wadr;
  yt_rsc_7_21_i_d_d <= yt_rsc_4_5_i_d_d_iff;
  yt_rsc_7_21_i_q_d <= yt_rsc_7_21_i_q_d_1;
  yt_rsc_7_21_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_7_21_i_wadr_d <= yt_rsc_4_5_i_wadr_d_iff;

  yt_rsc_7_22_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_253_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_7_22_clkr_en,
      clkw_en => yt_rsc_7_22_clkw_en,
      q => yt_rsc_7_22_i_q,
      radr => yt_rsc_7_22_i_radr,
      we => yt_rsc_7_22_we,
      d => yt_rsc_7_22_i_d,
      wadr => yt_rsc_7_22_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_7_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_7_16_i_clkr_en_d,
      d_d => yt_rsc_7_22_i_d_d,
      q_d => yt_rsc_7_22_i_q_d_1,
      radr_d => yt_rsc_7_22_i_radr_d,
      wadr_d => yt_rsc_7_22_i_wadr_d,
      we_d => yt_rsc_7_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_7_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_7_22_i_q <= yt_rsc_7_22_q;
  yt_rsc_7_22_radr <= yt_rsc_7_22_i_radr;
  yt_rsc_7_22_d <= yt_rsc_7_22_i_d;
  yt_rsc_7_22_wadr <= yt_rsc_7_22_i_wadr;
  yt_rsc_7_22_i_d_d <= yt_rsc_4_6_i_d_d_iff;
  yt_rsc_7_22_i_q_d <= yt_rsc_7_22_i_q_d_1;
  yt_rsc_7_22_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_7_22_i_wadr_d <= yt_rsc_4_6_i_wadr_d_iff;

  yt_rsc_7_23_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_254_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_7_23_clkr_en,
      clkw_en => yt_rsc_7_23_clkw_en,
      q => yt_rsc_7_23_i_q,
      radr => yt_rsc_7_23_i_radr,
      we => yt_rsc_7_23_we,
      d => yt_rsc_7_23_i_d,
      wadr => yt_rsc_7_23_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_7_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_7_16_i_clkr_en_d,
      d_d => yt_rsc_7_23_i_d_d,
      q_d => yt_rsc_7_23_i_q_d_1,
      radr_d => yt_rsc_7_23_i_radr_d,
      wadr_d => yt_rsc_7_23_i_wadr_d,
      we_d => yt_rsc_7_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_7_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_7_23_i_q <= yt_rsc_7_23_q;
  yt_rsc_7_23_radr <= yt_rsc_7_23_i_radr;
  yt_rsc_7_23_d <= yt_rsc_7_23_i_d;
  yt_rsc_7_23_wadr <= yt_rsc_7_23_i_wadr;
  yt_rsc_7_23_i_d_d <= yt_rsc_4_7_i_d_d_iff;
  yt_rsc_7_23_i_q_d <= yt_rsc_7_23_i_q_d_1;
  yt_rsc_7_23_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_7_23_i_wadr_d <= yt_rsc_4_0_i_wadr_d_iff;

  yt_rsc_7_24_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_255_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_7_24_clkr_en,
      clkw_en => yt_rsc_7_24_clkw_en,
      q => yt_rsc_7_24_i_q,
      radr => yt_rsc_7_24_i_radr,
      we => yt_rsc_7_24_we,
      d => yt_rsc_7_24_i_d,
      wadr => yt_rsc_7_24_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_7_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_7_16_i_clkr_en_d,
      d_d => yt_rsc_7_24_i_d_d,
      q_d => yt_rsc_7_24_i_q_d_1,
      radr_d => yt_rsc_7_24_i_radr_d,
      wadr_d => yt_rsc_7_24_i_wadr_d,
      we_d => yt_rsc_7_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_7_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_7_24_i_q <= yt_rsc_7_24_q;
  yt_rsc_7_24_radr <= yt_rsc_7_24_i_radr;
  yt_rsc_7_24_d <= yt_rsc_7_24_i_d;
  yt_rsc_7_24_wadr <= yt_rsc_7_24_i_wadr;
  yt_rsc_7_24_i_d_d <= yt_rsc_4_8_i_d_d_iff;
  yt_rsc_7_24_i_q_d <= yt_rsc_7_24_i_q_d_1;
  yt_rsc_7_24_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_7_24_i_wadr_d <= yt_rsc_4_1_i_wadr_d_iff;

  yt_rsc_7_25_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_256_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_7_25_clkr_en,
      clkw_en => yt_rsc_7_25_clkw_en,
      q => yt_rsc_7_25_i_q,
      radr => yt_rsc_7_25_i_radr,
      we => yt_rsc_7_25_we,
      d => yt_rsc_7_25_i_d,
      wadr => yt_rsc_7_25_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_7_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_7_16_i_clkr_en_d,
      d_d => yt_rsc_7_25_i_d_d,
      q_d => yt_rsc_7_25_i_q_d_1,
      radr_d => yt_rsc_7_25_i_radr_d,
      wadr_d => yt_rsc_7_25_i_wadr_d,
      we_d => yt_rsc_7_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_7_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_7_25_i_q <= yt_rsc_7_25_q;
  yt_rsc_7_25_radr <= yt_rsc_7_25_i_radr;
  yt_rsc_7_25_d <= yt_rsc_7_25_i_d;
  yt_rsc_7_25_wadr <= yt_rsc_7_25_i_wadr;
  yt_rsc_7_25_i_d_d <= yt_rsc_4_9_i_d_d_iff;
  yt_rsc_7_25_i_q_d <= yt_rsc_7_25_i_q_d_1;
  yt_rsc_7_25_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_7_25_i_wadr_d <= yt_rsc_4_9_i_wadr_d_iff;

  yt_rsc_7_26_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_257_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_7_26_clkr_en,
      clkw_en => yt_rsc_7_26_clkw_en,
      q => yt_rsc_7_26_i_q,
      radr => yt_rsc_7_26_i_radr,
      we => yt_rsc_7_26_we,
      d => yt_rsc_7_26_i_d,
      wadr => yt_rsc_7_26_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_7_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_7_16_i_clkr_en_d,
      d_d => yt_rsc_7_26_i_d_d,
      q_d => yt_rsc_7_26_i_q_d_1,
      radr_d => yt_rsc_7_26_i_radr_d,
      wadr_d => yt_rsc_7_26_i_wadr_d,
      we_d => yt_rsc_7_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_7_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_7_26_i_q <= yt_rsc_7_26_q;
  yt_rsc_7_26_radr <= yt_rsc_7_26_i_radr;
  yt_rsc_7_26_d <= yt_rsc_7_26_i_d;
  yt_rsc_7_26_wadr <= yt_rsc_7_26_i_wadr;
  yt_rsc_7_26_i_d_d <= yt_rsc_4_10_i_d_d_iff;
  yt_rsc_7_26_i_q_d <= yt_rsc_7_26_i_q_d_1;
  yt_rsc_7_26_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_7_26_i_wadr_d <= yt_rsc_4_10_i_wadr_d_iff;

  yt_rsc_7_27_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_258_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_7_27_clkr_en,
      clkw_en => yt_rsc_7_27_clkw_en,
      q => yt_rsc_7_27_i_q,
      radr => yt_rsc_7_27_i_radr,
      we => yt_rsc_7_27_we,
      d => yt_rsc_7_27_i_d,
      wadr => yt_rsc_7_27_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_7_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_7_16_i_clkr_en_d,
      d_d => yt_rsc_7_27_i_d_d,
      q_d => yt_rsc_7_27_i_q_d_1,
      radr_d => yt_rsc_7_27_i_radr_d,
      wadr_d => yt_rsc_7_27_i_wadr_d,
      we_d => yt_rsc_7_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_7_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_7_27_i_q <= yt_rsc_7_27_q;
  yt_rsc_7_27_radr <= yt_rsc_7_27_i_radr;
  yt_rsc_7_27_d <= yt_rsc_7_27_i_d;
  yt_rsc_7_27_wadr <= yt_rsc_7_27_i_wadr;
  yt_rsc_7_27_i_d_d <= yt_rsc_4_11_i_d_d_iff;
  yt_rsc_7_27_i_q_d <= yt_rsc_7_27_i_q_d_1;
  yt_rsc_7_27_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_7_27_i_wadr_d <= yt_rsc_4_11_i_wadr_d_iff;

  yt_rsc_7_28_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_259_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_7_28_clkr_en,
      clkw_en => yt_rsc_7_28_clkw_en,
      q => yt_rsc_7_28_i_q,
      radr => yt_rsc_7_28_i_radr,
      we => yt_rsc_7_28_we,
      d => yt_rsc_7_28_i_d,
      wadr => yt_rsc_7_28_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_7_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_7_16_i_clkr_en_d,
      d_d => yt_rsc_7_28_i_d_d,
      q_d => yt_rsc_7_28_i_q_d_1,
      radr_d => yt_rsc_7_28_i_radr_d,
      wadr_d => yt_rsc_7_28_i_wadr_d,
      we_d => yt_rsc_7_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_7_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_7_28_i_q <= yt_rsc_7_28_q;
  yt_rsc_7_28_radr <= yt_rsc_7_28_i_radr;
  yt_rsc_7_28_d <= yt_rsc_7_28_i_d;
  yt_rsc_7_28_wadr <= yt_rsc_7_28_i_wadr;
  yt_rsc_7_28_i_d_d <= yt_rsc_4_12_i_d_d_iff;
  yt_rsc_7_28_i_q_d <= yt_rsc_7_28_i_q_d_1;
  yt_rsc_7_28_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_7_28_i_wadr_d <= yt_rsc_4_3_i_wadr_d_iff;

  yt_rsc_7_29_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_260_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_7_29_clkr_en,
      clkw_en => yt_rsc_7_29_clkw_en,
      q => yt_rsc_7_29_i_q,
      radr => yt_rsc_7_29_i_radr,
      we => yt_rsc_7_29_we,
      d => yt_rsc_7_29_i_d,
      wadr => yt_rsc_7_29_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_7_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_7_16_i_clkr_en_d,
      d_d => yt_rsc_7_29_i_d_d,
      q_d => yt_rsc_7_29_i_q_d_1,
      radr_d => yt_rsc_7_29_i_radr_d,
      wadr_d => yt_rsc_7_29_i_wadr_d,
      we_d => yt_rsc_7_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_7_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_7_29_i_q <= yt_rsc_7_29_q;
  yt_rsc_7_29_radr <= yt_rsc_7_29_i_radr;
  yt_rsc_7_29_d <= yt_rsc_7_29_i_d;
  yt_rsc_7_29_wadr <= yt_rsc_7_29_i_wadr;
  yt_rsc_7_29_i_d_d <= yt_rsc_4_13_i_d_d_iff;
  yt_rsc_7_29_i_q_d <= yt_rsc_7_29_i_q_d_1;
  yt_rsc_7_29_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_7_29_i_wadr_d <= yt_rsc_4_4_i_wadr_d_iff;

  yt_rsc_7_30_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_261_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_7_30_clkr_en,
      clkw_en => yt_rsc_7_30_clkw_en,
      q => yt_rsc_7_30_i_q,
      radr => yt_rsc_7_30_i_radr,
      we => yt_rsc_7_30_we,
      d => yt_rsc_7_30_i_d,
      wadr => yt_rsc_7_30_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_7_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_7_16_i_clkr_en_d,
      d_d => yt_rsc_7_30_i_d_d,
      q_d => yt_rsc_7_30_i_q_d_1,
      radr_d => yt_rsc_7_30_i_radr_d,
      wadr_d => yt_rsc_7_30_i_wadr_d,
      we_d => yt_rsc_7_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_7_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_7_30_i_q <= yt_rsc_7_30_q;
  yt_rsc_7_30_radr <= yt_rsc_7_30_i_radr;
  yt_rsc_7_30_d <= yt_rsc_7_30_i_d;
  yt_rsc_7_30_wadr <= yt_rsc_7_30_i_wadr;
  yt_rsc_7_30_i_d_d <= yt_rsc_4_14_i_d_d_iff;
  yt_rsc_7_30_i_q_d <= yt_rsc_7_30_i_q_d_1;
  yt_rsc_7_30_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_7_30_i_wadr_d <= yt_rsc_4_5_i_wadr_d_iff;

  yt_rsc_7_31_i : peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_262_4_32_16_16_32_1_gen
    PORT MAP(
      clkr_en => yt_rsc_7_31_clkr_en,
      clkw_en => yt_rsc_7_31_clkw_en,
      q => yt_rsc_7_31_i_q,
      radr => yt_rsc_7_31_i_radr,
      we => yt_rsc_7_31_we,
      d => yt_rsc_7_31_i_d,
      wadr => yt_rsc_7_31_i_wadr,
      clkr => clk,
      clkr_en_d => yt_rsc_7_16_i_clkr_en_d,
      clkw_en_d => yt_rsc_7_16_i_clkr_en_d,
      d_d => yt_rsc_7_31_i_d_d,
      q_d => yt_rsc_7_31_i_q_d_1,
      radr_d => yt_rsc_7_31_i_radr_d,
      wadr_d => yt_rsc_7_31_i_wadr_d,
      we_d => yt_rsc_7_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => yt_rsc_7_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff
    );
  yt_rsc_7_31_i_q <= yt_rsc_7_31_q;
  yt_rsc_7_31_radr <= yt_rsc_7_31_i_radr;
  yt_rsc_7_31_d <= yt_rsc_7_31_i_d;
  yt_rsc_7_31_wadr <= yt_rsc_7_31_i_wadr;
  yt_rsc_7_31_i_d_d <= yt_rsc_4_15_i_d_d_iff;
  yt_rsc_7_31_i_q_d <= yt_rsc_7_31_i_q_d_1;
  yt_rsc_7_31_i_radr_d <= yt_rsc_0_0_i_radr_d_iff;
  yt_rsc_7_31_i_wadr_d <= yt_rsc_4_6_i_wadr_d_iff;

  xt_rsc_0_0_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_263_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_0_0_i_qa,
      wea => xt_rsc_0_0_wea,
      da => xt_rsc_0_0_i_da,
      adra => xt_rsc_0_0_i_adra,
      adra_d => xt_rsc_0_0_i_adra_d,
      da_d => xt_rsc_0_0_i_da_d,
      qa_d => xt_rsc_0_0_i_qa_d_1,
      wea_d => xt_rsc_0_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_0_i_wea_d_iff
    );
  xt_rsc_0_0_i_qa <= xt_rsc_0_0_qa;
  xt_rsc_0_0_da <= xt_rsc_0_0_i_da;
  xt_rsc_0_0_adra <= xt_rsc_0_0_i_adra;
  xt_rsc_0_0_i_adra_d <= xt_rsc_0_0_i_adra_d_iff;
  xt_rsc_0_0_i_da_d <= xt_rsc_0_0_i_da_d_iff;
  xt_rsc_0_0_i_qa_d <= xt_rsc_0_0_i_qa_d_1;

  xt_rsc_0_1_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_264_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_0_1_i_qa,
      wea => xt_rsc_0_1_wea,
      da => xt_rsc_0_1_i_da,
      adra => xt_rsc_0_1_i_adra,
      adra_d => xt_rsc_0_1_i_adra_d,
      da_d => xt_rsc_0_1_i_da_d,
      qa_d => xt_rsc_0_1_i_qa_d_1,
      wea_d => xt_rsc_0_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_0_i_wea_d_iff
    );
  xt_rsc_0_1_i_qa <= xt_rsc_0_1_qa;
  xt_rsc_0_1_da <= xt_rsc_0_1_i_da;
  xt_rsc_0_1_adra <= xt_rsc_0_1_i_adra;
  xt_rsc_0_1_i_adra_d <= xt_rsc_0_1_i_adra_d_iff;
  xt_rsc_0_1_i_da_d <= xt_rsc_0_1_i_da_d_iff;
  xt_rsc_0_1_i_qa_d <= xt_rsc_0_1_i_qa_d_1;

  xt_rsc_0_2_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_265_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_0_2_i_qa,
      wea => xt_rsc_0_2_wea,
      da => xt_rsc_0_2_i_da,
      adra => xt_rsc_0_2_i_adra,
      adra_d => xt_rsc_0_2_i_adra_d,
      da_d => xt_rsc_0_2_i_da_d,
      qa_d => xt_rsc_0_2_i_qa_d_1,
      wea_d => xt_rsc_0_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_0_i_wea_d_iff
    );
  xt_rsc_0_2_i_qa <= xt_rsc_0_2_qa;
  xt_rsc_0_2_da <= xt_rsc_0_2_i_da;
  xt_rsc_0_2_adra <= xt_rsc_0_2_i_adra;
  xt_rsc_0_2_i_adra_d <= xt_rsc_0_2_i_adra_d_iff;
  xt_rsc_0_2_i_da_d <= xt_rsc_0_2_i_da_d_iff;
  xt_rsc_0_2_i_qa_d <= xt_rsc_0_2_i_qa_d_1;

  xt_rsc_0_3_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_266_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_0_3_i_qa,
      wea => xt_rsc_0_3_wea,
      da => xt_rsc_0_3_i_da,
      adra => xt_rsc_0_3_i_adra,
      adra_d => xt_rsc_0_3_i_adra_d,
      da_d => xt_rsc_0_3_i_da_d,
      qa_d => xt_rsc_0_3_i_qa_d_1,
      wea_d => xt_rsc_0_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_0_i_wea_d_iff
    );
  xt_rsc_0_3_i_qa <= xt_rsc_0_3_qa;
  xt_rsc_0_3_da <= xt_rsc_0_3_i_da;
  xt_rsc_0_3_adra <= xt_rsc_0_3_i_adra;
  xt_rsc_0_3_i_adra_d <= xt_rsc_0_3_i_adra_d_iff;
  xt_rsc_0_3_i_da_d <= xt_rsc_0_3_i_da_d_iff;
  xt_rsc_0_3_i_qa_d <= xt_rsc_0_3_i_qa_d_1;

  xt_rsc_0_4_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_267_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_0_4_i_qa,
      wea => xt_rsc_0_4_wea,
      da => xt_rsc_0_4_i_da,
      adra => xt_rsc_0_4_i_adra,
      adra_d => xt_rsc_0_4_i_adra_d,
      da_d => xt_rsc_0_4_i_da_d,
      qa_d => xt_rsc_0_4_i_qa_d_1,
      wea_d => xt_rsc_0_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_0_i_wea_d_iff
    );
  xt_rsc_0_4_i_qa <= xt_rsc_0_4_qa;
  xt_rsc_0_4_da <= xt_rsc_0_4_i_da;
  xt_rsc_0_4_adra <= xt_rsc_0_4_i_adra;
  xt_rsc_0_4_i_adra_d <= xt_rsc_0_4_i_adra_d_iff;
  xt_rsc_0_4_i_da_d <= xt_rsc_0_4_i_da_d_iff;
  xt_rsc_0_4_i_qa_d <= xt_rsc_0_4_i_qa_d_1;

  xt_rsc_0_5_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_268_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_0_5_i_qa,
      wea => xt_rsc_0_5_wea,
      da => xt_rsc_0_5_i_da,
      adra => xt_rsc_0_5_i_adra,
      adra_d => xt_rsc_0_5_i_adra_d,
      da_d => xt_rsc_0_5_i_da_d,
      qa_d => xt_rsc_0_5_i_qa_d_1,
      wea_d => xt_rsc_0_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_0_i_wea_d_iff
    );
  xt_rsc_0_5_i_qa <= xt_rsc_0_5_qa;
  xt_rsc_0_5_da <= xt_rsc_0_5_i_da;
  xt_rsc_0_5_adra <= xt_rsc_0_5_i_adra;
  xt_rsc_0_5_i_adra_d <= xt_rsc_0_5_i_adra_d_iff;
  xt_rsc_0_5_i_da_d <= xt_rsc_0_5_i_da_d_iff;
  xt_rsc_0_5_i_qa_d <= xt_rsc_0_5_i_qa_d_1;

  xt_rsc_0_6_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_269_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_0_6_i_qa,
      wea => xt_rsc_0_6_wea,
      da => xt_rsc_0_6_i_da,
      adra => xt_rsc_0_6_i_adra,
      adra_d => xt_rsc_0_6_i_adra_d,
      da_d => xt_rsc_0_6_i_da_d,
      qa_d => xt_rsc_0_6_i_qa_d_1,
      wea_d => xt_rsc_0_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_0_i_wea_d_iff
    );
  xt_rsc_0_6_i_qa <= xt_rsc_0_6_qa;
  xt_rsc_0_6_da <= xt_rsc_0_6_i_da;
  xt_rsc_0_6_adra <= xt_rsc_0_6_i_adra;
  xt_rsc_0_6_i_adra_d <= xt_rsc_0_6_i_adra_d_iff;
  xt_rsc_0_6_i_da_d <= xt_rsc_0_6_i_da_d_iff;
  xt_rsc_0_6_i_qa_d <= xt_rsc_0_6_i_qa_d_1;

  xt_rsc_0_7_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_270_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_0_7_i_qa,
      wea => xt_rsc_0_7_wea,
      da => xt_rsc_0_7_i_da,
      adra => xt_rsc_0_7_i_adra,
      adra_d => xt_rsc_0_7_i_adra_d,
      da_d => xt_rsc_0_7_i_da_d,
      qa_d => xt_rsc_0_7_i_qa_d_1,
      wea_d => xt_rsc_0_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_0_i_wea_d_iff
    );
  xt_rsc_0_7_i_qa <= xt_rsc_0_7_qa;
  xt_rsc_0_7_da <= xt_rsc_0_7_i_da;
  xt_rsc_0_7_adra <= xt_rsc_0_7_i_adra;
  xt_rsc_0_7_i_adra_d <= xt_rsc_0_7_i_adra_d_iff;
  xt_rsc_0_7_i_da_d <= xt_rsc_0_7_i_da_d_iff;
  xt_rsc_0_7_i_qa_d <= xt_rsc_0_7_i_qa_d_1;

  xt_rsc_0_8_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_271_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_0_8_i_qa,
      wea => xt_rsc_0_8_wea,
      da => xt_rsc_0_8_i_da,
      adra => xt_rsc_0_8_i_adra,
      adra_d => xt_rsc_0_8_i_adra_d,
      da_d => xt_rsc_0_8_i_da_d,
      qa_d => xt_rsc_0_8_i_qa_d_1,
      wea_d => xt_rsc_0_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_0_i_wea_d_iff
    );
  xt_rsc_0_8_i_qa <= xt_rsc_0_8_qa;
  xt_rsc_0_8_da <= xt_rsc_0_8_i_da;
  xt_rsc_0_8_adra <= xt_rsc_0_8_i_adra;
  xt_rsc_0_8_i_adra_d <= xt_rsc_0_8_i_adra_d_iff;
  xt_rsc_0_8_i_da_d <= xt_rsc_0_8_i_da_d_iff;
  xt_rsc_0_8_i_qa_d <= xt_rsc_0_8_i_qa_d_1;

  xt_rsc_0_9_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_272_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_0_9_i_qa,
      wea => xt_rsc_0_9_wea,
      da => xt_rsc_0_9_i_da,
      adra => xt_rsc_0_9_i_adra,
      adra_d => xt_rsc_0_9_i_adra_d,
      da_d => xt_rsc_0_9_i_da_d,
      qa_d => xt_rsc_0_9_i_qa_d_1,
      wea_d => xt_rsc_0_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_0_i_wea_d_iff
    );
  xt_rsc_0_9_i_qa <= xt_rsc_0_9_qa;
  xt_rsc_0_9_da <= xt_rsc_0_9_i_da;
  xt_rsc_0_9_adra <= xt_rsc_0_9_i_adra;
  xt_rsc_0_9_i_adra_d <= xt_rsc_0_9_i_adra_d_iff;
  xt_rsc_0_9_i_da_d <= xt_rsc_0_9_i_da_d_iff;
  xt_rsc_0_9_i_qa_d <= xt_rsc_0_9_i_qa_d_1;

  xt_rsc_0_10_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_273_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_0_10_i_qa,
      wea => xt_rsc_0_10_wea,
      da => xt_rsc_0_10_i_da,
      adra => xt_rsc_0_10_i_adra,
      adra_d => xt_rsc_0_10_i_adra_d,
      da_d => xt_rsc_0_10_i_da_d,
      qa_d => xt_rsc_0_10_i_qa_d_1,
      wea_d => xt_rsc_0_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_0_i_wea_d_iff
    );
  xt_rsc_0_10_i_qa <= xt_rsc_0_10_qa;
  xt_rsc_0_10_da <= xt_rsc_0_10_i_da;
  xt_rsc_0_10_adra <= xt_rsc_0_10_i_adra;
  xt_rsc_0_10_i_adra_d <= xt_rsc_0_10_i_adra_d_iff;
  xt_rsc_0_10_i_da_d <= xt_rsc_0_10_i_da_d_iff;
  xt_rsc_0_10_i_qa_d <= xt_rsc_0_10_i_qa_d_1;

  xt_rsc_0_11_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_274_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_0_11_i_qa,
      wea => xt_rsc_0_11_wea,
      da => xt_rsc_0_11_i_da,
      adra => xt_rsc_0_11_i_adra,
      adra_d => xt_rsc_0_11_i_adra_d,
      da_d => xt_rsc_0_11_i_da_d,
      qa_d => xt_rsc_0_11_i_qa_d_1,
      wea_d => xt_rsc_0_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_0_i_wea_d_iff
    );
  xt_rsc_0_11_i_qa <= xt_rsc_0_11_qa;
  xt_rsc_0_11_da <= xt_rsc_0_11_i_da;
  xt_rsc_0_11_adra <= xt_rsc_0_11_i_adra;
  xt_rsc_0_11_i_adra_d <= xt_rsc_0_11_i_adra_d_iff;
  xt_rsc_0_11_i_da_d <= xt_rsc_0_11_i_da_d_iff;
  xt_rsc_0_11_i_qa_d <= xt_rsc_0_11_i_qa_d_1;

  xt_rsc_0_12_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_275_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_0_12_i_qa,
      wea => xt_rsc_0_12_wea,
      da => xt_rsc_0_12_i_da,
      adra => xt_rsc_0_12_i_adra,
      adra_d => xt_rsc_0_12_i_adra_d,
      da_d => xt_rsc_0_12_i_da_d,
      qa_d => xt_rsc_0_12_i_qa_d_1,
      wea_d => xt_rsc_0_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_0_i_wea_d_iff
    );
  xt_rsc_0_12_i_qa <= xt_rsc_0_12_qa;
  xt_rsc_0_12_da <= xt_rsc_0_12_i_da;
  xt_rsc_0_12_adra <= xt_rsc_0_12_i_adra;
  xt_rsc_0_12_i_adra_d <= xt_rsc_0_12_i_adra_d_iff;
  xt_rsc_0_12_i_da_d <= xt_rsc_0_12_i_da_d_iff;
  xt_rsc_0_12_i_qa_d <= xt_rsc_0_12_i_qa_d_1;

  xt_rsc_0_13_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_276_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_0_13_i_qa,
      wea => xt_rsc_0_13_wea,
      da => xt_rsc_0_13_i_da,
      adra => xt_rsc_0_13_i_adra,
      adra_d => xt_rsc_0_13_i_adra_d,
      da_d => xt_rsc_0_13_i_da_d,
      qa_d => xt_rsc_0_13_i_qa_d_1,
      wea_d => xt_rsc_0_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_0_i_wea_d_iff
    );
  xt_rsc_0_13_i_qa <= xt_rsc_0_13_qa;
  xt_rsc_0_13_da <= xt_rsc_0_13_i_da;
  xt_rsc_0_13_adra <= xt_rsc_0_13_i_adra;
  xt_rsc_0_13_i_adra_d <= xt_rsc_0_13_i_adra_d_iff;
  xt_rsc_0_13_i_da_d <= xt_rsc_0_13_i_da_d_iff;
  xt_rsc_0_13_i_qa_d <= xt_rsc_0_13_i_qa_d_1;

  xt_rsc_0_14_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_277_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_0_14_i_qa,
      wea => xt_rsc_0_14_wea,
      da => xt_rsc_0_14_i_da,
      adra => xt_rsc_0_14_i_adra,
      adra_d => xt_rsc_0_14_i_adra_d,
      da_d => xt_rsc_0_14_i_da_d,
      qa_d => xt_rsc_0_14_i_qa_d_1,
      wea_d => xt_rsc_0_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_0_i_wea_d_iff
    );
  xt_rsc_0_14_i_qa <= xt_rsc_0_14_qa;
  xt_rsc_0_14_da <= xt_rsc_0_14_i_da;
  xt_rsc_0_14_adra <= xt_rsc_0_14_i_adra;
  xt_rsc_0_14_i_adra_d <= xt_rsc_0_14_i_adra_d_iff;
  xt_rsc_0_14_i_da_d <= xt_rsc_0_14_i_da_d_iff;
  xt_rsc_0_14_i_qa_d <= xt_rsc_0_14_i_qa_d_1;

  xt_rsc_0_15_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_278_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_0_15_i_qa,
      wea => xt_rsc_0_15_wea,
      da => xt_rsc_0_15_i_da,
      adra => xt_rsc_0_15_i_adra,
      adra_d => xt_rsc_0_15_i_adra_d,
      da_d => xt_rsc_0_15_i_da_d,
      qa_d => xt_rsc_0_15_i_qa_d_1,
      wea_d => xt_rsc_0_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_0_i_wea_d_iff
    );
  xt_rsc_0_15_i_qa <= xt_rsc_0_15_qa;
  xt_rsc_0_15_da <= xt_rsc_0_15_i_da;
  xt_rsc_0_15_adra <= xt_rsc_0_15_i_adra;
  xt_rsc_0_15_i_adra_d <= xt_rsc_0_15_i_adra_d_iff;
  xt_rsc_0_15_i_da_d <= xt_rsc_0_15_i_da_d_iff;
  xt_rsc_0_15_i_qa_d <= xt_rsc_0_15_i_qa_d_1;

  xt_rsc_0_16_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_279_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_0_16_i_qa,
      wea => xt_rsc_0_16_wea,
      da => xt_rsc_0_16_i_da,
      adra => xt_rsc_0_16_i_adra,
      adra_d => xt_rsc_0_16_i_adra_d,
      da_d => xt_rsc_0_16_i_da_d,
      qa_d => xt_rsc_0_16_i_qa_d_1,
      wea_d => xt_rsc_0_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_16_i_wea_d_iff
    );
  xt_rsc_0_16_i_qa <= xt_rsc_0_16_qa;
  xt_rsc_0_16_da <= xt_rsc_0_16_i_da;
  xt_rsc_0_16_adra <= xt_rsc_0_16_i_adra;
  xt_rsc_0_16_i_adra_d <= xt_rsc_0_0_i_adra_d_iff;
  xt_rsc_0_16_i_da_d <= xt_rsc_0_0_i_da_d_iff;
  xt_rsc_0_16_i_qa_d <= xt_rsc_0_16_i_qa_d_1;

  xt_rsc_0_17_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_280_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_0_17_i_qa,
      wea => xt_rsc_0_17_wea,
      da => xt_rsc_0_17_i_da,
      adra => xt_rsc_0_17_i_adra,
      adra_d => xt_rsc_0_17_i_adra_d,
      da_d => xt_rsc_0_17_i_da_d,
      qa_d => xt_rsc_0_17_i_qa_d_1,
      wea_d => xt_rsc_0_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_16_i_wea_d_iff
    );
  xt_rsc_0_17_i_qa <= xt_rsc_0_17_qa;
  xt_rsc_0_17_da <= xt_rsc_0_17_i_da;
  xt_rsc_0_17_adra <= xt_rsc_0_17_i_adra;
  xt_rsc_0_17_i_adra_d <= xt_rsc_0_1_i_adra_d_iff;
  xt_rsc_0_17_i_da_d <= xt_rsc_0_1_i_da_d_iff;
  xt_rsc_0_17_i_qa_d <= xt_rsc_0_17_i_qa_d_1;

  xt_rsc_0_18_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_281_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_0_18_i_qa,
      wea => xt_rsc_0_18_wea,
      da => xt_rsc_0_18_i_da,
      adra => xt_rsc_0_18_i_adra,
      adra_d => xt_rsc_0_18_i_adra_d,
      da_d => xt_rsc_0_18_i_da_d,
      qa_d => xt_rsc_0_18_i_qa_d_1,
      wea_d => xt_rsc_0_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_16_i_wea_d_iff
    );
  xt_rsc_0_18_i_qa <= xt_rsc_0_18_qa;
  xt_rsc_0_18_da <= xt_rsc_0_18_i_da;
  xt_rsc_0_18_adra <= xt_rsc_0_18_i_adra;
  xt_rsc_0_18_i_adra_d <= xt_rsc_0_2_i_adra_d_iff;
  xt_rsc_0_18_i_da_d <= xt_rsc_0_2_i_da_d_iff;
  xt_rsc_0_18_i_qa_d <= xt_rsc_0_18_i_qa_d_1;

  xt_rsc_0_19_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_282_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_0_19_i_qa,
      wea => xt_rsc_0_19_wea,
      da => xt_rsc_0_19_i_da,
      adra => xt_rsc_0_19_i_adra,
      adra_d => xt_rsc_0_19_i_adra_d,
      da_d => xt_rsc_0_19_i_da_d,
      qa_d => xt_rsc_0_19_i_qa_d_1,
      wea_d => xt_rsc_0_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_16_i_wea_d_iff
    );
  xt_rsc_0_19_i_qa <= xt_rsc_0_19_qa;
  xt_rsc_0_19_da <= xt_rsc_0_19_i_da;
  xt_rsc_0_19_adra <= xt_rsc_0_19_i_adra;
  xt_rsc_0_19_i_adra_d <= xt_rsc_0_3_i_adra_d_iff;
  xt_rsc_0_19_i_da_d <= xt_rsc_0_3_i_da_d_iff;
  xt_rsc_0_19_i_qa_d <= xt_rsc_0_19_i_qa_d_1;

  xt_rsc_0_20_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_283_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_0_20_i_qa,
      wea => xt_rsc_0_20_wea,
      da => xt_rsc_0_20_i_da,
      adra => xt_rsc_0_20_i_adra,
      adra_d => xt_rsc_0_20_i_adra_d,
      da_d => xt_rsc_0_20_i_da_d,
      qa_d => xt_rsc_0_20_i_qa_d_1,
      wea_d => xt_rsc_0_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_16_i_wea_d_iff
    );
  xt_rsc_0_20_i_qa <= xt_rsc_0_20_qa;
  xt_rsc_0_20_da <= xt_rsc_0_20_i_da;
  xt_rsc_0_20_adra <= xt_rsc_0_20_i_adra;
  xt_rsc_0_20_i_adra_d <= xt_rsc_0_4_i_adra_d_iff;
  xt_rsc_0_20_i_da_d <= xt_rsc_0_4_i_da_d_iff;
  xt_rsc_0_20_i_qa_d <= xt_rsc_0_20_i_qa_d_1;

  xt_rsc_0_21_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_284_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_0_21_i_qa,
      wea => xt_rsc_0_21_wea,
      da => xt_rsc_0_21_i_da,
      adra => xt_rsc_0_21_i_adra,
      adra_d => xt_rsc_0_21_i_adra_d,
      da_d => xt_rsc_0_21_i_da_d,
      qa_d => xt_rsc_0_21_i_qa_d_1,
      wea_d => xt_rsc_0_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_16_i_wea_d_iff
    );
  xt_rsc_0_21_i_qa <= xt_rsc_0_21_qa;
  xt_rsc_0_21_da <= xt_rsc_0_21_i_da;
  xt_rsc_0_21_adra <= xt_rsc_0_21_i_adra;
  xt_rsc_0_21_i_adra_d <= xt_rsc_0_5_i_adra_d_iff;
  xt_rsc_0_21_i_da_d <= xt_rsc_0_5_i_da_d_iff;
  xt_rsc_0_21_i_qa_d <= xt_rsc_0_21_i_qa_d_1;

  xt_rsc_0_22_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_285_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_0_22_i_qa,
      wea => xt_rsc_0_22_wea,
      da => xt_rsc_0_22_i_da,
      adra => xt_rsc_0_22_i_adra,
      adra_d => xt_rsc_0_22_i_adra_d,
      da_d => xt_rsc_0_22_i_da_d,
      qa_d => xt_rsc_0_22_i_qa_d_1,
      wea_d => xt_rsc_0_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_16_i_wea_d_iff
    );
  xt_rsc_0_22_i_qa <= xt_rsc_0_22_qa;
  xt_rsc_0_22_da <= xt_rsc_0_22_i_da;
  xt_rsc_0_22_adra <= xt_rsc_0_22_i_adra;
  xt_rsc_0_22_i_adra_d <= xt_rsc_0_6_i_adra_d_iff;
  xt_rsc_0_22_i_da_d <= xt_rsc_0_6_i_da_d_iff;
  xt_rsc_0_22_i_qa_d <= xt_rsc_0_22_i_qa_d_1;

  xt_rsc_0_23_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_286_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_0_23_i_qa,
      wea => xt_rsc_0_23_wea,
      da => xt_rsc_0_23_i_da,
      adra => xt_rsc_0_23_i_adra,
      adra_d => xt_rsc_0_23_i_adra_d,
      da_d => xt_rsc_0_23_i_da_d,
      qa_d => xt_rsc_0_23_i_qa_d_1,
      wea_d => xt_rsc_0_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_16_i_wea_d_iff
    );
  xt_rsc_0_23_i_qa <= xt_rsc_0_23_qa;
  xt_rsc_0_23_da <= xt_rsc_0_23_i_da;
  xt_rsc_0_23_adra <= xt_rsc_0_23_i_adra;
  xt_rsc_0_23_i_adra_d <= xt_rsc_0_7_i_adra_d_iff;
  xt_rsc_0_23_i_da_d <= xt_rsc_0_7_i_da_d_iff;
  xt_rsc_0_23_i_qa_d <= xt_rsc_0_23_i_qa_d_1;

  xt_rsc_0_24_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_287_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_0_24_i_qa,
      wea => xt_rsc_0_24_wea,
      da => xt_rsc_0_24_i_da,
      adra => xt_rsc_0_24_i_adra,
      adra_d => xt_rsc_0_24_i_adra_d,
      da_d => xt_rsc_0_24_i_da_d,
      qa_d => xt_rsc_0_24_i_qa_d_1,
      wea_d => xt_rsc_0_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_16_i_wea_d_iff
    );
  xt_rsc_0_24_i_qa <= xt_rsc_0_24_qa;
  xt_rsc_0_24_da <= xt_rsc_0_24_i_da;
  xt_rsc_0_24_adra <= xt_rsc_0_24_i_adra;
  xt_rsc_0_24_i_adra_d <= xt_rsc_0_8_i_adra_d_iff;
  xt_rsc_0_24_i_da_d <= xt_rsc_0_8_i_da_d_iff;
  xt_rsc_0_24_i_qa_d <= xt_rsc_0_24_i_qa_d_1;

  xt_rsc_0_25_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_288_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_0_25_i_qa,
      wea => xt_rsc_0_25_wea,
      da => xt_rsc_0_25_i_da,
      adra => xt_rsc_0_25_i_adra,
      adra_d => xt_rsc_0_25_i_adra_d,
      da_d => xt_rsc_0_25_i_da_d,
      qa_d => xt_rsc_0_25_i_qa_d_1,
      wea_d => xt_rsc_0_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_16_i_wea_d_iff
    );
  xt_rsc_0_25_i_qa <= xt_rsc_0_25_qa;
  xt_rsc_0_25_da <= xt_rsc_0_25_i_da;
  xt_rsc_0_25_adra <= xt_rsc_0_25_i_adra;
  xt_rsc_0_25_i_adra_d <= xt_rsc_0_9_i_adra_d_iff;
  xt_rsc_0_25_i_da_d <= xt_rsc_0_9_i_da_d_iff;
  xt_rsc_0_25_i_qa_d <= xt_rsc_0_25_i_qa_d_1;

  xt_rsc_0_26_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_289_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_0_26_i_qa,
      wea => xt_rsc_0_26_wea,
      da => xt_rsc_0_26_i_da,
      adra => xt_rsc_0_26_i_adra,
      adra_d => xt_rsc_0_26_i_adra_d,
      da_d => xt_rsc_0_26_i_da_d,
      qa_d => xt_rsc_0_26_i_qa_d_1,
      wea_d => xt_rsc_0_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_16_i_wea_d_iff
    );
  xt_rsc_0_26_i_qa <= xt_rsc_0_26_qa;
  xt_rsc_0_26_da <= xt_rsc_0_26_i_da;
  xt_rsc_0_26_adra <= xt_rsc_0_26_i_adra;
  xt_rsc_0_26_i_adra_d <= xt_rsc_0_10_i_adra_d_iff;
  xt_rsc_0_26_i_da_d <= xt_rsc_0_10_i_da_d_iff;
  xt_rsc_0_26_i_qa_d <= xt_rsc_0_26_i_qa_d_1;

  xt_rsc_0_27_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_290_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_0_27_i_qa,
      wea => xt_rsc_0_27_wea,
      da => xt_rsc_0_27_i_da,
      adra => xt_rsc_0_27_i_adra,
      adra_d => xt_rsc_0_27_i_adra_d,
      da_d => xt_rsc_0_27_i_da_d,
      qa_d => xt_rsc_0_27_i_qa_d_1,
      wea_d => xt_rsc_0_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_16_i_wea_d_iff
    );
  xt_rsc_0_27_i_qa <= xt_rsc_0_27_qa;
  xt_rsc_0_27_da <= xt_rsc_0_27_i_da;
  xt_rsc_0_27_adra <= xt_rsc_0_27_i_adra;
  xt_rsc_0_27_i_adra_d <= xt_rsc_0_11_i_adra_d_iff;
  xt_rsc_0_27_i_da_d <= xt_rsc_0_11_i_da_d_iff;
  xt_rsc_0_27_i_qa_d <= xt_rsc_0_27_i_qa_d_1;

  xt_rsc_0_28_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_291_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_0_28_i_qa,
      wea => xt_rsc_0_28_wea,
      da => xt_rsc_0_28_i_da,
      adra => xt_rsc_0_28_i_adra,
      adra_d => xt_rsc_0_28_i_adra_d,
      da_d => xt_rsc_0_28_i_da_d,
      qa_d => xt_rsc_0_28_i_qa_d_1,
      wea_d => xt_rsc_0_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_16_i_wea_d_iff
    );
  xt_rsc_0_28_i_qa <= xt_rsc_0_28_qa;
  xt_rsc_0_28_da <= xt_rsc_0_28_i_da;
  xt_rsc_0_28_adra <= xt_rsc_0_28_i_adra;
  xt_rsc_0_28_i_adra_d <= xt_rsc_0_12_i_adra_d_iff;
  xt_rsc_0_28_i_da_d <= xt_rsc_0_12_i_da_d_iff;
  xt_rsc_0_28_i_qa_d <= xt_rsc_0_28_i_qa_d_1;

  xt_rsc_0_29_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_292_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_0_29_i_qa,
      wea => xt_rsc_0_29_wea,
      da => xt_rsc_0_29_i_da,
      adra => xt_rsc_0_29_i_adra,
      adra_d => xt_rsc_0_29_i_adra_d,
      da_d => xt_rsc_0_29_i_da_d,
      qa_d => xt_rsc_0_29_i_qa_d_1,
      wea_d => xt_rsc_0_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_16_i_wea_d_iff
    );
  xt_rsc_0_29_i_qa <= xt_rsc_0_29_qa;
  xt_rsc_0_29_da <= xt_rsc_0_29_i_da;
  xt_rsc_0_29_adra <= xt_rsc_0_29_i_adra;
  xt_rsc_0_29_i_adra_d <= xt_rsc_0_13_i_adra_d_iff;
  xt_rsc_0_29_i_da_d <= xt_rsc_0_13_i_da_d_iff;
  xt_rsc_0_29_i_qa_d <= xt_rsc_0_29_i_qa_d_1;

  xt_rsc_0_30_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_293_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_0_30_i_qa,
      wea => xt_rsc_0_30_wea,
      da => xt_rsc_0_30_i_da,
      adra => xt_rsc_0_30_i_adra,
      adra_d => xt_rsc_0_30_i_adra_d,
      da_d => xt_rsc_0_30_i_da_d,
      qa_d => xt_rsc_0_30_i_qa_d_1,
      wea_d => xt_rsc_0_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_16_i_wea_d_iff
    );
  xt_rsc_0_30_i_qa <= xt_rsc_0_30_qa;
  xt_rsc_0_30_da <= xt_rsc_0_30_i_da;
  xt_rsc_0_30_adra <= xt_rsc_0_30_i_adra;
  xt_rsc_0_30_i_adra_d <= xt_rsc_0_14_i_adra_d_iff;
  xt_rsc_0_30_i_da_d <= xt_rsc_0_14_i_da_d_iff;
  xt_rsc_0_30_i_qa_d <= xt_rsc_0_30_i_qa_d_1;

  xt_rsc_0_31_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_294_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_0_31_i_qa,
      wea => xt_rsc_0_31_wea,
      da => xt_rsc_0_31_i_da,
      adra => xt_rsc_0_31_i_adra,
      adra_d => xt_rsc_0_31_i_adra_d,
      da_d => xt_rsc_0_31_i_da_d,
      qa_d => xt_rsc_0_31_i_qa_d_1,
      wea_d => xt_rsc_0_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_16_i_wea_d_iff
    );
  xt_rsc_0_31_i_qa <= xt_rsc_0_31_qa;
  xt_rsc_0_31_da <= xt_rsc_0_31_i_da;
  xt_rsc_0_31_adra <= xt_rsc_0_31_i_adra;
  xt_rsc_0_31_i_adra_d <= xt_rsc_0_15_i_adra_d_iff;
  xt_rsc_0_31_i_da_d <= xt_rsc_0_15_i_da_d_iff;
  xt_rsc_0_31_i_qa_d <= xt_rsc_0_31_i_qa_d_1;

  xt_rsc_1_0_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_295_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_1_0_i_qa,
      wea => xt_rsc_1_0_wea,
      da => xt_rsc_1_0_i_da,
      adra => xt_rsc_1_0_i_adra,
      adra_d => xt_rsc_1_0_i_adra_d,
      da_d => xt_rsc_1_0_i_da_d,
      qa_d => xt_rsc_1_0_i_qa_d_1,
      wea_d => xt_rsc_1_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_0_i_wea_d_iff
    );
  xt_rsc_1_0_i_qa <= xt_rsc_1_0_qa;
  xt_rsc_1_0_da <= xt_rsc_1_0_i_da;
  xt_rsc_1_0_adra <= xt_rsc_1_0_i_adra;
  xt_rsc_1_0_i_adra_d <= xt_rsc_0_0_i_adra_d_iff;
  xt_rsc_1_0_i_da_d <= xt_rsc_0_0_i_da_d_iff;
  xt_rsc_1_0_i_qa_d <= xt_rsc_1_0_i_qa_d_1;

  xt_rsc_1_1_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_296_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_1_1_i_qa,
      wea => xt_rsc_1_1_wea,
      da => xt_rsc_1_1_i_da,
      adra => xt_rsc_1_1_i_adra,
      adra_d => xt_rsc_1_1_i_adra_d,
      da_d => xt_rsc_1_1_i_da_d,
      qa_d => xt_rsc_1_1_i_qa_d_1,
      wea_d => xt_rsc_1_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_0_i_wea_d_iff
    );
  xt_rsc_1_1_i_qa <= xt_rsc_1_1_qa;
  xt_rsc_1_1_da <= xt_rsc_1_1_i_da;
  xt_rsc_1_1_adra <= xt_rsc_1_1_i_adra;
  xt_rsc_1_1_i_adra_d <= xt_rsc_0_1_i_adra_d_iff;
  xt_rsc_1_1_i_da_d <= xt_rsc_0_1_i_da_d_iff;
  xt_rsc_1_1_i_qa_d <= xt_rsc_1_1_i_qa_d_1;

  xt_rsc_1_2_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_297_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_1_2_i_qa,
      wea => xt_rsc_1_2_wea,
      da => xt_rsc_1_2_i_da,
      adra => xt_rsc_1_2_i_adra,
      adra_d => xt_rsc_1_2_i_adra_d,
      da_d => xt_rsc_1_2_i_da_d,
      qa_d => xt_rsc_1_2_i_qa_d_1,
      wea_d => xt_rsc_1_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_0_i_wea_d_iff
    );
  xt_rsc_1_2_i_qa <= xt_rsc_1_2_qa;
  xt_rsc_1_2_da <= xt_rsc_1_2_i_da;
  xt_rsc_1_2_adra <= xt_rsc_1_2_i_adra;
  xt_rsc_1_2_i_adra_d <= xt_rsc_0_2_i_adra_d_iff;
  xt_rsc_1_2_i_da_d <= xt_rsc_0_2_i_da_d_iff;
  xt_rsc_1_2_i_qa_d <= xt_rsc_1_2_i_qa_d_1;

  xt_rsc_1_3_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_298_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_1_3_i_qa,
      wea => xt_rsc_1_3_wea,
      da => xt_rsc_1_3_i_da,
      adra => xt_rsc_1_3_i_adra,
      adra_d => xt_rsc_1_3_i_adra_d,
      da_d => xt_rsc_1_3_i_da_d,
      qa_d => xt_rsc_1_3_i_qa_d_1,
      wea_d => xt_rsc_1_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_0_i_wea_d_iff
    );
  xt_rsc_1_3_i_qa <= xt_rsc_1_3_qa;
  xt_rsc_1_3_da <= xt_rsc_1_3_i_da;
  xt_rsc_1_3_adra <= xt_rsc_1_3_i_adra;
  xt_rsc_1_3_i_adra_d <= xt_rsc_0_3_i_adra_d_iff;
  xt_rsc_1_3_i_da_d <= xt_rsc_0_3_i_da_d_iff;
  xt_rsc_1_3_i_qa_d <= xt_rsc_1_3_i_qa_d_1;

  xt_rsc_1_4_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_299_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_1_4_i_qa,
      wea => xt_rsc_1_4_wea,
      da => xt_rsc_1_4_i_da,
      adra => xt_rsc_1_4_i_adra,
      adra_d => xt_rsc_1_4_i_adra_d,
      da_d => xt_rsc_1_4_i_da_d,
      qa_d => xt_rsc_1_4_i_qa_d_1,
      wea_d => xt_rsc_1_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_0_i_wea_d_iff
    );
  xt_rsc_1_4_i_qa <= xt_rsc_1_4_qa;
  xt_rsc_1_4_da <= xt_rsc_1_4_i_da;
  xt_rsc_1_4_adra <= xt_rsc_1_4_i_adra;
  xt_rsc_1_4_i_adra_d <= xt_rsc_0_4_i_adra_d_iff;
  xt_rsc_1_4_i_da_d <= xt_rsc_0_4_i_da_d_iff;
  xt_rsc_1_4_i_qa_d <= xt_rsc_1_4_i_qa_d_1;

  xt_rsc_1_5_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_300_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_1_5_i_qa,
      wea => xt_rsc_1_5_wea,
      da => xt_rsc_1_5_i_da,
      adra => xt_rsc_1_5_i_adra,
      adra_d => xt_rsc_1_5_i_adra_d,
      da_d => xt_rsc_1_5_i_da_d,
      qa_d => xt_rsc_1_5_i_qa_d_1,
      wea_d => xt_rsc_1_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_0_i_wea_d_iff
    );
  xt_rsc_1_5_i_qa <= xt_rsc_1_5_qa;
  xt_rsc_1_5_da <= xt_rsc_1_5_i_da;
  xt_rsc_1_5_adra <= xt_rsc_1_5_i_adra;
  xt_rsc_1_5_i_adra_d <= xt_rsc_0_5_i_adra_d_iff;
  xt_rsc_1_5_i_da_d <= xt_rsc_0_5_i_da_d_iff;
  xt_rsc_1_5_i_qa_d <= xt_rsc_1_5_i_qa_d_1;

  xt_rsc_1_6_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_301_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_1_6_i_qa,
      wea => xt_rsc_1_6_wea,
      da => xt_rsc_1_6_i_da,
      adra => xt_rsc_1_6_i_adra,
      adra_d => xt_rsc_1_6_i_adra_d,
      da_d => xt_rsc_1_6_i_da_d,
      qa_d => xt_rsc_1_6_i_qa_d_1,
      wea_d => xt_rsc_1_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_0_i_wea_d_iff
    );
  xt_rsc_1_6_i_qa <= xt_rsc_1_6_qa;
  xt_rsc_1_6_da <= xt_rsc_1_6_i_da;
  xt_rsc_1_6_adra <= xt_rsc_1_6_i_adra;
  xt_rsc_1_6_i_adra_d <= xt_rsc_0_6_i_adra_d_iff;
  xt_rsc_1_6_i_da_d <= xt_rsc_0_6_i_da_d_iff;
  xt_rsc_1_6_i_qa_d <= xt_rsc_1_6_i_qa_d_1;

  xt_rsc_1_7_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_302_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_1_7_i_qa,
      wea => xt_rsc_1_7_wea,
      da => xt_rsc_1_7_i_da,
      adra => xt_rsc_1_7_i_adra,
      adra_d => xt_rsc_1_7_i_adra_d,
      da_d => xt_rsc_1_7_i_da_d,
      qa_d => xt_rsc_1_7_i_qa_d_1,
      wea_d => xt_rsc_1_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_0_i_wea_d_iff
    );
  xt_rsc_1_7_i_qa <= xt_rsc_1_7_qa;
  xt_rsc_1_7_da <= xt_rsc_1_7_i_da;
  xt_rsc_1_7_adra <= xt_rsc_1_7_i_adra;
  xt_rsc_1_7_i_adra_d <= xt_rsc_0_7_i_adra_d_iff;
  xt_rsc_1_7_i_da_d <= xt_rsc_0_7_i_da_d_iff;
  xt_rsc_1_7_i_qa_d <= xt_rsc_1_7_i_qa_d_1;

  xt_rsc_1_8_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_303_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_1_8_i_qa,
      wea => xt_rsc_1_8_wea,
      da => xt_rsc_1_8_i_da,
      adra => xt_rsc_1_8_i_adra,
      adra_d => xt_rsc_1_8_i_adra_d,
      da_d => xt_rsc_1_8_i_da_d,
      qa_d => xt_rsc_1_8_i_qa_d_1,
      wea_d => xt_rsc_1_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_0_i_wea_d_iff
    );
  xt_rsc_1_8_i_qa <= xt_rsc_1_8_qa;
  xt_rsc_1_8_da <= xt_rsc_1_8_i_da;
  xt_rsc_1_8_adra <= xt_rsc_1_8_i_adra;
  xt_rsc_1_8_i_adra_d <= xt_rsc_0_8_i_adra_d_iff;
  xt_rsc_1_8_i_da_d <= xt_rsc_0_8_i_da_d_iff;
  xt_rsc_1_8_i_qa_d <= xt_rsc_1_8_i_qa_d_1;

  xt_rsc_1_9_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_304_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_1_9_i_qa,
      wea => xt_rsc_1_9_wea,
      da => xt_rsc_1_9_i_da,
      adra => xt_rsc_1_9_i_adra,
      adra_d => xt_rsc_1_9_i_adra_d,
      da_d => xt_rsc_1_9_i_da_d,
      qa_d => xt_rsc_1_9_i_qa_d_1,
      wea_d => xt_rsc_1_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_0_i_wea_d_iff
    );
  xt_rsc_1_9_i_qa <= xt_rsc_1_9_qa;
  xt_rsc_1_9_da <= xt_rsc_1_9_i_da;
  xt_rsc_1_9_adra <= xt_rsc_1_9_i_adra;
  xt_rsc_1_9_i_adra_d <= xt_rsc_0_9_i_adra_d_iff;
  xt_rsc_1_9_i_da_d <= xt_rsc_0_9_i_da_d_iff;
  xt_rsc_1_9_i_qa_d <= xt_rsc_1_9_i_qa_d_1;

  xt_rsc_1_10_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_305_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_1_10_i_qa,
      wea => xt_rsc_1_10_wea,
      da => xt_rsc_1_10_i_da,
      adra => xt_rsc_1_10_i_adra,
      adra_d => xt_rsc_1_10_i_adra_d,
      da_d => xt_rsc_1_10_i_da_d,
      qa_d => xt_rsc_1_10_i_qa_d_1,
      wea_d => xt_rsc_1_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_0_i_wea_d_iff
    );
  xt_rsc_1_10_i_qa <= xt_rsc_1_10_qa;
  xt_rsc_1_10_da <= xt_rsc_1_10_i_da;
  xt_rsc_1_10_adra <= xt_rsc_1_10_i_adra;
  xt_rsc_1_10_i_adra_d <= xt_rsc_0_10_i_adra_d_iff;
  xt_rsc_1_10_i_da_d <= xt_rsc_0_10_i_da_d_iff;
  xt_rsc_1_10_i_qa_d <= xt_rsc_1_10_i_qa_d_1;

  xt_rsc_1_11_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_306_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_1_11_i_qa,
      wea => xt_rsc_1_11_wea,
      da => xt_rsc_1_11_i_da,
      adra => xt_rsc_1_11_i_adra,
      adra_d => xt_rsc_1_11_i_adra_d,
      da_d => xt_rsc_1_11_i_da_d,
      qa_d => xt_rsc_1_11_i_qa_d_1,
      wea_d => xt_rsc_1_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_0_i_wea_d_iff
    );
  xt_rsc_1_11_i_qa <= xt_rsc_1_11_qa;
  xt_rsc_1_11_da <= xt_rsc_1_11_i_da;
  xt_rsc_1_11_adra <= xt_rsc_1_11_i_adra;
  xt_rsc_1_11_i_adra_d <= xt_rsc_0_11_i_adra_d_iff;
  xt_rsc_1_11_i_da_d <= xt_rsc_0_11_i_da_d_iff;
  xt_rsc_1_11_i_qa_d <= xt_rsc_1_11_i_qa_d_1;

  xt_rsc_1_12_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_307_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_1_12_i_qa,
      wea => xt_rsc_1_12_wea,
      da => xt_rsc_1_12_i_da,
      adra => xt_rsc_1_12_i_adra,
      adra_d => xt_rsc_1_12_i_adra_d,
      da_d => xt_rsc_1_12_i_da_d,
      qa_d => xt_rsc_1_12_i_qa_d_1,
      wea_d => xt_rsc_1_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_0_i_wea_d_iff
    );
  xt_rsc_1_12_i_qa <= xt_rsc_1_12_qa;
  xt_rsc_1_12_da <= xt_rsc_1_12_i_da;
  xt_rsc_1_12_adra <= xt_rsc_1_12_i_adra;
  xt_rsc_1_12_i_adra_d <= xt_rsc_0_12_i_adra_d_iff;
  xt_rsc_1_12_i_da_d <= xt_rsc_0_12_i_da_d_iff;
  xt_rsc_1_12_i_qa_d <= xt_rsc_1_12_i_qa_d_1;

  xt_rsc_1_13_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_308_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_1_13_i_qa,
      wea => xt_rsc_1_13_wea,
      da => xt_rsc_1_13_i_da,
      adra => xt_rsc_1_13_i_adra,
      adra_d => xt_rsc_1_13_i_adra_d,
      da_d => xt_rsc_1_13_i_da_d,
      qa_d => xt_rsc_1_13_i_qa_d_1,
      wea_d => xt_rsc_1_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_0_i_wea_d_iff
    );
  xt_rsc_1_13_i_qa <= xt_rsc_1_13_qa;
  xt_rsc_1_13_da <= xt_rsc_1_13_i_da;
  xt_rsc_1_13_adra <= xt_rsc_1_13_i_adra;
  xt_rsc_1_13_i_adra_d <= xt_rsc_0_13_i_adra_d_iff;
  xt_rsc_1_13_i_da_d <= xt_rsc_0_13_i_da_d_iff;
  xt_rsc_1_13_i_qa_d <= xt_rsc_1_13_i_qa_d_1;

  xt_rsc_1_14_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_309_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_1_14_i_qa,
      wea => xt_rsc_1_14_wea,
      da => xt_rsc_1_14_i_da,
      adra => xt_rsc_1_14_i_adra,
      adra_d => xt_rsc_1_14_i_adra_d,
      da_d => xt_rsc_1_14_i_da_d,
      qa_d => xt_rsc_1_14_i_qa_d_1,
      wea_d => xt_rsc_1_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_0_i_wea_d_iff
    );
  xt_rsc_1_14_i_qa <= xt_rsc_1_14_qa;
  xt_rsc_1_14_da <= xt_rsc_1_14_i_da;
  xt_rsc_1_14_adra <= xt_rsc_1_14_i_adra;
  xt_rsc_1_14_i_adra_d <= xt_rsc_0_14_i_adra_d_iff;
  xt_rsc_1_14_i_da_d <= xt_rsc_0_14_i_da_d_iff;
  xt_rsc_1_14_i_qa_d <= xt_rsc_1_14_i_qa_d_1;

  xt_rsc_1_15_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_310_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_1_15_i_qa,
      wea => xt_rsc_1_15_wea,
      da => xt_rsc_1_15_i_da,
      adra => xt_rsc_1_15_i_adra,
      adra_d => xt_rsc_1_15_i_adra_d,
      da_d => xt_rsc_1_15_i_da_d,
      qa_d => xt_rsc_1_15_i_qa_d_1,
      wea_d => xt_rsc_1_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_0_i_wea_d_iff
    );
  xt_rsc_1_15_i_qa <= xt_rsc_1_15_qa;
  xt_rsc_1_15_da <= xt_rsc_1_15_i_da;
  xt_rsc_1_15_adra <= xt_rsc_1_15_i_adra;
  xt_rsc_1_15_i_adra_d <= xt_rsc_0_15_i_adra_d_iff;
  xt_rsc_1_15_i_da_d <= xt_rsc_0_15_i_da_d_iff;
  xt_rsc_1_15_i_qa_d <= xt_rsc_1_15_i_qa_d_1;

  xt_rsc_1_16_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_311_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_1_16_i_qa,
      wea => xt_rsc_1_16_wea,
      da => xt_rsc_1_16_i_da,
      adra => xt_rsc_1_16_i_adra,
      adra_d => xt_rsc_1_16_i_adra_d,
      da_d => xt_rsc_1_16_i_da_d,
      qa_d => xt_rsc_1_16_i_qa_d_1,
      wea_d => xt_rsc_1_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_16_i_wea_d_iff
    );
  xt_rsc_1_16_i_qa <= xt_rsc_1_16_qa;
  xt_rsc_1_16_da <= xt_rsc_1_16_i_da;
  xt_rsc_1_16_adra <= xt_rsc_1_16_i_adra;
  xt_rsc_1_16_i_adra_d <= xt_rsc_0_0_i_adra_d_iff;
  xt_rsc_1_16_i_da_d <= xt_rsc_0_0_i_da_d_iff;
  xt_rsc_1_16_i_qa_d <= xt_rsc_1_16_i_qa_d_1;

  xt_rsc_1_17_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_312_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_1_17_i_qa,
      wea => xt_rsc_1_17_wea,
      da => xt_rsc_1_17_i_da,
      adra => xt_rsc_1_17_i_adra,
      adra_d => xt_rsc_1_17_i_adra_d,
      da_d => xt_rsc_1_17_i_da_d,
      qa_d => xt_rsc_1_17_i_qa_d_1,
      wea_d => xt_rsc_1_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_16_i_wea_d_iff
    );
  xt_rsc_1_17_i_qa <= xt_rsc_1_17_qa;
  xt_rsc_1_17_da <= xt_rsc_1_17_i_da;
  xt_rsc_1_17_adra <= xt_rsc_1_17_i_adra;
  xt_rsc_1_17_i_adra_d <= xt_rsc_0_1_i_adra_d_iff;
  xt_rsc_1_17_i_da_d <= xt_rsc_0_1_i_da_d_iff;
  xt_rsc_1_17_i_qa_d <= xt_rsc_1_17_i_qa_d_1;

  xt_rsc_1_18_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_313_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_1_18_i_qa,
      wea => xt_rsc_1_18_wea,
      da => xt_rsc_1_18_i_da,
      adra => xt_rsc_1_18_i_adra,
      adra_d => xt_rsc_1_18_i_adra_d,
      da_d => xt_rsc_1_18_i_da_d,
      qa_d => xt_rsc_1_18_i_qa_d_1,
      wea_d => xt_rsc_1_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_16_i_wea_d_iff
    );
  xt_rsc_1_18_i_qa <= xt_rsc_1_18_qa;
  xt_rsc_1_18_da <= xt_rsc_1_18_i_da;
  xt_rsc_1_18_adra <= xt_rsc_1_18_i_adra;
  xt_rsc_1_18_i_adra_d <= xt_rsc_0_2_i_adra_d_iff;
  xt_rsc_1_18_i_da_d <= xt_rsc_0_2_i_da_d_iff;
  xt_rsc_1_18_i_qa_d <= xt_rsc_1_18_i_qa_d_1;

  xt_rsc_1_19_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_314_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_1_19_i_qa,
      wea => xt_rsc_1_19_wea,
      da => xt_rsc_1_19_i_da,
      adra => xt_rsc_1_19_i_adra,
      adra_d => xt_rsc_1_19_i_adra_d,
      da_d => xt_rsc_1_19_i_da_d,
      qa_d => xt_rsc_1_19_i_qa_d_1,
      wea_d => xt_rsc_1_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_16_i_wea_d_iff
    );
  xt_rsc_1_19_i_qa <= xt_rsc_1_19_qa;
  xt_rsc_1_19_da <= xt_rsc_1_19_i_da;
  xt_rsc_1_19_adra <= xt_rsc_1_19_i_adra;
  xt_rsc_1_19_i_adra_d <= xt_rsc_0_3_i_adra_d_iff;
  xt_rsc_1_19_i_da_d <= xt_rsc_0_3_i_da_d_iff;
  xt_rsc_1_19_i_qa_d <= xt_rsc_1_19_i_qa_d_1;

  xt_rsc_1_20_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_315_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_1_20_i_qa,
      wea => xt_rsc_1_20_wea,
      da => xt_rsc_1_20_i_da,
      adra => xt_rsc_1_20_i_adra,
      adra_d => xt_rsc_1_20_i_adra_d,
      da_d => xt_rsc_1_20_i_da_d,
      qa_d => xt_rsc_1_20_i_qa_d_1,
      wea_d => xt_rsc_1_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_16_i_wea_d_iff
    );
  xt_rsc_1_20_i_qa <= xt_rsc_1_20_qa;
  xt_rsc_1_20_da <= xt_rsc_1_20_i_da;
  xt_rsc_1_20_adra <= xt_rsc_1_20_i_adra;
  xt_rsc_1_20_i_adra_d <= xt_rsc_0_4_i_adra_d_iff;
  xt_rsc_1_20_i_da_d <= xt_rsc_0_4_i_da_d_iff;
  xt_rsc_1_20_i_qa_d <= xt_rsc_1_20_i_qa_d_1;

  xt_rsc_1_21_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_316_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_1_21_i_qa,
      wea => xt_rsc_1_21_wea,
      da => xt_rsc_1_21_i_da,
      adra => xt_rsc_1_21_i_adra,
      adra_d => xt_rsc_1_21_i_adra_d,
      da_d => xt_rsc_1_21_i_da_d,
      qa_d => xt_rsc_1_21_i_qa_d_1,
      wea_d => xt_rsc_1_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_16_i_wea_d_iff
    );
  xt_rsc_1_21_i_qa <= xt_rsc_1_21_qa;
  xt_rsc_1_21_da <= xt_rsc_1_21_i_da;
  xt_rsc_1_21_adra <= xt_rsc_1_21_i_adra;
  xt_rsc_1_21_i_adra_d <= xt_rsc_0_5_i_adra_d_iff;
  xt_rsc_1_21_i_da_d <= xt_rsc_0_5_i_da_d_iff;
  xt_rsc_1_21_i_qa_d <= xt_rsc_1_21_i_qa_d_1;

  xt_rsc_1_22_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_317_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_1_22_i_qa,
      wea => xt_rsc_1_22_wea,
      da => xt_rsc_1_22_i_da,
      adra => xt_rsc_1_22_i_adra,
      adra_d => xt_rsc_1_22_i_adra_d,
      da_d => xt_rsc_1_22_i_da_d,
      qa_d => xt_rsc_1_22_i_qa_d_1,
      wea_d => xt_rsc_1_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_16_i_wea_d_iff
    );
  xt_rsc_1_22_i_qa <= xt_rsc_1_22_qa;
  xt_rsc_1_22_da <= xt_rsc_1_22_i_da;
  xt_rsc_1_22_adra <= xt_rsc_1_22_i_adra;
  xt_rsc_1_22_i_adra_d <= xt_rsc_0_6_i_adra_d_iff;
  xt_rsc_1_22_i_da_d <= xt_rsc_0_6_i_da_d_iff;
  xt_rsc_1_22_i_qa_d <= xt_rsc_1_22_i_qa_d_1;

  xt_rsc_1_23_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_318_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_1_23_i_qa,
      wea => xt_rsc_1_23_wea,
      da => xt_rsc_1_23_i_da,
      adra => xt_rsc_1_23_i_adra,
      adra_d => xt_rsc_1_23_i_adra_d,
      da_d => xt_rsc_1_23_i_da_d,
      qa_d => xt_rsc_1_23_i_qa_d_1,
      wea_d => xt_rsc_1_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_16_i_wea_d_iff
    );
  xt_rsc_1_23_i_qa <= xt_rsc_1_23_qa;
  xt_rsc_1_23_da <= xt_rsc_1_23_i_da;
  xt_rsc_1_23_adra <= xt_rsc_1_23_i_adra;
  xt_rsc_1_23_i_adra_d <= xt_rsc_0_7_i_adra_d_iff;
  xt_rsc_1_23_i_da_d <= xt_rsc_0_7_i_da_d_iff;
  xt_rsc_1_23_i_qa_d <= xt_rsc_1_23_i_qa_d_1;

  xt_rsc_1_24_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_319_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_1_24_i_qa,
      wea => xt_rsc_1_24_wea,
      da => xt_rsc_1_24_i_da,
      adra => xt_rsc_1_24_i_adra,
      adra_d => xt_rsc_1_24_i_adra_d,
      da_d => xt_rsc_1_24_i_da_d,
      qa_d => xt_rsc_1_24_i_qa_d_1,
      wea_d => xt_rsc_1_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_16_i_wea_d_iff
    );
  xt_rsc_1_24_i_qa <= xt_rsc_1_24_qa;
  xt_rsc_1_24_da <= xt_rsc_1_24_i_da;
  xt_rsc_1_24_adra <= xt_rsc_1_24_i_adra;
  xt_rsc_1_24_i_adra_d <= xt_rsc_0_8_i_adra_d_iff;
  xt_rsc_1_24_i_da_d <= xt_rsc_0_8_i_da_d_iff;
  xt_rsc_1_24_i_qa_d <= xt_rsc_1_24_i_qa_d_1;

  xt_rsc_1_25_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_320_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_1_25_i_qa,
      wea => xt_rsc_1_25_wea,
      da => xt_rsc_1_25_i_da,
      adra => xt_rsc_1_25_i_adra,
      adra_d => xt_rsc_1_25_i_adra_d,
      da_d => xt_rsc_1_25_i_da_d,
      qa_d => xt_rsc_1_25_i_qa_d_1,
      wea_d => xt_rsc_1_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_16_i_wea_d_iff
    );
  xt_rsc_1_25_i_qa <= xt_rsc_1_25_qa;
  xt_rsc_1_25_da <= xt_rsc_1_25_i_da;
  xt_rsc_1_25_adra <= xt_rsc_1_25_i_adra;
  xt_rsc_1_25_i_adra_d <= xt_rsc_0_9_i_adra_d_iff;
  xt_rsc_1_25_i_da_d <= xt_rsc_0_9_i_da_d_iff;
  xt_rsc_1_25_i_qa_d <= xt_rsc_1_25_i_qa_d_1;

  xt_rsc_1_26_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_321_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_1_26_i_qa,
      wea => xt_rsc_1_26_wea,
      da => xt_rsc_1_26_i_da,
      adra => xt_rsc_1_26_i_adra,
      adra_d => xt_rsc_1_26_i_adra_d,
      da_d => xt_rsc_1_26_i_da_d,
      qa_d => xt_rsc_1_26_i_qa_d_1,
      wea_d => xt_rsc_1_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_16_i_wea_d_iff
    );
  xt_rsc_1_26_i_qa <= xt_rsc_1_26_qa;
  xt_rsc_1_26_da <= xt_rsc_1_26_i_da;
  xt_rsc_1_26_adra <= xt_rsc_1_26_i_adra;
  xt_rsc_1_26_i_adra_d <= xt_rsc_0_10_i_adra_d_iff;
  xt_rsc_1_26_i_da_d <= xt_rsc_0_10_i_da_d_iff;
  xt_rsc_1_26_i_qa_d <= xt_rsc_1_26_i_qa_d_1;

  xt_rsc_1_27_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_322_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_1_27_i_qa,
      wea => xt_rsc_1_27_wea,
      da => xt_rsc_1_27_i_da,
      adra => xt_rsc_1_27_i_adra,
      adra_d => xt_rsc_1_27_i_adra_d,
      da_d => xt_rsc_1_27_i_da_d,
      qa_d => xt_rsc_1_27_i_qa_d_1,
      wea_d => xt_rsc_1_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_16_i_wea_d_iff
    );
  xt_rsc_1_27_i_qa <= xt_rsc_1_27_qa;
  xt_rsc_1_27_da <= xt_rsc_1_27_i_da;
  xt_rsc_1_27_adra <= xt_rsc_1_27_i_adra;
  xt_rsc_1_27_i_adra_d <= xt_rsc_0_11_i_adra_d_iff;
  xt_rsc_1_27_i_da_d <= xt_rsc_0_11_i_da_d_iff;
  xt_rsc_1_27_i_qa_d <= xt_rsc_1_27_i_qa_d_1;

  xt_rsc_1_28_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_323_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_1_28_i_qa,
      wea => xt_rsc_1_28_wea,
      da => xt_rsc_1_28_i_da,
      adra => xt_rsc_1_28_i_adra,
      adra_d => xt_rsc_1_28_i_adra_d,
      da_d => xt_rsc_1_28_i_da_d,
      qa_d => xt_rsc_1_28_i_qa_d_1,
      wea_d => xt_rsc_1_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_16_i_wea_d_iff
    );
  xt_rsc_1_28_i_qa <= xt_rsc_1_28_qa;
  xt_rsc_1_28_da <= xt_rsc_1_28_i_da;
  xt_rsc_1_28_adra <= xt_rsc_1_28_i_adra;
  xt_rsc_1_28_i_adra_d <= xt_rsc_0_12_i_adra_d_iff;
  xt_rsc_1_28_i_da_d <= xt_rsc_0_12_i_da_d_iff;
  xt_rsc_1_28_i_qa_d <= xt_rsc_1_28_i_qa_d_1;

  xt_rsc_1_29_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_324_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_1_29_i_qa,
      wea => xt_rsc_1_29_wea,
      da => xt_rsc_1_29_i_da,
      adra => xt_rsc_1_29_i_adra,
      adra_d => xt_rsc_1_29_i_adra_d,
      da_d => xt_rsc_1_29_i_da_d,
      qa_d => xt_rsc_1_29_i_qa_d_1,
      wea_d => xt_rsc_1_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_16_i_wea_d_iff
    );
  xt_rsc_1_29_i_qa <= xt_rsc_1_29_qa;
  xt_rsc_1_29_da <= xt_rsc_1_29_i_da;
  xt_rsc_1_29_adra <= xt_rsc_1_29_i_adra;
  xt_rsc_1_29_i_adra_d <= xt_rsc_0_13_i_adra_d_iff;
  xt_rsc_1_29_i_da_d <= xt_rsc_0_13_i_da_d_iff;
  xt_rsc_1_29_i_qa_d <= xt_rsc_1_29_i_qa_d_1;

  xt_rsc_1_30_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_325_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_1_30_i_qa,
      wea => xt_rsc_1_30_wea,
      da => xt_rsc_1_30_i_da,
      adra => xt_rsc_1_30_i_adra,
      adra_d => xt_rsc_1_30_i_adra_d,
      da_d => xt_rsc_1_30_i_da_d,
      qa_d => xt_rsc_1_30_i_qa_d_1,
      wea_d => xt_rsc_1_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_16_i_wea_d_iff
    );
  xt_rsc_1_30_i_qa <= xt_rsc_1_30_qa;
  xt_rsc_1_30_da <= xt_rsc_1_30_i_da;
  xt_rsc_1_30_adra <= xt_rsc_1_30_i_adra;
  xt_rsc_1_30_i_adra_d <= xt_rsc_0_14_i_adra_d_iff;
  xt_rsc_1_30_i_da_d <= xt_rsc_0_14_i_da_d_iff;
  xt_rsc_1_30_i_qa_d <= xt_rsc_1_30_i_qa_d_1;

  xt_rsc_1_31_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_326_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_1_31_i_qa,
      wea => xt_rsc_1_31_wea,
      da => xt_rsc_1_31_i_da,
      adra => xt_rsc_1_31_i_adra,
      adra_d => xt_rsc_1_31_i_adra_d,
      da_d => xt_rsc_1_31_i_da_d,
      qa_d => xt_rsc_1_31_i_qa_d_1,
      wea_d => xt_rsc_1_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_16_i_wea_d_iff
    );
  xt_rsc_1_31_i_qa <= xt_rsc_1_31_qa;
  xt_rsc_1_31_da <= xt_rsc_1_31_i_da;
  xt_rsc_1_31_adra <= xt_rsc_1_31_i_adra;
  xt_rsc_1_31_i_adra_d <= xt_rsc_0_15_i_adra_d_iff;
  xt_rsc_1_31_i_da_d <= xt_rsc_0_15_i_da_d_iff;
  xt_rsc_1_31_i_qa_d <= xt_rsc_1_31_i_qa_d_1;

  xt_rsc_2_0_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_327_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_2_0_i_qa,
      wea => xt_rsc_2_0_wea,
      da => xt_rsc_2_0_i_da,
      adra => xt_rsc_2_0_i_adra,
      adra_d => xt_rsc_2_0_i_adra_d,
      da_d => xt_rsc_2_0_i_da_d,
      qa_d => xt_rsc_2_0_i_qa_d_1,
      wea_d => xt_rsc_2_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_2_0_i_wea_d_iff
    );
  xt_rsc_2_0_i_qa <= xt_rsc_2_0_qa;
  xt_rsc_2_0_da <= xt_rsc_2_0_i_da;
  xt_rsc_2_0_adra <= xt_rsc_2_0_i_adra;
  xt_rsc_2_0_i_adra_d <= xt_rsc_0_0_i_adra_d_iff;
  xt_rsc_2_0_i_da_d <= xt_rsc_0_0_i_da_d_iff;
  xt_rsc_2_0_i_qa_d <= xt_rsc_2_0_i_qa_d_1;

  xt_rsc_2_1_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_328_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_2_1_i_qa,
      wea => xt_rsc_2_1_wea,
      da => xt_rsc_2_1_i_da,
      adra => xt_rsc_2_1_i_adra,
      adra_d => xt_rsc_2_1_i_adra_d,
      da_d => xt_rsc_2_1_i_da_d,
      qa_d => xt_rsc_2_1_i_qa_d_1,
      wea_d => xt_rsc_2_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_2_0_i_wea_d_iff
    );
  xt_rsc_2_1_i_qa <= xt_rsc_2_1_qa;
  xt_rsc_2_1_da <= xt_rsc_2_1_i_da;
  xt_rsc_2_1_adra <= xt_rsc_2_1_i_adra;
  xt_rsc_2_1_i_adra_d <= xt_rsc_0_1_i_adra_d_iff;
  xt_rsc_2_1_i_da_d <= xt_rsc_0_1_i_da_d_iff;
  xt_rsc_2_1_i_qa_d <= xt_rsc_2_1_i_qa_d_1;

  xt_rsc_2_2_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_329_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_2_2_i_qa,
      wea => xt_rsc_2_2_wea,
      da => xt_rsc_2_2_i_da,
      adra => xt_rsc_2_2_i_adra,
      adra_d => xt_rsc_2_2_i_adra_d,
      da_d => xt_rsc_2_2_i_da_d,
      qa_d => xt_rsc_2_2_i_qa_d_1,
      wea_d => xt_rsc_2_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_2_0_i_wea_d_iff
    );
  xt_rsc_2_2_i_qa <= xt_rsc_2_2_qa;
  xt_rsc_2_2_da <= xt_rsc_2_2_i_da;
  xt_rsc_2_2_adra <= xt_rsc_2_2_i_adra;
  xt_rsc_2_2_i_adra_d <= xt_rsc_0_2_i_adra_d_iff;
  xt_rsc_2_2_i_da_d <= xt_rsc_0_2_i_da_d_iff;
  xt_rsc_2_2_i_qa_d <= xt_rsc_2_2_i_qa_d_1;

  xt_rsc_2_3_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_330_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_2_3_i_qa,
      wea => xt_rsc_2_3_wea,
      da => xt_rsc_2_3_i_da,
      adra => xt_rsc_2_3_i_adra,
      adra_d => xt_rsc_2_3_i_adra_d,
      da_d => xt_rsc_2_3_i_da_d,
      qa_d => xt_rsc_2_3_i_qa_d_1,
      wea_d => xt_rsc_2_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_2_0_i_wea_d_iff
    );
  xt_rsc_2_3_i_qa <= xt_rsc_2_3_qa;
  xt_rsc_2_3_da <= xt_rsc_2_3_i_da;
  xt_rsc_2_3_adra <= xt_rsc_2_3_i_adra;
  xt_rsc_2_3_i_adra_d <= xt_rsc_0_3_i_adra_d_iff;
  xt_rsc_2_3_i_da_d <= xt_rsc_0_3_i_da_d_iff;
  xt_rsc_2_3_i_qa_d <= xt_rsc_2_3_i_qa_d_1;

  xt_rsc_2_4_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_331_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_2_4_i_qa,
      wea => xt_rsc_2_4_wea,
      da => xt_rsc_2_4_i_da,
      adra => xt_rsc_2_4_i_adra,
      adra_d => xt_rsc_2_4_i_adra_d,
      da_d => xt_rsc_2_4_i_da_d,
      qa_d => xt_rsc_2_4_i_qa_d_1,
      wea_d => xt_rsc_2_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_2_0_i_wea_d_iff
    );
  xt_rsc_2_4_i_qa <= xt_rsc_2_4_qa;
  xt_rsc_2_4_da <= xt_rsc_2_4_i_da;
  xt_rsc_2_4_adra <= xt_rsc_2_4_i_adra;
  xt_rsc_2_4_i_adra_d <= xt_rsc_0_4_i_adra_d_iff;
  xt_rsc_2_4_i_da_d <= xt_rsc_0_4_i_da_d_iff;
  xt_rsc_2_4_i_qa_d <= xt_rsc_2_4_i_qa_d_1;

  xt_rsc_2_5_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_332_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_2_5_i_qa,
      wea => xt_rsc_2_5_wea,
      da => xt_rsc_2_5_i_da,
      adra => xt_rsc_2_5_i_adra,
      adra_d => xt_rsc_2_5_i_adra_d,
      da_d => xt_rsc_2_5_i_da_d,
      qa_d => xt_rsc_2_5_i_qa_d_1,
      wea_d => xt_rsc_2_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_2_0_i_wea_d_iff
    );
  xt_rsc_2_5_i_qa <= xt_rsc_2_5_qa;
  xt_rsc_2_5_da <= xt_rsc_2_5_i_da;
  xt_rsc_2_5_adra <= xt_rsc_2_5_i_adra;
  xt_rsc_2_5_i_adra_d <= xt_rsc_0_5_i_adra_d_iff;
  xt_rsc_2_5_i_da_d <= xt_rsc_0_5_i_da_d_iff;
  xt_rsc_2_5_i_qa_d <= xt_rsc_2_5_i_qa_d_1;

  xt_rsc_2_6_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_333_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_2_6_i_qa,
      wea => xt_rsc_2_6_wea,
      da => xt_rsc_2_6_i_da,
      adra => xt_rsc_2_6_i_adra,
      adra_d => xt_rsc_2_6_i_adra_d,
      da_d => xt_rsc_2_6_i_da_d,
      qa_d => xt_rsc_2_6_i_qa_d_1,
      wea_d => xt_rsc_2_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_2_0_i_wea_d_iff
    );
  xt_rsc_2_6_i_qa <= xt_rsc_2_6_qa;
  xt_rsc_2_6_da <= xt_rsc_2_6_i_da;
  xt_rsc_2_6_adra <= xt_rsc_2_6_i_adra;
  xt_rsc_2_6_i_adra_d <= xt_rsc_0_6_i_adra_d_iff;
  xt_rsc_2_6_i_da_d <= xt_rsc_0_6_i_da_d_iff;
  xt_rsc_2_6_i_qa_d <= xt_rsc_2_6_i_qa_d_1;

  xt_rsc_2_7_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_334_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_2_7_i_qa,
      wea => xt_rsc_2_7_wea,
      da => xt_rsc_2_7_i_da,
      adra => xt_rsc_2_7_i_adra,
      adra_d => xt_rsc_2_7_i_adra_d,
      da_d => xt_rsc_2_7_i_da_d,
      qa_d => xt_rsc_2_7_i_qa_d_1,
      wea_d => xt_rsc_2_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_2_0_i_wea_d_iff
    );
  xt_rsc_2_7_i_qa <= xt_rsc_2_7_qa;
  xt_rsc_2_7_da <= xt_rsc_2_7_i_da;
  xt_rsc_2_7_adra <= xt_rsc_2_7_i_adra;
  xt_rsc_2_7_i_adra_d <= xt_rsc_0_7_i_adra_d_iff;
  xt_rsc_2_7_i_da_d <= xt_rsc_0_7_i_da_d_iff;
  xt_rsc_2_7_i_qa_d <= xt_rsc_2_7_i_qa_d_1;

  xt_rsc_2_8_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_335_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_2_8_i_qa,
      wea => xt_rsc_2_8_wea,
      da => xt_rsc_2_8_i_da,
      adra => xt_rsc_2_8_i_adra,
      adra_d => xt_rsc_2_8_i_adra_d,
      da_d => xt_rsc_2_8_i_da_d,
      qa_d => xt_rsc_2_8_i_qa_d_1,
      wea_d => xt_rsc_2_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_2_0_i_wea_d_iff
    );
  xt_rsc_2_8_i_qa <= xt_rsc_2_8_qa;
  xt_rsc_2_8_da <= xt_rsc_2_8_i_da;
  xt_rsc_2_8_adra <= xt_rsc_2_8_i_adra;
  xt_rsc_2_8_i_adra_d <= xt_rsc_0_8_i_adra_d_iff;
  xt_rsc_2_8_i_da_d <= xt_rsc_0_8_i_da_d_iff;
  xt_rsc_2_8_i_qa_d <= xt_rsc_2_8_i_qa_d_1;

  xt_rsc_2_9_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_336_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_2_9_i_qa,
      wea => xt_rsc_2_9_wea,
      da => xt_rsc_2_9_i_da,
      adra => xt_rsc_2_9_i_adra,
      adra_d => xt_rsc_2_9_i_adra_d,
      da_d => xt_rsc_2_9_i_da_d,
      qa_d => xt_rsc_2_9_i_qa_d_1,
      wea_d => xt_rsc_2_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_2_0_i_wea_d_iff
    );
  xt_rsc_2_9_i_qa <= xt_rsc_2_9_qa;
  xt_rsc_2_9_da <= xt_rsc_2_9_i_da;
  xt_rsc_2_9_adra <= xt_rsc_2_9_i_adra;
  xt_rsc_2_9_i_adra_d <= xt_rsc_0_9_i_adra_d_iff;
  xt_rsc_2_9_i_da_d <= xt_rsc_0_9_i_da_d_iff;
  xt_rsc_2_9_i_qa_d <= xt_rsc_2_9_i_qa_d_1;

  xt_rsc_2_10_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_337_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_2_10_i_qa,
      wea => xt_rsc_2_10_wea,
      da => xt_rsc_2_10_i_da,
      adra => xt_rsc_2_10_i_adra,
      adra_d => xt_rsc_2_10_i_adra_d,
      da_d => xt_rsc_2_10_i_da_d,
      qa_d => xt_rsc_2_10_i_qa_d_1,
      wea_d => xt_rsc_2_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_2_0_i_wea_d_iff
    );
  xt_rsc_2_10_i_qa <= xt_rsc_2_10_qa;
  xt_rsc_2_10_da <= xt_rsc_2_10_i_da;
  xt_rsc_2_10_adra <= xt_rsc_2_10_i_adra;
  xt_rsc_2_10_i_adra_d <= xt_rsc_0_10_i_adra_d_iff;
  xt_rsc_2_10_i_da_d <= xt_rsc_0_10_i_da_d_iff;
  xt_rsc_2_10_i_qa_d <= xt_rsc_2_10_i_qa_d_1;

  xt_rsc_2_11_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_338_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_2_11_i_qa,
      wea => xt_rsc_2_11_wea,
      da => xt_rsc_2_11_i_da,
      adra => xt_rsc_2_11_i_adra,
      adra_d => xt_rsc_2_11_i_adra_d,
      da_d => xt_rsc_2_11_i_da_d,
      qa_d => xt_rsc_2_11_i_qa_d_1,
      wea_d => xt_rsc_2_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_2_0_i_wea_d_iff
    );
  xt_rsc_2_11_i_qa <= xt_rsc_2_11_qa;
  xt_rsc_2_11_da <= xt_rsc_2_11_i_da;
  xt_rsc_2_11_adra <= xt_rsc_2_11_i_adra;
  xt_rsc_2_11_i_adra_d <= xt_rsc_0_11_i_adra_d_iff;
  xt_rsc_2_11_i_da_d <= xt_rsc_0_11_i_da_d_iff;
  xt_rsc_2_11_i_qa_d <= xt_rsc_2_11_i_qa_d_1;

  xt_rsc_2_12_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_339_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_2_12_i_qa,
      wea => xt_rsc_2_12_wea,
      da => xt_rsc_2_12_i_da,
      adra => xt_rsc_2_12_i_adra,
      adra_d => xt_rsc_2_12_i_adra_d,
      da_d => xt_rsc_2_12_i_da_d,
      qa_d => xt_rsc_2_12_i_qa_d_1,
      wea_d => xt_rsc_2_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_2_0_i_wea_d_iff
    );
  xt_rsc_2_12_i_qa <= xt_rsc_2_12_qa;
  xt_rsc_2_12_da <= xt_rsc_2_12_i_da;
  xt_rsc_2_12_adra <= xt_rsc_2_12_i_adra;
  xt_rsc_2_12_i_adra_d <= xt_rsc_0_12_i_adra_d_iff;
  xt_rsc_2_12_i_da_d <= xt_rsc_0_12_i_da_d_iff;
  xt_rsc_2_12_i_qa_d <= xt_rsc_2_12_i_qa_d_1;

  xt_rsc_2_13_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_340_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_2_13_i_qa,
      wea => xt_rsc_2_13_wea,
      da => xt_rsc_2_13_i_da,
      adra => xt_rsc_2_13_i_adra,
      adra_d => xt_rsc_2_13_i_adra_d,
      da_d => xt_rsc_2_13_i_da_d,
      qa_d => xt_rsc_2_13_i_qa_d_1,
      wea_d => xt_rsc_2_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_2_0_i_wea_d_iff
    );
  xt_rsc_2_13_i_qa <= xt_rsc_2_13_qa;
  xt_rsc_2_13_da <= xt_rsc_2_13_i_da;
  xt_rsc_2_13_adra <= xt_rsc_2_13_i_adra;
  xt_rsc_2_13_i_adra_d <= xt_rsc_0_13_i_adra_d_iff;
  xt_rsc_2_13_i_da_d <= xt_rsc_0_13_i_da_d_iff;
  xt_rsc_2_13_i_qa_d <= xt_rsc_2_13_i_qa_d_1;

  xt_rsc_2_14_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_341_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_2_14_i_qa,
      wea => xt_rsc_2_14_wea,
      da => xt_rsc_2_14_i_da,
      adra => xt_rsc_2_14_i_adra,
      adra_d => xt_rsc_2_14_i_adra_d,
      da_d => xt_rsc_2_14_i_da_d,
      qa_d => xt_rsc_2_14_i_qa_d_1,
      wea_d => xt_rsc_2_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_2_0_i_wea_d_iff
    );
  xt_rsc_2_14_i_qa <= xt_rsc_2_14_qa;
  xt_rsc_2_14_da <= xt_rsc_2_14_i_da;
  xt_rsc_2_14_adra <= xt_rsc_2_14_i_adra;
  xt_rsc_2_14_i_adra_d <= xt_rsc_0_14_i_adra_d_iff;
  xt_rsc_2_14_i_da_d <= xt_rsc_0_14_i_da_d_iff;
  xt_rsc_2_14_i_qa_d <= xt_rsc_2_14_i_qa_d_1;

  xt_rsc_2_15_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_342_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_2_15_i_qa,
      wea => xt_rsc_2_15_wea,
      da => xt_rsc_2_15_i_da,
      adra => xt_rsc_2_15_i_adra,
      adra_d => xt_rsc_2_15_i_adra_d,
      da_d => xt_rsc_2_15_i_da_d,
      qa_d => xt_rsc_2_15_i_qa_d_1,
      wea_d => xt_rsc_2_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_2_0_i_wea_d_iff
    );
  xt_rsc_2_15_i_qa <= xt_rsc_2_15_qa;
  xt_rsc_2_15_da <= xt_rsc_2_15_i_da;
  xt_rsc_2_15_adra <= xt_rsc_2_15_i_adra;
  xt_rsc_2_15_i_adra_d <= xt_rsc_0_15_i_adra_d_iff;
  xt_rsc_2_15_i_da_d <= xt_rsc_0_15_i_da_d_iff;
  xt_rsc_2_15_i_qa_d <= xt_rsc_2_15_i_qa_d_1;

  xt_rsc_2_16_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_343_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_2_16_i_qa,
      wea => xt_rsc_2_16_wea,
      da => xt_rsc_2_16_i_da,
      adra => xt_rsc_2_16_i_adra,
      adra_d => xt_rsc_2_16_i_adra_d,
      da_d => xt_rsc_2_16_i_da_d,
      qa_d => xt_rsc_2_16_i_qa_d_1,
      wea_d => xt_rsc_2_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_2_16_i_wea_d_iff
    );
  xt_rsc_2_16_i_qa <= xt_rsc_2_16_qa;
  xt_rsc_2_16_da <= xt_rsc_2_16_i_da;
  xt_rsc_2_16_adra <= xt_rsc_2_16_i_adra;
  xt_rsc_2_16_i_adra_d <= xt_rsc_0_0_i_adra_d_iff;
  xt_rsc_2_16_i_da_d <= xt_rsc_0_0_i_da_d_iff;
  xt_rsc_2_16_i_qa_d <= xt_rsc_2_16_i_qa_d_1;

  xt_rsc_2_17_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_344_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_2_17_i_qa,
      wea => xt_rsc_2_17_wea,
      da => xt_rsc_2_17_i_da,
      adra => xt_rsc_2_17_i_adra,
      adra_d => xt_rsc_2_17_i_adra_d,
      da_d => xt_rsc_2_17_i_da_d,
      qa_d => xt_rsc_2_17_i_qa_d_1,
      wea_d => xt_rsc_2_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_2_16_i_wea_d_iff
    );
  xt_rsc_2_17_i_qa <= xt_rsc_2_17_qa;
  xt_rsc_2_17_da <= xt_rsc_2_17_i_da;
  xt_rsc_2_17_adra <= xt_rsc_2_17_i_adra;
  xt_rsc_2_17_i_adra_d <= xt_rsc_0_1_i_adra_d_iff;
  xt_rsc_2_17_i_da_d <= xt_rsc_0_1_i_da_d_iff;
  xt_rsc_2_17_i_qa_d <= xt_rsc_2_17_i_qa_d_1;

  xt_rsc_2_18_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_345_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_2_18_i_qa,
      wea => xt_rsc_2_18_wea,
      da => xt_rsc_2_18_i_da,
      adra => xt_rsc_2_18_i_adra,
      adra_d => xt_rsc_2_18_i_adra_d,
      da_d => xt_rsc_2_18_i_da_d,
      qa_d => xt_rsc_2_18_i_qa_d_1,
      wea_d => xt_rsc_2_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_2_16_i_wea_d_iff
    );
  xt_rsc_2_18_i_qa <= xt_rsc_2_18_qa;
  xt_rsc_2_18_da <= xt_rsc_2_18_i_da;
  xt_rsc_2_18_adra <= xt_rsc_2_18_i_adra;
  xt_rsc_2_18_i_adra_d <= xt_rsc_0_2_i_adra_d_iff;
  xt_rsc_2_18_i_da_d <= xt_rsc_0_2_i_da_d_iff;
  xt_rsc_2_18_i_qa_d <= xt_rsc_2_18_i_qa_d_1;

  xt_rsc_2_19_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_346_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_2_19_i_qa,
      wea => xt_rsc_2_19_wea,
      da => xt_rsc_2_19_i_da,
      adra => xt_rsc_2_19_i_adra,
      adra_d => xt_rsc_2_19_i_adra_d,
      da_d => xt_rsc_2_19_i_da_d,
      qa_d => xt_rsc_2_19_i_qa_d_1,
      wea_d => xt_rsc_2_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_2_16_i_wea_d_iff
    );
  xt_rsc_2_19_i_qa <= xt_rsc_2_19_qa;
  xt_rsc_2_19_da <= xt_rsc_2_19_i_da;
  xt_rsc_2_19_adra <= xt_rsc_2_19_i_adra;
  xt_rsc_2_19_i_adra_d <= xt_rsc_0_3_i_adra_d_iff;
  xt_rsc_2_19_i_da_d <= xt_rsc_0_3_i_da_d_iff;
  xt_rsc_2_19_i_qa_d <= xt_rsc_2_19_i_qa_d_1;

  xt_rsc_2_20_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_347_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_2_20_i_qa,
      wea => xt_rsc_2_20_wea,
      da => xt_rsc_2_20_i_da,
      adra => xt_rsc_2_20_i_adra,
      adra_d => xt_rsc_2_20_i_adra_d,
      da_d => xt_rsc_2_20_i_da_d,
      qa_d => xt_rsc_2_20_i_qa_d_1,
      wea_d => xt_rsc_2_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_2_16_i_wea_d_iff
    );
  xt_rsc_2_20_i_qa <= xt_rsc_2_20_qa;
  xt_rsc_2_20_da <= xt_rsc_2_20_i_da;
  xt_rsc_2_20_adra <= xt_rsc_2_20_i_adra;
  xt_rsc_2_20_i_adra_d <= xt_rsc_0_4_i_adra_d_iff;
  xt_rsc_2_20_i_da_d <= xt_rsc_0_4_i_da_d_iff;
  xt_rsc_2_20_i_qa_d <= xt_rsc_2_20_i_qa_d_1;

  xt_rsc_2_21_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_348_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_2_21_i_qa,
      wea => xt_rsc_2_21_wea,
      da => xt_rsc_2_21_i_da,
      adra => xt_rsc_2_21_i_adra,
      adra_d => xt_rsc_2_21_i_adra_d,
      da_d => xt_rsc_2_21_i_da_d,
      qa_d => xt_rsc_2_21_i_qa_d_1,
      wea_d => xt_rsc_2_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_2_16_i_wea_d_iff
    );
  xt_rsc_2_21_i_qa <= xt_rsc_2_21_qa;
  xt_rsc_2_21_da <= xt_rsc_2_21_i_da;
  xt_rsc_2_21_adra <= xt_rsc_2_21_i_adra;
  xt_rsc_2_21_i_adra_d <= xt_rsc_0_5_i_adra_d_iff;
  xt_rsc_2_21_i_da_d <= xt_rsc_0_5_i_da_d_iff;
  xt_rsc_2_21_i_qa_d <= xt_rsc_2_21_i_qa_d_1;

  xt_rsc_2_22_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_349_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_2_22_i_qa,
      wea => xt_rsc_2_22_wea,
      da => xt_rsc_2_22_i_da,
      adra => xt_rsc_2_22_i_adra,
      adra_d => xt_rsc_2_22_i_adra_d,
      da_d => xt_rsc_2_22_i_da_d,
      qa_d => xt_rsc_2_22_i_qa_d_1,
      wea_d => xt_rsc_2_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_2_16_i_wea_d_iff
    );
  xt_rsc_2_22_i_qa <= xt_rsc_2_22_qa;
  xt_rsc_2_22_da <= xt_rsc_2_22_i_da;
  xt_rsc_2_22_adra <= xt_rsc_2_22_i_adra;
  xt_rsc_2_22_i_adra_d <= xt_rsc_0_6_i_adra_d_iff;
  xt_rsc_2_22_i_da_d <= xt_rsc_0_6_i_da_d_iff;
  xt_rsc_2_22_i_qa_d <= xt_rsc_2_22_i_qa_d_1;

  xt_rsc_2_23_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_350_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_2_23_i_qa,
      wea => xt_rsc_2_23_wea,
      da => xt_rsc_2_23_i_da,
      adra => xt_rsc_2_23_i_adra,
      adra_d => xt_rsc_2_23_i_adra_d,
      da_d => xt_rsc_2_23_i_da_d,
      qa_d => xt_rsc_2_23_i_qa_d_1,
      wea_d => xt_rsc_2_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_2_16_i_wea_d_iff
    );
  xt_rsc_2_23_i_qa <= xt_rsc_2_23_qa;
  xt_rsc_2_23_da <= xt_rsc_2_23_i_da;
  xt_rsc_2_23_adra <= xt_rsc_2_23_i_adra;
  xt_rsc_2_23_i_adra_d <= xt_rsc_0_7_i_adra_d_iff;
  xt_rsc_2_23_i_da_d <= xt_rsc_0_7_i_da_d_iff;
  xt_rsc_2_23_i_qa_d <= xt_rsc_2_23_i_qa_d_1;

  xt_rsc_2_24_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_351_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_2_24_i_qa,
      wea => xt_rsc_2_24_wea,
      da => xt_rsc_2_24_i_da,
      adra => xt_rsc_2_24_i_adra,
      adra_d => xt_rsc_2_24_i_adra_d,
      da_d => xt_rsc_2_24_i_da_d,
      qa_d => xt_rsc_2_24_i_qa_d_1,
      wea_d => xt_rsc_2_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_2_16_i_wea_d_iff
    );
  xt_rsc_2_24_i_qa <= xt_rsc_2_24_qa;
  xt_rsc_2_24_da <= xt_rsc_2_24_i_da;
  xt_rsc_2_24_adra <= xt_rsc_2_24_i_adra;
  xt_rsc_2_24_i_adra_d <= xt_rsc_0_8_i_adra_d_iff;
  xt_rsc_2_24_i_da_d <= xt_rsc_0_8_i_da_d_iff;
  xt_rsc_2_24_i_qa_d <= xt_rsc_2_24_i_qa_d_1;

  xt_rsc_2_25_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_352_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_2_25_i_qa,
      wea => xt_rsc_2_25_wea,
      da => xt_rsc_2_25_i_da,
      adra => xt_rsc_2_25_i_adra,
      adra_d => xt_rsc_2_25_i_adra_d,
      da_d => xt_rsc_2_25_i_da_d,
      qa_d => xt_rsc_2_25_i_qa_d_1,
      wea_d => xt_rsc_2_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_2_16_i_wea_d_iff
    );
  xt_rsc_2_25_i_qa <= xt_rsc_2_25_qa;
  xt_rsc_2_25_da <= xt_rsc_2_25_i_da;
  xt_rsc_2_25_adra <= xt_rsc_2_25_i_adra;
  xt_rsc_2_25_i_adra_d <= xt_rsc_0_9_i_adra_d_iff;
  xt_rsc_2_25_i_da_d <= xt_rsc_0_9_i_da_d_iff;
  xt_rsc_2_25_i_qa_d <= xt_rsc_2_25_i_qa_d_1;

  xt_rsc_2_26_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_353_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_2_26_i_qa,
      wea => xt_rsc_2_26_wea,
      da => xt_rsc_2_26_i_da,
      adra => xt_rsc_2_26_i_adra,
      adra_d => xt_rsc_2_26_i_adra_d,
      da_d => xt_rsc_2_26_i_da_d,
      qa_d => xt_rsc_2_26_i_qa_d_1,
      wea_d => xt_rsc_2_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_2_16_i_wea_d_iff
    );
  xt_rsc_2_26_i_qa <= xt_rsc_2_26_qa;
  xt_rsc_2_26_da <= xt_rsc_2_26_i_da;
  xt_rsc_2_26_adra <= xt_rsc_2_26_i_adra;
  xt_rsc_2_26_i_adra_d <= xt_rsc_0_10_i_adra_d_iff;
  xt_rsc_2_26_i_da_d <= xt_rsc_0_10_i_da_d_iff;
  xt_rsc_2_26_i_qa_d <= xt_rsc_2_26_i_qa_d_1;

  xt_rsc_2_27_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_354_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_2_27_i_qa,
      wea => xt_rsc_2_27_wea,
      da => xt_rsc_2_27_i_da,
      adra => xt_rsc_2_27_i_adra,
      adra_d => xt_rsc_2_27_i_adra_d,
      da_d => xt_rsc_2_27_i_da_d,
      qa_d => xt_rsc_2_27_i_qa_d_1,
      wea_d => xt_rsc_2_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_2_16_i_wea_d_iff
    );
  xt_rsc_2_27_i_qa <= xt_rsc_2_27_qa;
  xt_rsc_2_27_da <= xt_rsc_2_27_i_da;
  xt_rsc_2_27_adra <= xt_rsc_2_27_i_adra;
  xt_rsc_2_27_i_adra_d <= xt_rsc_0_11_i_adra_d_iff;
  xt_rsc_2_27_i_da_d <= xt_rsc_0_11_i_da_d_iff;
  xt_rsc_2_27_i_qa_d <= xt_rsc_2_27_i_qa_d_1;

  xt_rsc_2_28_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_355_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_2_28_i_qa,
      wea => xt_rsc_2_28_wea,
      da => xt_rsc_2_28_i_da,
      adra => xt_rsc_2_28_i_adra,
      adra_d => xt_rsc_2_28_i_adra_d,
      da_d => xt_rsc_2_28_i_da_d,
      qa_d => xt_rsc_2_28_i_qa_d_1,
      wea_d => xt_rsc_2_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_2_16_i_wea_d_iff
    );
  xt_rsc_2_28_i_qa <= xt_rsc_2_28_qa;
  xt_rsc_2_28_da <= xt_rsc_2_28_i_da;
  xt_rsc_2_28_adra <= xt_rsc_2_28_i_adra;
  xt_rsc_2_28_i_adra_d <= xt_rsc_0_12_i_adra_d_iff;
  xt_rsc_2_28_i_da_d <= xt_rsc_0_12_i_da_d_iff;
  xt_rsc_2_28_i_qa_d <= xt_rsc_2_28_i_qa_d_1;

  xt_rsc_2_29_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_356_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_2_29_i_qa,
      wea => xt_rsc_2_29_wea,
      da => xt_rsc_2_29_i_da,
      adra => xt_rsc_2_29_i_adra,
      adra_d => xt_rsc_2_29_i_adra_d,
      da_d => xt_rsc_2_29_i_da_d,
      qa_d => xt_rsc_2_29_i_qa_d_1,
      wea_d => xt_rsc_2_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_2_16_i_wea_d_iff
    );
  xt_rsc_2_29_i_qa <= xt_rsc_2_29_qa;
  xt_rsc_2_29_da <= xt_rsc_2_29_i_da;
  xt_rsc_2_29_adra <= xt_rsc_2_29_i_adra;
  xt_rsc_2_29_i_adra_d <= xt_rsc_0_13_i_adra_d_iff;
  xt_rsc_2_29_i_da_d <= xt_rsc_0_13_i_da_d_iff;
  xt_rsc_2_29_i_qa_d <= xt_rsc_2_29_i_qa_d_1;

  xt_rsc_2_30_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_357_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_2_30_i_qa,
      wea => xt_rsc_2_30_wea,
      da => xt_rsc_2_30_i_da,
      adra => xt_rsc_2_30_i_adra,
      adra_d => xt_rsc_2_30_i_adra_d,
      da_d => xt_rsc_2_30_i_da_d,
      qa_d => xt_rsc_2_30_i_qa_d_1,
      wea_d => xt_rsc_2_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_2_16_i_wea_d_iff
    );
  xt_rsc_2_30_i_qa <= xt_rsc_2_30_qa;
  xt_rsc_2_30_da <= xt_rsc_2_30_i_da;
  xt_rsc_2_30_adra <= xt_rsc_2_30_i_adra;
  xt_rsc_2_30_i_adra_d <= xt_rsc_0_14_i_adra_d_iff;
  xt_rsc_2_30_i_da_d <= xt_rsc_0_14_i_da_d_iff;
  xt_rsc_2_30_i_qa_d <= xt_rsc_2_30_i_qa_d_1;

  xt_rsc_2_31_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_358_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_2_31_i_qa,
      wea => xt_rsc_2_31_wea,
      da => xt_rsc_2_31_i_da,
      adra => xt_rsc_2_31_i_adra,
      adra_d => xt_rsc_2_31_i_adra_d,
      da_d => xt_rsc_2_31_i_da_d,
      qa_d => xt_rsc_2_31_i_qa_d_1,
      wea_d => xt_rsc_2_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_2_16_i_wea_d_iff
    );
  xt_rsc_2_31_i_qa <= xt_rsc_2_31_qa;
  xt_rsc_2_31_da <= xt_rsc_2_31_i_da;
  xt_rsc_2_31_adra <= xt_rsc_2_31_i_adra;
  xt_rsc_2_31_i_adra_d <= xt_rsc_0_15_i_adra_d_iff;
  xt_rsc_2_31_i_da_d <= xt_rsc_0_15_i_da_d_iff;
  xt_rsc_2_31_i_qa_d <= xt_rsc_2_31_i_qa_d_1;

  xt_rsc_3_0_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_359_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_3_0_i_qa,
      wea => xt_rsc_3_0_wea,
      da => xt_rsc_3_0_i_da,
      adra => xt_rsc_3_0_i_adra,
      adra_d => xt_rsc_3_0_i_adra_d,
      da_d => xt_rsc_3_0_i_da_d,
      qa_d => xt_rsc_3_0_i_qa_d_1,
      wea_d => xt_rsc_3_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_3_0_i_wea_d_iff
    );
  xt_rsc_3_0_i_qa <= xt_rsc_3_0_qa;
  xt_rsc_3_0_da <= xt_rsc_3_0_i_da;
  xt_rsc_3_0_adra <= xt_rsc_3_0_i_adra;
  xt_rsc_3_0_i_adra_d <= xt_rsc_0_0_i_adra_d_iff;
  xt_rsc_3_0_i_da_d <= xt_rsc_0_0_i_da_d_iff;
  xt_rsc_3_0_i_qa_d <= xt_rsc_3_0_i_qa_d_1;

  xt_rsc_3_1_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_360_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_3_1_i_qa,
      wea => xt_rsc_3_1_wea,
      da => xt_rsc_3_1_i_da,
      adra => xt_rsc_3_1_i_adra,
      adra_d => xt_rsc_3_1_i_adra_d,
      da_d => xt_rsc_3_1_i_da_d,
      qa_d => xt_rsc_3_1_i_qa_d_1,
      wea_d => xt_rsc_3_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_3_0_i_wea_d_iff
    );
  xt_rsc_3_1_i_qa <= xt_rsc_3_1_qa;
  xt_rsc_3_1_da <= xt_rsc_3_1_i_da;
  xt_rsc_3_1_adra <= xt_rsc_3_1_i_adra;
  xt_rsc_3_1_i_adra_d <= xt_rsc_0_1_i_adra_d_iff;
  xt_rsc_3_1_i_da_d <= xt_rsc_0_1_i_da_d_iff;
  xt_rsc_3_1_i_qa_d <= xt_rsc_3_1_i_qa_d_1;

  xt_rsc_3_2_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_361_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_3_2_i_qa,
      wea => xt_rsc_3_2_wea,
      da => xt_rsc_3_2_i_da,
      adra => xt_rsc_3_2_i_adra,
      adra_d => xt_rsc_3_2_i_adra_d,
      da_d => xt_rsc_3_2_i_da_d,
      qa_d => xt_rsc_3_2_i_qa_d_1,
      wea_d => xt_rsc_3_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_3_0_i_wea_d_iff
    );
  xt_rsc_3_2_i_qa <= xt_rsc_3_2_qa;
  xt_rsc_3_2_da <= xt_rsc_3_2_i_da;
  xt_rsc_3_2_adra <= xt_rsc_3_2_i_adra;
  xt_rsc_3_2_i_adra_d <= xt_rsc_0_2_i_adra_d_iff;
  xt_rsc_3_2_i_da_d <= xt_rsc_0_2_i_da_d_iff;
  xt_rsc_3_2_i_qa_d <= xt_rsc_3_2_i_qa_d_1;

  xt_rsc_3_3_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_362_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_3_3_i_qa,
      wea => xt_rsc_3_3_wea,
      da => xt_rsc_3_3_i_da,
      adra => xt_rsc_3_3_i_adra,
      adra_d => xt_rsc_3_3_i_adra_d,
      da_d => xt_rsc_3_3_i_da_d,
      qa_d => xt_rsc_3_3_i_qa_d_1,
      wea_d => xt_rsc_3_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_3_0_i_wea_d_iff
    );
  xt_rsc_3_3_i_qa <= xt_rsc_3_3_qa;
  xt_rsc_3_3_da <= xt_rsc_3_3_i_da;
  xt_rsc_3_3_adra <= xt_rsc_3_3_i_adra;
  xt_rsc_3_3_i_adra_d <= xt_rsc_0_3_i_adra_d_iff;
  xt_rsc_3_3_i_da_d <= xt_rsc_0_3_i_da_d_iff;
  xt_rsc_3_3_i_qa_d <= xt_rsc_3_3_i_qa_d_1;

  xt_rsc_3_4_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_363_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_3_4_i_qa,
      wea => xt_rsc_3_4_wea,
      da => xt_rsc_3_4_i_da,
      adra => xt_rsc_3_4_i_adra,
      adra_d => xt_rsc_3_4_i_adra_d,
      da_d => xt_rsc_3_4_i_da_d,
      qa_d => xt_rsc_3_4_i_qa_d_1,
      wea_d => xt_rsc_3_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_3_0_i_wea_d_iff
    );
  xt_rsc_3_4_i_qa <= xt_rsc_3_4_qa;
  xt_rsc_3_4_da <= xt_rsc_3_4_i_da;
  xt_rsc_3_4_adra <= xt_rsc_3_4_i_adra;
  xt_rsc_3_4_i_adra_d <= xt_rsc_0_4_i_adra_d_iff;
  xt_rsc_3_4_i_da_d <= xt_rsc_0_4_i_da_d_iff;
  xt_rsc_3_4_i_qa_d <= xt_rsc_3_4_i_qa_d_1;

  xt_rsc_3_5_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_364_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_3_5_i_qa,
      wea => xt_rsc_3_5_wea,
      da => xt_rsc_3_5_i_da,
      adra => xt_rsc_3_5_i_adra,
      adra_d => xt_rsc_3_5_i_adra_d,
      da_d => xt_rsc_3_5_i_da_d,
      qa_d => xt_rsc_3_5_i_qa_d_1,
      wea_d => xt_rsc_3_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_3_0_i_wea_d_iff
    );
  xt_rsc_3_5_i_qa <= xt_rsc_3_5_qa;
  xt_rsc_3_5_da <= xt_rsc_3_5_i_da;
  xt_rsc_3_5_adra <= xt_rsc_3_5_i_adra;
  xt_rsc_3_5_i_adra_d <= xt_rsc_0_5_i_adra_d_iff;
  xt_rsc_3_5_i_da_d <= xt_rsc_0_5_i_da_d_iff;
  xt_rsc_3_5_i_qa_d <= xt_rsc_3_5_i_qa_d_1;

  xt_rsc_3_6_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_365_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_3_6_i_qa,
      wea => xt_rsc_3_6_wea,
      da => xt_rsc_3_6_i_da,
      adra => xt_rsc_3_6_i_adra,
      adra_d => xt_rsc_3_6_i_adra_d,
      da_d => xt_rsc_3_6_i_da_d,
      qa_d => xt_rsc_3_6_i_qa_d_1,
      wea_d => xt_rsc_3_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_3_0_i_wea_d_iff
    );
  xt_rsc_3_6_i_qa <= xt_rsc_3_6_qa;
  xt_rsc_3_6_da <= xt_rsc_3_6_i_da;
  xt_rsc_3_6_adra <= xt_rsc_3_6_i_adra;
  xt_rsc_3_6_i_adra_d <= xt_rsc_0_6_i_adra_d_iff;
  xt_rsc_3_6_i_da_d <= xt_rsc_0_6_i_da_d_iff;
  xt_rsc_3_6_i_qa_d <= xt_rsc_3_6_i_qa_d_1;

  xt_rsc_3_7_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_366_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_3_7_i_qa,
      wea => xt_rsc_3_7_wea,
      da => xt_rsc_3_7_i_da,
      adra => xt_rsc_3_7_i_adra,
      adra_d => xt_rsc_3_7_i_adra_d,
      da_d => xt_rsc_3_7_i_da_d,
      qa_d => xt_rsc_3_7_i_qa_d_1,
      wea_d => xt_rsc_3_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_3_0_i_wea_d_iff
    );
  xt_rsc_3_7_i_qa <= xt_rsc_3_7_qa;
  xt_rsc_3_7_da <= xt_rsc_3_7_i_da;
  xt_rsc_3_7_adra <= xt_rsc_3_7_i_adra;
  xt_rsc_3_7_i_adra_d <= xt_rsc_0_7_i_adra_d_iff;
  xt_rsc_3_7_i_da_d <= xt_rsc_0_7_i_da_d_iff;
  xt_rsc_3_7_i_qa_d <= xt_rsc_3_7_i_qa_d_1;

  xt_rsc_3_8_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_367_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_3_8_i_qa,
      wea => xt_rsc_3_8_wea,
      da => xt_rsc_3_8_i_da,
      adra => xt_rsc_3_8_i_adra,
      adra_d => xt_rsc_3_8_i_adra_d,
      da_d => xt_rsc_3_8_i_da_d,
      qa_d => xt_rsc_3_8_i_qa_d_1,
      wea_d => xt_rsc_3_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_3_0_i_wea_d_iff
    );
  xt_rsc_3_8_i_qa <= xt_rsc_3_8_qa;
  xt_rsc_3_8_da <= xt_rsc_3_8_i_da;
  xt_rsc_3_8_adra <= xt_rsc_3_8_i_adra;
  xt_rsc_3_8_i_adra_d <= xt_rsc_0_8_i_adra_d_iff;
  xt_rsc_3_8_i_da_d <= xt_rsc_0_8_i_da_d_iff;
  xt_rsc_3_8_i_qa_d <= xt_rsc_3_8_i_qa_d_1;

  xt_rsc_3_9_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_368_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_3_9_i_qa,
      wea => xt_rsc_3_9_wea,
      da => xt_rsc_3_9_i_da,
      adra => xt_rsc_3_9_i_adra,
      adra_d => xt_rsc_3_9_i_adra_d,
      da_d => xt_rsc_3_9_i_da_d,
      qa_d => xt_rsc_3_9_i_qa_d_1,
      wea_d => xt_rsc_3_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_3_0_i_wea_d_iff
    );
  xt_rsc_3_9_i_qa <= xt_rsc_3_9_qa;
  xt_rsc_3_9_da <= xt_rsc_3_9_i_da;
  xt_rsc_3_9_adra <= xt_rsc_3_9_i_adra;
  xt_rsc_3_9_i_adra_d <= xt_rsc_0_9_i_adra_d_iff;
  xt_rsc_3_9_i_da_d <= xt_rsc_0_9_i_da_d_iff;
  xt_rsc_3_9_i_qa_d <= xt_rsc_3_9_i_qa_d_1;

  xt_rsc_3_10_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_369_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_3_10_i_qa,
      wea => xt_rsc_3_10_wea,
      da => xt_rsc_3_10_i_da,
      adra => xt_rsc_3_10_i_adra,
      adra_d => xt_rsc_3_10_i_adra_d,
      da_d => xt_rsc_3_10_i_da_d,
      qa_d => xt_rsc_3_10_i_qa_d_1,
      wea_d => xt_rsc_3_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_3_0_i_wea_d_iff
    );
  xt_rsc_3_10_i_qa <= xt_rsc_3_10_qa;
  xt_rsc_3_10_da <= xt_rsc_3_10_i_da;
  xt_rsc_3_10_adra <= xt_rsc_3_10_i_adra;
  xt_rsc_3_10_i_adra_d <= xt_rsc_0_10_i_adra_d_iff;
  xt_rsc_3_10_i_da_d <= xt_rsc_0_10_i_da_d_iff;
  xt_rsc_3_10_i_qa_d <= xt_rsc_3_10_i_qa_d_1;

  xt_rsc_3_11_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_370_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_3_11_i_qa,
      wea => xt_rsc_3_11_wea,
      da => xt_rsc_3_11_i_da,
      adra => xt_rsc_3_11_i_adra,
      adra_d => xt_rsc_3_11_i_adra_d,
      da_d => xt_rsc_3_11_i_da_d,
      qa_d => xt_rsc_3_11_i_qa_d_1,
      wea_d => xt_rsc_3_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_3_0_i_wea_d_iff
    );
  xt_rsc_3_11_i_qa <= xt_rsc_3_11_qa;
  xt_rsc_3_11_da <= xt_rsc_3_11_i_da;
  xt_rsc_3_11_adra <= xt_rsc_3_11_i_adra;
  xt_rsc_3_11_i_adra_d <= xt_rsc_0_11_i_adra_d_iff;
  xt_rsc_3_11_i_da_d <= xt_rsc_0_11_i_da_d_iff;
  xt_rsc_3_11_i_qa_d <= xt_rsc_3_11_i_qa_d_1;

  xt_rsc_3_12_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_371_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_3_12_i_qa,
      wea => xt_rsc_3_12_wea,
      da => xt_rsc_3_12_i_da,
      adra => xt_rsc_3_12_i_adra,
      adra_d => xt_rsc_3_12_i_adra_d,
      da_d => xt_rsc_3_12_i_da_d,
      qa_d => xt_rsc_3_12_i_qa_d_1,
      wea_d => xt_rsc_3_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_3_0_i_wea_d_iff
    );
  xt_rsc_3_12_i_qa <= xt_rsc_3_12_qa;
  xt_rsc_3_12_da <= xt_rsc_3_12_i_da;
  xt_rsc_3_12_adra <= xt_rsc_3_12_i_adra;
  xt_rsc_3_12_i_adra_d <= xt_rsc_0_12_i_adra_d_iff;
  xt_rsc_3_12_i_da_d <= xt_rsc_0_12_i_da_d_iff;
  xt_rsc_3_12_i_qa_d <= xt_rsc_3_12_i_qa_d_1;

  xt_rsc_3_13_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_372_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_3_13_i_qa,
      wea => xt_rsc_3_13_wea,
      da => xt_rsc_3_13_i_da,
      adra => xt_rsc_3_13_i_adra,
      adra_d => xt_rsc_3_13_i_adra_d,
      da_d => xt_rsc_3_13_i_da_d,
      qa_d => xt_rsc_3_13_i_qa_d_1,
      wea_d => xt_rsc_3_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_3_0_i_wea_d_iff
    );
  xt_rsc_3_13_i_qa <= xt_rsc_3_13_qa;
  xt_rsc_3_13_da <= xt_rsc_3_13_i_da;
  xt_rsc_3_13_adra <= xt_rsc_3_13_i_adra;
  xt_rsc_3_13_i_adra_d <= xt_rsc_0_13_i_adra_d_iff;
  xt_rsc_3_13_i_da_d <= xt_rsc_0_13_i_da_d_iff;
  xt_rsc_3_13_i_qa_d <= xt_rsc_3_13_i_qa_d_1;

  xt_rsc_3_14_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_373_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_3_14_i_qa,
      wea => xt_rsc_3_14_wea,
      da => xt_rsc_3_14_i_da,
      adra => xt_rsc_3_14_i_adra,
      adra_d => xt_rsc_3_14_i_adra_d,
      da_d => xt_rsc_3_14_i_da_d,
      qa_d => xt_rsc_3_14_i_qa_d_1,
      wea_d => xt_rsc_3_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_3_0_i_wea_d_iff
    );
  xt_rsc_3_14_i_qa <= xt_rsc_3_14_qa;
  xt_rsc_3_14_da <= xt_rsc_3_14_i_da;
  xt_rsc_3_14_adra <= xt_rsc_3_14_i_adra;
  xt_rsc_3_14_i_adra_d <= xt_rsc_0_14_i_adra_d_iff;
  xt_rsc_3_14_i_da_d <= xt_rsc_0_14_i_da_d_iff;
  xt_rsc_3_14_i_qa_d <= xt_rsc_3_14_i_qa_d_1;

  xt_rsc_3_15_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_374_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_3_15_i_qa,
      wea => xt_rsc_3_15_wea,
      da => xt_rsc_3_15_i_da,
      adra => xt_rsc_3_15_i_adra,
      adra_d => xt_rsc_3_15_i_adra_d,
      da_d => xt_rsc_3_15_i_da_d,
      qa_d => xt_rsc_3_15_i_qa_d_1,
      wea_d => xt_rsc_3_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_3_0_i_wea_d_iff
    );
  xt_rsc_3_15_i_qa <= xt_rsc_3_15_qa;
  xt_rsc_3_15_da <= xt_rsc_3_15_i_da;
  xt_rsc_3_15_adra <= xt_rsc_3_15_i_adra;
  xt_rsc_3_15_i_adra_d <= xt_rsc_0_15_i_adra_d_iff;
  xt_rsc_3_15_i_da_d <= xt_rsc_0_15_i_da_d_iff;
  xt_rsc_3_15_i_qa_d <= xt_rsc_3_15_i_qa_d_1;

  xt_rsc_3_16_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_375_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_3_16_i_qa,
      wea => xt_rsc_3_16_wea,
      da => xt_rsc_3_16_i_da,
      adra => xt_rsc_3_16_i_adra,
      adra_d => xt_rsc_3_16_i_adra_d,
      da_d => xt_rsc_3_16_i_da_d,
      qa_d => xt_rsc_3_16_i_qa_d_1,
      wea_d => xt_rsc_3_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_3_16_i_wea_d_iff
    );
  xt_rsc_3_16_i_qa <= xt_rsc_3_16_qa;
  xt_rsc_3_16_da <= xt_rsc_3_16_i_da;
  xt_rsc_3_16_adra <= xt_rsc_3_16_i_adra;
  xt_rsc_3_16_i_adra_d <= xt_rsc_0_0_i_adra_d_iff;
  xt_rsc_3_16_i_da_d <= xt_rsc_0_0_i_da_d_iff;
  xt_rsc_3_16_i_qa_d <= xt_rsc_3_16_i_qa_d_1;

  xt_rsc_3_17_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_376_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_3_17_i_qa,
      wea => xt_rsc_3_17_wea,
      da => xt_rsc_3_17_i_da,
      adra => xt_rsc_3_17_i_adra,
      adra_d => xt_rsc_3_17_i_adra_d,
      da_d => xt_rsc_3_17_i_da_d,
      qa_d => xt_rsc_3_17_i_qa_d_1,
      wea_d => xt_rsc_3_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_3_16_i_wea_d_iff
    );
  xt_rsc_3_17_i_qa <= xt_rsc_3_17_qa;
  xt_rsc_3_17_da <= xt_rsc_3_17_i_da;
  xt_rsc_3_17_adra <= xt_rsc_3_17_i_adra;
  xt_rsc_3_17_i_adra_d <= xt_rsc_0_1_i_adra_d_iff;
  xt_rsc_3_17_i_da_d <= xt_rsc_0_1_i_da_d_iff;
  xt_rsc_3_17_i_qa_d <= xt_rsc_3_17_i_qa_d_1;

  xt_rsc_3_18_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_377_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_3_18_i_qa,
      wea => xt_rsc_3_18_wea,
      da => xt_rsc_3_18_i_da,
      adra => xt_rsc_3_18_i_adra,
      adra_d => xt_rsc_3_18_i_adra_d,
      da_d => xt_rsc_3_18_i_da_d,
      qa_d => xt_rsc_3_18_i_qa_d_1,
      wea_d => xt_rsc_3_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_3_16_i_wea_d_iff
    );
  xt_rsc_3_18_i_qa <= xt_rsc_3_18_qa;
  xt_rsc_3_18_da <= xt_rsc_3_18_i_da;
  xt_rsc_3_18_adra <= xt_rsc_3_18_i_adra;
  xt_rsc_3_18_i_adra_d <= xt_rsc_0_2_i_adra_d_iff;
  xt_rsc_3_18_i_da_d <= xt_rsc_0_2_i_da_d_iff;
  xt_rsc_3_18_i_qa_d <= xt_rsc_3_18_i_qa_d_1;

  xt_rsc_3_19_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_378_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_3_19_i_qa,
      wea => xt_rsc_3_19_wea,
      da => xt_rsc_3_19_i_da,
      adra => xt_rsc_3_19_i_adra,
      adra_d => xt_rsc_3_19_i_adra_d,
      da_d => xt_rsc_3_19_i_da_d,
      qa_d => xt_rsc_3_19_i_qa_d_1,
      wea_d => xt_rsc_3_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_3_16_i_wea_d_iff
    );
  xt_rsc_3_19_i_qa <= xt_rsc_3_19_qa;
  xt_rsc_3_19_da <= xt_rsc_3_19_i_da;
  xt_rsc_3_19_adra <= xt_rsc_3_19_i_adra;
  xt_rsc_3_19_i_adra_d <= xt_rsc_0_3_i_adra_d_iff;
  xt_rsc_3_19_i_da_d <= xt_rsc_0_3_i_da_d_iff;
  xt_rsc_3_19_i_qa_d <= xt_rsc_3_19_i_qa_d_1;

  xt_rsc_3_20_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_379_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_3_20_i_qa,
      wea => xt_rsc_3_20_wea,
      da => xt_rsc_3_20_i_da,
      adra => xt_rsc_3_20_i_adra,
      adra_d => xt_rsc_3_20_i_adra_d,
      da_d => xt_rsc_3_20_i_da_d,
      qa_d => xt_rsc_3_20_i_qa_d_1,
      wea_d => xt_rsc_3_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_3_16_i_wea_d_iff
    );
  xt_rsc_3_20_i_qa <= xt_rsc_3_20_qa;
  xt_rsc_3_20_da <= xt_rsc_3_20_i_da;
  xt_rsc_3_20_adra <= xt_rsc_3_20_i_adra;
  xt_rsc_3_20_i_adra_d <= xt_rsc_0_4_i_adra_d_iff;
  xt_rsc_3_20_i_da_d <= xt_rsc_0_4_i_da_d_iff;
  xt_rsc_3_20_i_qa_d <= xt_rsc_3_20_i_qa_d_1;

  xt_rsc_3_21_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_380_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_3_21_i_qa,
      wea => xt_rsc_3_21_wea,
      da => xt_rsc_3_21_i_da,
      adra => xt_rsc_3_21_i_adra,
      adra_d => xt_rsc_3_21_i_adra_d,
      da_d => xt_rsc_3_21_i_da_d,
      qa_d => xt_rsc_3_21_i_qa_d_1,
      wea_d => xt_rsc_3_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_3_16_i_wea_d_iff
    );
  xt_rsc_3_21_i_qa <= xt_rsc_3_21_qa;
  xt_rsc_3_21_da <= xt_rsc_3_21_i_da;
  xt_rsc_3_21_adra <= xt_rsc_3_21_i_adra;
  xt_rsc_3_21_i_adra_d <= xt_rsc_0_5_i_adra_d_iff;
  xt_rsc_3_21_i_da_d <= xt_rsc_0_5_i_da_d_iff;
  xt_rsc_3_21_i_qa_d <= xt_rsc_3_21_i_qa_d_1;

  xt_rsc_3_22_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_381_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_3_22_i_qa,
      wea => xt_rsc_3_22_wea,
      da => xt_rsc_3_22_i_da,
      adra => xt_rsc_3_22_i_adra,
      adra_d => xt_rsc_3_22_i_adra_d,
      da_d => xt_rsc_3_22_i_da_d,
      qa_d => xt_rsc_3_22_i_qa_d_1,
      wea_d => xt_rsc_3_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_3_16_i_wea_d_iff
    );
  xt_rsc_3_22_i_qa <= xt_rsc_3_22_qa;
  xt_rsc_3_22_da <= xt_rsc_3_22_i_da;
  xt_rsc_3_22_adra <= xt_rsc_3_22_i_adra;
  xt_rsc_3_22_i_adra_d <= xt_rsc_0_6_i_adra_d_iff;
  xt_rsc_3_22_i_da_d <= xt_rsc_0_6_i_da_d_iff;
  xt_rsc_3_22_i_qa_d <= xt_rsc_3_22_i_qa_d_1;

  xt_rsc_3_23_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_382_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_3_23_i_qa,
      wea => xt_rsc_3_23_wea,
      da => xt_rsc_3_23_i_da,
      adra => xt_rsc_3_23_i_adra,
      adra_d => xt_rsc_3_23_i_adra_d,
      da_d => xt_rsc_3_23_i_da_d,
      qa_d => xt_rsc_3_23_i_qa_d_1,
      wea_d => xt_rsc_3_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_3_16_i_wea_d_iff
    );
  xt_rsc_3_23_i_qa <= xt_rsc_3_23_qa;
  xt_rsc_3_23_da <= xt_rsc_3_23_i_da;
  xt_rsc_3_23_adra <= xt_rsc_3_23_i_adra;
  xt_rsc_3_23_i_adra_d <= xt_rsc_0_7_i_adra_d_iff;
  xt_rsc_3_23_i_da_d <= xt_rsc_0_7_i_da_d_iff;
  xt_rsc_3_23_i_qa_d <= xt_rsc_3_23_i_qa_d_1;

  xt_rsc_3_24_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_383_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_3_24_i_qa,
      wea => xt_rsc_3_24_wea,
      da => xt_rsc_3_24_i_da,
      adra => xt_rsc_3_24_i_adra,
      adra_d => xt_rsc_3_24_i_adra_d,
      da_d => xt_rsc_3_24_i_da_d,
      qa_d => xt_rsc_3_24_i_qa_d_1,
      wea_d => xt_rsc_3_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_3_16_i_wea_d_iff
    );
  xt_rsc_3_24_i_qa <= xt_rsc_3_24_qa;
  xt_rsc_3_24_da <= xt_rsc_3_24_i_da;
  xt_rsc_3_24_adra <= xt_rsc_3_24_i_adra;
  xt_rsc_3_24_i_adra_d <= xt_rsc_0_8_i_adra_d_iff;
  xt_rsc_3_24_i_da_d <= xt_rsc_0_8_i_da_d_iff;
  xt_rsc_3_24_i_qa_d <= xt_rsc_3_24_i_qa_d_1;

  xt_rsc_3_25_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_384_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_3_25_i_qa,
      wea => xt_rsc_3_25_wea,
      da => xt_rsc_3_25_i_da,
      adra => xt_rsc_3_25_i_adra,
      adra_d => xt_rsc_3_25_i_adra_d,
      da_d => xt_rsc_3_25_i_da_d,
      qa_d => xt_rsc_3_25_i_qa_d_1,
      wea_d => xt_rsc_3_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_3_16_i_wea_d_iff
    );
  xt_rsc_3_25_i_qa <= xt_rsc_3_25_qa;
  xt_rsc_3_25_da <= xt_rsc_3_25_i_da;
  xt_rsc_3_25_adra <= xt_rsc_3_25_i_adra;
  xt_rsc_3_25_i_adra_d <= xt_rsc_0_9_i_adra_d_iff;
  xt_rsc_3_25_i_da_d <= xt_rsc_0_9_i_da_d_iff;
  xt_rsc_3_25_i_qa_d <= xt_rsc_3_25_i_qa_d_1;

  xt_rsc_3_26_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_385_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_3_26_i_qa,
      wea => xt_rsc_3_26_wea,
      da => xt_rsc_3_26_i_da,
      adra => xt_rsc_3_26_i_adra,
      adra_d => xt_rsc_3_26_i_adra_d,
      da_d => xt_rsc_3_26_i_da_d,
      qa_d => xt_rsc_3_26_i_qa_d_1,
      wea_d => xt_rsc_3_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_3_16_i_wea_d_iff
    );
  xt_rsc_3_26_i_qa <= xt_rsc_3_26_qa;
  xt_rsc_3_26_da <= xt_rsc_3_26_i_da;
  xt_rsc_3_26_adra <= xt_rsc_3_26_i_adra;
  xt_rsc_3_26_i_adra_d <= xt_rsc_0_10_i_adra_d_iff;
  xt_rsc_3_26_i_da_d <= xt_rsc_0_10_i_da_d_iff;
  xt_rsc_3_26_i_qa_d <= xt_rsc_3_26_i_qa_d_1;

  xt_rsc_3_27_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_386_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_3_27_i_qa,
      wea => xt_rsc_3_27_wea,
      da => xt_rsc_3_27_i_da,
      adra => xt_rsc_3_27_i_adra,
      adra_d => xt_rsc_3_27_i_adra_d,
      da_d => xt_rsc_3_27_i_da_d,
      qa_d => xt_rsc_3_27_i_qa_d_1,
      wea_d => xt_rsc_3_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_3_16_i_wea_d_iff
    );
  xt_rsc_3_27_i_qa <= xt_rsc_3_27_qa;
  xt_rsc_3_27_da <= xt_rsc_3_27_i_da;
  xt_rsc_3_27_adra <= xt_rsc_3_27_i_adra;
  xt_rsc_3_27_i_adra_d <= xt_rsc_0_11_i_adra_d_iff;
  xt_rsc_3_27_i_da_d <= xt_rsc_0_11_i_da_d_iff;
  xt_rsc_3_27_i_qa_d <= xt_rsc_3_27_i_qa_d_1;

  xt_rsc_3_28_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_387_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_3_28_i_qa,
      wea => xt_rsc_3_28_wea,
      da => xt_rsc_3_28_i_da,
      adra => xt_rsc_3_28_i_adra,
      adra_d => xt_rsc_3_28_i_adra_d,
      da_d => xt_rsc_3_28_i_da_d,
      qa_d => xt_rsc_3_28_i_qa_d_1,
      wea_d => xt_rsc_3_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_3_16_i_wea_d_iff
    );
  xt_rsc_3_28_i_qa <= xt_rsc_3_28_qa;
  xt_rsc_3_28_da <= xt_rsc_3_28_i_da;
  xt_rsc_3_28_adra <= xt_rsc_3_28_i_adra;
  xt_rsc_3_28_i_adra_d <= xt_rsc_0_12_i_adra_d_iff;
  xt_rsc_3_28_i_da_d <= xt_rsc_0_12_i_da_d_iff;
  xt_rsc_3_28_i_qa_d <= xt_rsc_3_28_i_qa_d_1;

  xt_rsc_3_29_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_388_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_3_29_i_qa,
      wea => xt_rsc_3_29_wea,
      da => xt_rsc_3_29_i_da,
      adra => xt_rsc_3_29_i_adra,
      adra_d => xt_rsc_3_29_i_adra_d,
      da_d => xt_rsc_3_29_i_da_d,
      qa_d => xt_rsc_3_29_i_qa_d_1,
      wea_d => xt_rsc_3_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_3_16_i_wea_d_iff
    );
  xt_rsc_3_29_i_qa <= xt_rsc_3_29_qa;
  xt_rsc_3_29_da <= xt_rsc_3_29_i_da;
  xt_rsc_3_29_adra <= xt_rsc_3_29_i_adra;
  xt_rsc_3_29_i_adra_d <= xt_rsc_0_13_i_adra_d_iff;
  xt_rsc_3_29_i_da_d <= xt_rsc_0_13_i_da_d_iff;
  xt_rsc_3_29_i_qa_d <= xt_rsc_3_29_i_qa_d_1;

  xt_rsc_3_30_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_389_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_3_30_i_qa,
      wea => xt_rsc_3_30_wea,
      da => xt_rsc_3_30_i_da,
      adra => xt_rsc_3_30_i_adra,
      adra_d => xt_rsc_3_30_i_adra_d,
      da_d => xt_rsc_3_30_i_da_d,
      qa_d => xt_rsc_3_30_i_qa_d_1,
      wea_d => xt_rsc_3_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_3_16_i_wea_d_iff
    );
  xt_rsc_3_30_i_qa <= xt_rsc_3_30_qa;
  xt_rsc_3_30_da <= xt_rsc_3_30_i_da;
  xt_rsc_3_30_adra <= xt_rsc_3_30_i_adra;
  xt_rsc_3_30_i_adra_d <= xt_rsc_0_14_i_adra_d_iff;
  xt_rsc_3_30_i_da_d <= xt_rsc_0_14_i_da_d_iff;
  xt_rsc_3_30_i_qa_d <= xt_rsc_3_30_i_qa_d_1;

  xt_rsc_3_31_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_390_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_3_31_i_qa,
      wea => xt_rsc_3_31_wea,
      da => xt_rsc_3_31_i_da,
      adra => xt_rsc_3_31_i_adra,
      adra_d => xt_rsc_3_31_i_adra_d,
      da_d => xt_rsc_3_31_i_da_d,
      qa_d => xt_rsc_3_31_i_qa_d_1,
      wea_d => xt_rsc_3_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_3_16_i_wea_d_iff
    );
  xt_rsc_3_31_i_qa <= xt_rsc_3_31_qa;
  xt_rsc_3_31_da <= xt_rsc_3_31_i_da;
  xt_rsc_3_31_adra <= xt_rsc_3_31_i_adra;
  xt_rsc_3_31_i_adra_d <= xt_rsc_0_15_i_adra_d_iff;
  xt_rsc_3_31_i_da_d <= xt_rsc_0_15_i_da_d_iff;
  xt_rsc_3_31_i_qa_d <= xt_rsc_3_31_i_qa_d_1;

  xt_rsc_4_0_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_391_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_4_0_i_qa,
      wea => xt_rsc_4_0_wea,
      da => xt_rsc_4_0_i_da,
      adra => xt_rsc_4_0_i_adra,
      adra_d => xt_rsc_4_0_i_adra_d,
      da_d => xt_rsc_4_0_i_da_d,
      qa_d => xt_rsc_4_0_i_qa_d_1,
      wea_d => xt_rsc_0_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_0_i_wea_d_iff
    );
  xt_rsc_4_0_i_qa <= xt_rsc_4_0_qa;
  xt_rsc_4_0_da <= xt_rsc_4_0_i_da;
  xt_rsc_4_0_adra <= xt_rsc_4_0_i_adra;
  xt_rsc_4_0_i_adra_d <= xt_rsc_0_8_i_adra_d_iff;
  xt_rsc_4_0_i_da_d <= xt_rsc_4_0_i_da_d_iff;
  xt_rsc_4_0_i_qa_d <= xt_rsc_4_0_i_qa_d_1;

  xt_rsc_4_1_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_392_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_4_1_i_qa,
      wea => xt_rsc_4_1_wea,
      da => xt_rsc_4_1_i_da,
      adra => xt_rsc_4_1_i_adra,
      adra_d => xt_rsc_4_1_i_adra_d,
      da_d => xt_rsc_4_1_i_da_d,
      qa_d => xt_rsc_4_1_i_qa_d_1,
      wea_d => xt_rsc_0_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_0_i_wea_d_iff
    );
  xt_rsc_4_1_i_qa <= xt_rsc_4_1_qa;
  xt_rsc_4_1_da <= xt_rsc_4_1_i_da;
  xt_rsc_4_1_adra <= xt_rsc_4_1_i_adra;
  xt_rsc_4_1_i_adra_d <= xt_rsc_4_1_i_adra_d_iff;
  xt_rsc_4_1_i_da_d <= xt_rsc_4_1_i_da_d_iff;
  xt_rsc_4_1_i_qa_d <= xt_rsc_4_1_i_qa_d_1;

  xt_rsc_4_2_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_393_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_4_2_i_qa,
      wea => xt_rsc_4_2_wea,
      da => xt_rsc_4_2_i_da,
      adra => xt_rsc_4_2_i_adra,
      adra_d => xt_rsc_4_2_i_adra_d,
      da_d => xt_rsc_4_2_i_da_d,
      qa_d => xt_rsc_4_2_i_qa_d_1,
      wea_d => xt_rsc_0_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_0_i_wea_d_iff
    );
  xt_rsc_4_2_i_qa <= xt_rsc_4_2_qa;
  xt_rsc_4_2_da <= xt_rsc_4_2_i_da;
  xt_rsc_4_2_adra <= xt_rsc_4_2_i_adra;
  xt_rsc_4_2_i_adra_d <= xt_rsc_4_2_i_adra_d_iff;
  xt_rsc_4_2_i_da_d <= xt_rsc_4_2_i_da_d_iff;
  xt_rsc_4_2_i_qa_d <= xt_rsc_4_2_i_qa_d_1;

  xt_rsc_4_3_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_394_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_4_3_i_qa,
      wea => xt_rsc_4_3_wea,
      da => xt_rsc_4_3_i_da,
      adra => xt_rsc_4_3_i_adra,
      adra_d => xt_rsc_4_3_i_adra_d,
      da_d => xt_rsc_4_3_i_da_d,
      qa_d => xt_rsc_4_3_i_qa_d_1,
      wea_d => xt_rsc_0_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_0_i_wea_d_iff
    );
  xt_rsc_4_3_i_qa <= xt_rsc_4_3_qa;
  xt_rsc_4_3_da <= xt_rsc_4_3_i_da;
  xt_rsc_4_3_adra <= xt_rsc_4_3_i_adra;
  xt_rsc_4_3_i_adra_d <= xt_rsc_0_12_i_adra_d_iff;
  xt_rsc_4_3_i_da_d <= xt_rsc_4_3_i_da_d_iff;
  xt_rsc_4_3_i_qa_d <= xt_rsc_4_3_i_qa_d_1;

  xt_rsc_4_4_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_395_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_4_4_i_qa,
      wea => xt_rsc_4_4_wea,
      da => xt_rsc_4_4_i_da,
      adra => xt_rsc_4_4_i_adra,
      adra_d => xt_rsc_4_4_i_adra_d,
      da_d => xt_rsc_4_4_i_da_d,
      qa_d => xt_rsc_4_4_i_qa_d_1,
      wea_d => xt_rsc_0_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_0_i_wea_d_iff
    );
  xt_rsc_4_4_i_qa <= xt_rsc_4_4_qa;
  xt_rsc_4_4_da <= xt_rsc_4_4_i_da;
  xt_rsc_4_4_adra <= xt_rsc_4_4_i_adra;
  xt_rsc_4_4_i_adra_d <= xt_rsc_0_13_i_adra_d_iff;
  xt_rsc_4_4_i_da_d <= xt_rsc_4_4_i_da_d_iff;
  xt_rsc_4_4_i_qa_d <= xt_rsc_4_4_i_qa_d_1;

  xt_rsc_4_5_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_396_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_4_5_i_qa,
      wea => xt_rsc_4_5_wea,
      da => xt_rsc_4_5_i_da,
      adra => xt_rsc_4_5_i_adra,
      adra_d => xt_rsc_4_5_i_adra_d,
      da_d => xt_rsc_4_5_i_da_d,
      qa_d => xt_rsc_4_5_i_qa_d_1,
      wea_d => xt_rsc_0_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_0_i_wea_d_iff
    );
  xt_rsc_4_5_i_qa <= xt_rsc_4_5_qa;
  xt_rsc_4_5_da <= xt_rsc_4_5_i_da;
  xt_rsc_4_5_adra <= xt_rsc_4_5_i_adra;
  xt_rsc_4_5_i_adra_d <= xt_rsc_0_14_i_adra_d_iff;
  xt_rsc_4_5_i_da_d <= xt_rsc_4_5_i_da_d_iff;
  xt_rsc_4_5_i_qa_d <= xt_rsc_4_5_i_qa_d_1;

  xt_rsc_4_6_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_397_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_4_6_i_qa,
      wea => xt_rsc_4_6_wea,
      da => xt_rsc_4_6_i_da,
      adra => xt_rsc_4_6_i_adra,
      adra_d => xt_rsc_4_6_i_adra_d,
      da_d => xt_rsc_4_6_i_da_d,
      qa_d => xt_rsc_4_6_i_qa_d_1,
      wea_d => xt_rsc_0_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_0_i_wea_d_iff
    );
  xt_rsc_4_6_i_qa <= xt_rsc_4_6_qa;
  xt_rsc_4_6_da <= xt_rsc_4_6_i_da;
  xt_rsc_4_6_adra <= xt_rsc_4_6_i_adra;
  xt_rsc_4_6_i_adra_d <= xt_rsc_0_15_i_adra_d_iff;
  xt_rsc_4_6_i_da_d <= xt_rsc_4_6_i_da_d_iff;
  xt_rsc_4_6_i_qa_d <= xt_rsc_4_6_i_qa_d_1;

  xt_rsc_4_7_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_398_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_4_7_i_qa,
      wea => xt_rsc_4_7_wea,
      da => xt_rsc_4_7_i_da,
      adra => xt_rsc_4_7_i_adra,
      adra_d => xt_rsc_4_7_i_adra_d,
      da_d => xt_rsc_4_7_i_da_d,
      qa_d => xt_rsc_4_7_i_qa_d_1,
      wea_d => xt_rsc_0_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_0_i_wea_d_iff
    );
  xt_rsc_4_7_i_qa <= xt_rsc_4_7_qa;
  xt_rsc_4_7_da <= xt_rsc_4_7_i_da;
  xt_rsc_4_7_adra <= xt_rsc_4_7_i_adra;
  xt_rsc_4_7_i_adra_d <= xt_rsc_0_0_i_adra_d_iff;
  xt_rsc_4_7_i_da_d <= xt_rsc_4_7_i_da_d_iff;
  xt_rsc_4_7_i_qa_d <= xt_rsc_4_7_i_qa_d_1;

  xt_rsc_4_8_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_399_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_4_8_i_qa,
      wea => xt_rsc_4_8_wea,
      da => xt_rsc_4_8_i_da,
      adra => xt_rsc_4_8_i_adra,
      adra_d => xt_rsc_4_8_i_adra_d,
      da_d => xt_rsc_4_8_i_da_d,
      qa_d => xt_rsc_4_8_i_qa_d_1,
      wea_d => xt_rsc_0_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_0_i_wea_d_iff
    );
  xt_rsc_4_8_i_qa <= xt_rsc_4_8_qa;
  xt_rsc_4_8_da <= xt_rsc_4_8_i_da;
  xt_rsc_4_8_adra <= xt_rsc_4_8_i_adra;
  xt_rsc_4_8_i_adra_d <= xt_rsc_0_1_i_adra_d_iff;
  xt_rsc_4_8_i_da_d <= xt_rsc_4_8_i_da_d_iff;
  xt_rsc_4_8_i_qa_d <= xt_rsc_4_8_i_qa_d_1;

  xt_rsc_4_9_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_400_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_4_9_i_qa,
      wea => xt_rsc_4_9_wea,
      da => xt_rsc_4_9_i_da,
      adra => xt_rsc_4_9_i_adra,
      adra_d => xt_rsc_4_9_i_adra_d,
      da_d => xt_rsc_4_9_i_da_d,
      qa_d => xt_rsc_4_9_i_qa_d_1,
      wea_d => xt_rsc_0_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_0_i_wea_d_iff
    );
  xt_rsc_4_9_i_qa <= xt_rsc_4_9_qa;
  xt_rsc_4_9_da <= xt_rsc_4_9_i_da;
  xt_rsc_4_9_adra <= xt_rsc_4_9_i_adra;
  xt_rsc_4_9_i_adra_d <= xt_rsc_4_9_i_adra_d_iff;
  xt_rsc_4_9_i_da_d <= xt_rsc_4_9_i_da_d_iff;
  xt_rsc_4_9_i_qa_d <= xt_rsc_4_9_i_qa_d_1;

  xt_rsc_4_10_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_401_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_4_10_i_qa,
      wea => xt_rsc_4_10_wea,
      da => xt_rsc_4_10_i_da,
      adra => xt_rsc_4_10_i_adra,
      adra_d => xt_rsc_4_10_i_adra_d,
      da_d => xt_rsc_4_10_i_da_d,
      qa_d => xt_rsc_4_10_i_qa_d_1,
      wea_d => xt_rsc_0_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_0_i_wea_d_iff
    );
  xt_rsc_4_10_i_qa <= xt_rsc_4_10_qa;
  xt_rsc_4_10_da <= xt_rsc_4_10_i_da;
  xt_rsc_4_10_adra <= xt_rsc_4_10_i_adra;
  xt_rsc_4_10_i_adra_d <= xt_rsc_4_10_i_adra_d_iff;
  xt_rsc_4_10_i_da_d <= xt_rsc_4_10_i_da_d_iff;
  xt_rsc_4_10_i_qa_d <= xt_rsc_4_10_i_qa_d_1;

  xt_rsc_4_11_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_402_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_4_11_i_qa,
      wea => xt_rsc_4_11_wea,
      da => xt_rsc_4_11_i_da,
      adra => xt_rsc_4_11_i_adra,
      adra_d => xt_rsc_4_11_i_adra_d,
      da_d => xt_rsc_4_11_i_da_d,
      qa_d => xt_rsc_4_11_i_qa_d_1,
      wea_d => xt_rsc_0_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_0_i_wea_d_iff
    );
  xt_rsc_4_11_i_qa <= xt_rsc_4_11_qa;
  xt_rsc_4_11_da <= xt_rsc_4_11_i_da;
  xt_rsc_4_11_adra <= xt_rsc_4_11_i_adra;
  xt_rsc_4_11_i_adra_d <= xt_rsc_0_3_i_adra_d_iff;
  xt_rsc_4_11_i_da_d <= xt_rsc_4_11_i_da_d_iff;
  xt_rsc_4_11_i_qa_d <= xt_rsc_4_11_i_qa_d_1;

  xt_rsc_4_12_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_403_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_4_12_i_qa,
      wea => xt_rsc_4_12_wea,
      da => xt_rsc_4_12_i_da,
      adra => xt_rsc_4_12_i_adra,
      adra_d => xt_rsc_4_12_i_adra_d,
      da_d => xt_rsc_4_12_i_da_d,
      qa_d => xt_rsc_4_12_i_qa_d_1,
      wea_d => xt_rsc_0_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_0_i_wea_d_iff
    );
  xt_rsc_4_12_i_qa <= xt_rsc_4_12_qa;
  xt_rsc_4_12_da <= xt_rsc_4_12_i_da;
  xt_rsc_4_12_adra <= xt_rsc_4_12_i_adra;
  xt_rsc_4_12_i_adra_d <= xt_rsc_0_4_i_adra_d_iff;
  xt_rsc_4_12_i_da_d <= xt_rsc_4_12_i_da_d_iff;
  xt_rsc_4_12_i_qa_d <= xt_rsc_4_12_i_qa_d_1;

  xt_rsc_4_13_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_404_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_4_13_i_qa,
      wea => xt_rsc_4_13_wea,
      da => xt_rsc_4_13_i_da,
      adra => xt_rsc_4_13_i_adra,
      adra_d => xt_rsc_4_13_i_adra_d,
      da_d => xt_rsc_4_13_i_da_d,
      qa_d => xt_rsc_4_13_i_qa_d_1,
      wea_d => xt_rsc_0_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_0_i_wea_d_iff
    );
  xt_rsc_4_13_i_qa <= xt_rsc_4_13_qa;
  xt_rsc_4_13_da <= xt_rsc_4_13_i_da;
  xt_rsc_4_13_adra <= xt_rsc_4_13_i_adra;
  xt_rsc_4_13_i_adra_d <= xt_rsc_0_5_i_adra_d_iff;
  xt_rsc_4_13_i_da_d <= xt_rsc_4_13_i_da_d_iff;
  xt_rsc_4_13_i_qa_d <= xt_rsc_4_13_i_qa_d_1;

  xt_rsc_4_14_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_405_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_4_14_i_qa,
      wea => xt_rsc_4_14_wea,
      da => xt_rsc_4_14_i_da,
      adra => xt_rsc_4_14_i_adra,
      adra_d => xt_rsc_4_14_i_adra_d,
      da_d => xt_rsc_4_14_i_da_d,
      qa_d => xt_rsc_4_14_i_qa_d_1,
      wea_d => xt_rsc_0_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_0_i_wea_d_iff
    );
  xt_rsc_4_14_i_qa <= xt_rsc_4_14_qa;
  xt_rsc_4_14_da <= xt_rsc_4_14_i_da;
  xt_rsc_4_14_adra <= xt_rsc_4_14_i_adra;
  xt_rsc_4_14_i_adra_d <= xt_rsc_0_6_i_adra_d_iff;
  xt_rsc_4_14_i_da_d <= xt_rsc_4_14_i_da_d_iff;
  xt_rsc_4_14_i_qa_d <= xt_rsc_4_14_i_qa_d_1;

  xt_rsc_4_15_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_406_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_4_15_i_qa,
      wea => xt_rsc_4_15_wea,
      da => xt_rsc_4_15_i_da,
      adra => xt_rsc_4_15_i_adra,
      adra_d => xt_rsc_4_15_i_adra_d,
      da_d => xt_rsc_4_15_i_da_d,
      qa_d => xt_rsc_4_15_i_qa_d_1,
      wea_d => xt_rsc_0_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_0_i_wea_d_iff
    );
  xt_rsc_4_15_i_qa <= xt_rsc_4_15_qa;
  xt_rsc_4_15_da <= xt_rsc_4_15_i_da;
  xt_rsc_4_15_adra <= xt_rsc_4_15_i_adra;
  xt_rsc_4_15_i_adra_d <= xt_rsc_0_7_i_adra_d_iff;
  xt_rsc_4_15_i_da_d <= xt_rsc_4_15_i_da_d_iff;
  xt_rsc_4_15_i_qa_d <= xt_rsc_4_15_i_qa_d_1;

  xt_rsc_4_16_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_407_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_4_16_i_qa,
      wea => xt_rsc_4_16_wea,
      da => xt_rsc_4_16_i_da,
      adra => xt_rsc_4_16_i_adra,
      adra_d => xt_rsc_4_16_i_adra_d,
      da_d => xt_rsc_4_16_i_da_d,
      qa_d => xt_rsc_4_16_i_qa_d_1,
      wea_d => xt_rsc_0_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_16_i_wea_d_iff
    );
  xt_rsc_4_16_i_qa <= xt_rsc_4_16_qa;
  xt_rsc_4_16_da <= xt_rsc_4_16_i_da;
  xt_rsc_4_16_adra <= xt_rsc_4_16_i_adra;
  xt_rsc_4_16_i_adra_d <= xt_rsc_0_8_i_adra_d_iff;
  xt_rsc_4_16_i_da_d <= xt_rsc_4_0_i_da_d_iff;
  xt_rsc_4_16_i_qa_d <= xt_rsc_4_16_i_qa_d_1;

  xt_rsc_4_17_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_408_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_4_17_i_qa,
      wea => xt_rsc_4_17_wea,
      da => xt_rsc_4_17_i_da,
      adra => xt_rsc_4_17_i_adra,
      adra_d => xt_rsc_4_17_i_adra_d,
      da_d => xt_rsc_4_17_i_da_d,
      qa_d => xt_rsc_4_17_i_qa_d_1,
      wea_d => xt_rsc_0_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_16_i_wea_d_iff
    );
  xt_rsc_4_17_i_qa <= xt_rsc_4_17_qa;
  xt_rsc_4_17_da <= xt_rsc_4_17_i_da;
  xt_rsc_4_17_adra <= xt_rsc_4_17_i_adra;
  xt_rsc_4_17_i_adra_d <= xt_rsc_4_1_i_adra_d_iff;
  xt_rsc_4_17_i_da_d <= xt_rsc_4_1_i_da_d_iff;
  xt_rsc_4_17_i_qa_d <= xt_rsc_4_17_i_qa_d_1;

  xt_rsc_4_18_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_409_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_4_18_i_qa,
      wea => xt_rsc_4_18_wea,
      da => xt_rsc_4_18_i_da,
      adra => xt_rsc_4_18_i_adra,
      adra_d => xt_rsc_4_18_i_adra_d,
      da_d => xt_rsc_4_18_i_da_d,
      qa_d => xt_rsc_4_18_i_qa_d_1,
      wea_d => xt_rsc_0_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_16_i_wea_d_iff
    );
  xt_rsc_4_18_i_qa <= xt_rsc_4_18_qa;
  xt_rsc_4_18_da <= xt_rsc_4_18_i_da;
  xt_rsc_4_18_adra <= xt_rsc_4_18_i_adra;
  xt_rsc_4_18_i_adra_d <= xt_rsc_4_2_i_adra_d_iff;
  xt_rsc_4_18_i_da_d <= xt_rsc_4_2_i_da_d_iff;
  xt_rsc_4_18_i_qa_d <= xt_rsc_4_18_i_qa_d_1;

  xt_rsc_4_19_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_410_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_4_19_i_qa,
      wea => xt_rsc_4_19_wea,
      da => xt_rsc_4_19_i_da,
      adra => xt_rsc_4_19_i_adra,
      adra_d => xt_rsc_4_19_i_adra_d,
      da_d => xt_rsc_4_19_i_da_d,
      qa_d => xt_rsc_4_19_i_qa_d_1,
      wea_d => xt_rsc_0_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_16_i_wea_d_iff
    );
  xt_rsc_4_19_i_qa <= xt_rsc_4_19_qa;
  xt_rsc_4_19_da <= xt_rsc_4_19_i_da;
  xt_rsc_4_19_adra <= xt_rsc_4_19_i_adra;
  xt_rsc_4_19_i_adra_d <= xt_rsc_0_12_i_adra_d_iff;
  xt_rsc_4_19_i_da_d <= xt_rsc_4_3_i_da_d_iff;
  xt_rsc_4_19_i_qa_d <= xt_rsc_4_19_i_qa_d_1;

  xt_rsc_4_20_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_411_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_4_20_i_qa,
      wea => xt_rsc_4_20_wea,
      da => xt_rsc_4_20_i_da,
      adra => xt_rsc_4_20_i_adra,
      adra_d => xt_rsc_4_20_i_adra_d,
      da_d => xt_rsc_4_20_i_da_d,
      qa_d => xt_rsc_4_20_i_qa_d_1,
      wea_d => xt_rsc_0_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_16_i_wea_d_iff
    );
  xt_rsc_4_20_i_qa <= xt_rsc_4_20_qa;
  xt_rsc_4_20_da <= xt_rsc_4_20_i_da;
  xt_rsc_4_20_adra <= xt_rsc_4_20_i_adra;
  xt_rsc_4_20_i_adra_d <= xt_rsc_0_13_i_adra_d_iff;
  xt_rsc_4_20_i_da_d <= xt_rsc_4_4_i_da_d_iff;
  xt_rsc_4_20_i_qa_d <= xt_rsc_4_20_i_qa_d_1;

  xt_rsc_4_21_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_412_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_4_21_i_qa,
      wea => xt_rsc_4_21_wea,
      da => xt_rsc_4_21_i_da,
      adra => xt_rsc_4_21_i_adra,
      adra_d => xt_rsc_4_21_i_adra_d,
      da_d => xt_rsc_4_21_i_da_d,
      qa_d => xt_rsc_4_21_i_qa_d_1,
      wea_d => xt_rsc_0_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_16_i_wea_d_iff
    );
  xt_rsc_4_21_i_qa <= xt_rsc_4_21_qa;
  xt_rsc_4_21_da <= xt_rsc_4_21_i_da;
  xt_rsc_4_21_adra <= xt_rsc_4_21_i_adra;
  xt_rsc_4_21_i_adra_d <= xt_rsc_0_14_i_adra_d_iff;
  xt_rsc_4_21_i_da_d <= xt_rsc_4_5_i_da_d_iff;
  xt_rsc_4_21_i_qa_d <= xt_rsc_4_21_i_qa_d_1;

  xt_rsc_4_22_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_413_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_4_22_i_qa,
      wea => xt_rsc_4_22_wea,
      da => xt_rsc_4_22_i_da,
      adra => xt_rsc_4_22_i_adra,
      adra_d => xt_rsc_4_22_i_adra_d,
      da_d => xt_rsc_4_22_i_da_d,
      qa_d => xt_rsc_4_22_i_qa_d_1,
      wea_d => xt_rsc_0_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_16_i_wea_d_iff
    );
  xt_rsc_4_22_i_qa <= xt_rsc_4_22_qa;
  xt_rsc_4_22_da <= xt_rsc_4_22_i_da;
  xt_rsc_4_22_adra <= xt_rsc_4_22_i_adra;
  xt_rsc_4_22_i_adra_d <= xt_rsc_0_15_i_adra_d_iff;
  xt_rsc_4_22_i_da_d <= xt_rsc_4_6_i_da_d_iff;
  xt_rsc_4_22_i_qa_d <= xt_rsc_4_22_i_qa_d_1;

  xt_rsc_4_23_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_414_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_4_23_i_qa,
      wea => xt_rsc_4_23_wea,
      da => xt_rsc_4_23_i_da,
      adra => xt_rsc_4_23_i_adra,
      adra_d => xt_rsc_4_23_i_adra_d,
      da_d => xt_rsc_4_23_i_da_d,
      qa_d => xt_rsc_4_23_i_qa_d_1,
      wea_d => xt_rsc_0_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_16_i_wea_d_iff
    );
  xt_rsc_4_23_i_qa <= xt_rsc_4_23_qa;
  xt_rsc_4_23_da <= xt_rsc_4_23_i_da;
  xt_rsc_4_23_adra <= xt_rsc_4_23_i_adra;
  xt_rsc_4_23_i_adra_d <= xt_rsc_0_0_i_adra_d_iff;
  xt_rsc_4_23_i_da_d <= xt_rsc_4_7_i_da_d_iff;
  xt_rsc_4_23_i_qa_d <= xt_rsc_4_23_i_qa_d_1;

  xt_rsc_4_24_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_415_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_4_24_i_qa,
      wea => xt_rsc_4_24_wea,
      da => xt_rsc_4_24_i_da,
      adra => xt_rsc_4_24_i_adra,
      adra_d => xt_rsc_4_24_i_adra_d,
      da_d => xt_rsc_4_24_i_da_d,
      qa_d => xt_rsc_4_24_i_qa_d_1,
      wea_d => xt_rsc_0_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_16_i_wea_d_iff
    );
  xt_rsc_4_24_i_qa <= xt_rsc_4_24_qa;
  xt_rsc_4_24_da <= xt_rsc_4_24_i_da;
  xt_rsc_4_24_adra <= xt_rsc_4_24_i_adra;
  xt_rsc_4_24_i_adra_d <= xt_rsc_0_1_i_adra_d_iff;
  xt_rsc_4_24_i_da_d <= xt_rsc_4_8_i_da_d_iff;
  xt_rsc_4_24_i_qa_d <= xt_rsc_4_24_i_qa_d_1;

  xt_rsc_4_25_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_416_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_4_25_i_qa,
      wea => xt_rsc_4_25_wea,
      da => xt_rsc_4_25_i_da,
      adra => xt_rsc_4_25_i_adra,
      adra_d => xt_rsc_4_25_i_adra_d,
      da_d => xt_rsc_4_25_i_da_d,
      qa_d => xt_rsc_4_25_i_qa_d_1,
      wea_d => xt_rsc_0_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_16_i_wea_d_iff
    );
  xt_rsc_4_25_i_qa <= xt_rsc_4_25_qa;
  xt_rsc_4_25_da <= xt_rsc_4_25_i_da;
  xt_rsc_4_25_adra <= xt_rsc_4_25_i_adra;
  xt_rsc_4_25_i_adra_d <= xt_rsc_4_9_i_adra_d_iff;
  xt_rsc_4_25_i_da_d <= xt_rsc_4_9_i_da_d_iff;
  xt_rsc_4_25_i_qa_d <= xt_rsc_4_25_i_qa_d_1;

  xt_rsc_4_26_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_417_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_4_26_i_qa,
      wea => xt_rsc_4_26_wea,
      da => xt_rsc_4_26_i_da,
      adra => xt_rsc_4_26_i_adra,
      adra_d => xt_rsc_4_26_i_adra_d,
      da_d => xt_rsc_4_26_i_da_d,
      qa_d => xt_rsc_4_26_i_qa_d_1,
      wea_d => xt_rsc_0_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_16_i_wea_d_iff
    );
  xt_rsc_4_26_i_qa <= xt_rsc_4_26_qa;
  xt_rsc_4_26_da <= xt_rsc_4_26_i_da;
  xt_rsc_4_26_adra <= xt_rsc_4_26_i_adra;
  xt_rsc_4_26_i_adra_d <= xt_rsc_4_10_i_adra_d_iff;
  xt_rsc_4_26_i_da_d <= xt_rsc_4_10_i_da_d_iff;
  xt_rsc_4_26_i_qa_d <= xt_rsc_4_26_i_qa_d_1;

  xt_rsc_4_27_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_418_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_4_27_i_qa,
      wea => xt_rsc_4_27_wea,
      da => xt_rsc_4_27_i_da,
      adra => xt_rsc_4_27_i_adra,
      adra_d => xt_rsc_4_27_i_adra_d,
      da_d => xt_rsc_4_27_i_da_d,
      qa_d => xt_rsc_4_27_i_qa_d_1,
      wea_d => xt_rsc_0_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_16_i_wea_d_iff
    );
  xt_rsc_4_27_i_qa <= xt_rsc_4_27_qa;
  xt_rsc_4_27_da <= xt_rsc_4_27_i_da;
  xt_rsc_4_27_adra <= xt_rsc_4_27_i_adra;
  xt_rsc_4_27_i_adra_d <= xt_rsc_0_3_i_adra_d_iff;
  xt_rsc_4_27_i_da_d <= xt_rsc_4_11_i_da_d_iff;
  xt_rsc_4_27_i_qa_d <= xt_rsc_4_27_i_qa_d_1;

  xt_rsc_4_28_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_419_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_4_28_i_qa,
      wea => xt_rsc_4_28_wea,
      da => xt_rsc_4_28_i_da,
      adra => xt_rsc_4_28_i_adra,
      adra_d => xt_rsc_4_28_i_adra_d,
      da_d => xt_rsc_4_28_i_da_d,
      qa_d => xt_rsc_4_28_i_qa_d_1,
      wea_d => xt_rsc_0_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_16_i_wea_d_iff
    );
  xt_rsc_4_28_i_qa <= xt_rsc_4_28_qa;
  xt_rsc_4_28_da <= xt_rsc_4_28_i_da;
  xt_rsc_4_28_adra <= xt_rsc_4_28_i_adra;
  xt_rsc_4_28_i_adra_d <= xt_rsc_0_4_i_adra_d_iff;
  xt_rsc_4_28_i_da_d <= xt_rsc_4_12_i_da_d_iff;
  xt_rsc_4_28_i_qa_d <= xt_rsc_4_28_i_qa_d_1;

  xt_rsc_4_29_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_420_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_4_29_i_qa,
      wea => xt_rsc_4_29_wea,
      da => xt_rsc_4_29_i_da,
      adra => xt_rsc_4_29_i_adra,
      adra_d => xt_rsc_4_29_i_adra_d,
      da_d => xt_rsc_4_29_i_da_d,
      qa_d => xt_rsc_4_29_i_qa_d_1,
      wea_d => xt_rsc_0_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_16_i_wea_d_iff
    );
  xt_rsc_4_29_i_qa <= xt_rsc_4_29_qa;
  xt_rsc_4_29_da <= xt_rsc_4_29_i_da;
  xt_rsc_4_29_adra <= xt_rsc_4_29_i_adra;
  xt_rsc_4_29_i_adra_d <= xt_rsc_0_5_i_adra_d_iff;
  xt_rsc_4_29_i_da_d <= xt_rsc_4_13_i_da_d_iff;
  xt_rsc_4_29_i_qa_d <= xt_rsc_4_29_i_qa_d_1;

  xt_rsc_4_30_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_421_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_4_30_i_qa,
      wea => xt_rsc_4_30_wea,
      da => xt_rsc_4_30_i_da,
      adra => xt_rsc_4_30_i_adra,
      adra_d => xt_rsc_4_30_i_adra_d,
      da_d => xt_rsc_4_30_i_da_d,
      qa_d => xt_rsc_4_30_i_qa_d_1,
      wea_d => xt_rsc_0_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_16_i_wea_d_iff
    );
  xt_rsc_4_30_i_qa <= xt_rsc_4_30_qa;
  xt_rsc_4_30_da <= xt_rsc_4_30_i_da;
  xt_rsc_4_30_adra <= xt_rsc_4_30_i_adra;
  xt_rsc_4_30_i_adra_d <= xt_rsc_0_6_i_adra_d_iff;
  xt_rsc_4_30_i_da_d <= xt_rsc_4_14_i_da_d_iff;
  xt_rsc_4_30_i_qa_d <= xt_rsc_4_30_i_qa_d_1;

  xt_rsc_4_31_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_422_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_4_31_i_qa,
      wea => xt_rsc_4_31_wea,
      da => xt_rsc_4_31_i_da,
      adra => xt_rsc_4_31_i_adra,
      adra_d => xt_rsc_4_31_i_adra_d,
      da_d => xt_rsc_4_31_i_da_d,
      qa_d => xt_rsc_4_31_i_qa_d_1,
      wea_d => xt_rsc_0_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_16_i_wea_d_iff
    );
  xt_rsc_4_31_i_qa <= xt_rsc_4_31_qa;
  xt_rsc_4_31_da <= xt_rsc_4_31_i_da;
  xt_rsc_4_31_adra <= xt_rsc_4_31_i_adra;
  xt_rsc_4_31_i_adra_d <= xt_rsc_0_7_i_adra_d_iff;
  xt_rsc_4_31_i_da_d <= xt_rsc_4_15_i_da_d_iff;
  xt_rsc_4_31_i_qa_d <= xt_rsc_4_31_i_qa_d_1;

  xt_rsc_5_0_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_423_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_5_0_i_qa,
      wea => xt_rsc_5_0_wea,
      da => xt_rsc_5_0_i_da,
      adra => xt_rsc_5_0_i_adra,
      adra_d => xt_rsc_5_0_i_adra_d,
      da_d => xt_rsc_5_0_i_da_d,
      qa_d => xt_rsc_5_0_i_qa_d_1,
      wea_d => xt_rsc_1_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_0_i_wea_d_iff
    );
  xt_rsc_5_0_i_qa <= xt_rsc_5_0_qa;
  xt_rsc_5_0_da <= xt_rsc_5_0_i_da;
  xt_rsc_5_0_adra <= xt_rsc_5_0_i_adra;
  xt_rsc_5_0_i_adra_d <= xt_rsc_0_8_i_adra_d_iff;
  xt_rsc_5_0_i_da_d <= xt_rsc_4_0_i_da_d_iff;
  xt_rsc_5_0_i_qa_d <= xt_rsc_5_0_i_qa_d_1;

  xt_rsc_5_1_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_424_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_5_1_i_qa,
      wea => xt_rsc_5_1_wea,
      da => xt_rsc_5_1_i_da,
      adra => xt_rsc_5_1_i_adra,
      adra_d => xt_rsc_5_1_i_adra_d,
      da_d => xt_rsc_5_1_i_da_d,
      qa_d => xt_rsc_5_1_i_qa_d_1,
      wea_d => xt_rsc_1_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_0_i_wea_d_iff
    );
  xt_rsc_5_1_i_qa <= xt_rsc_5_1_qa;
  xt_rsc_5_1_da <= xt_rsc_5_1_i_da;
  xt_rsc_5_1_adra <= xt_rsc_5_1_i_adra;
  xt_rsc_5_1_i_adra_d <= xt_rsc_4_1_i_adra_d_iff;
  xt_rsc_5_1_i_da_d <= xt_rsc_4_1_i_da_d_iff;
  xt_rsc_5_1_i_qa_d <= xt_rsc_5_1_i_qa_d_1;

  xt_rsc_5_2_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_425_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_5_2_i_qa,
      wea => xt_rsc_5_2_wea,
      da => xt_rsc_5_2_i_da,
      adra => xt_rsc_5_2_i_adra,
      adra_d => xt_rsc_5_2_i_adra_d,
      da_d => xt_rsc_5_2_i_da_d,
      qa_d => xt_rsc_5_2_i_qa_d_1,
      wea_d => xt_rsc_1_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_0_i_wea_d_iff
    );
  xt_rsc_5_2_i_qa <= xt_rsc_5_2_qa;
  xt_rsc_5_2_da <= xt_rsc_5_2_i_da;
  xt_rsc_5_2_adra <= xt_rsc_5_2_i_adra;
  xt_rsc_5_2_i_adra_d <= xt_rsc_4_2_i_adra_d_iff;
  xt_rsc_5_2_i_da_d <= xt_rsc_4_2_i_da_d_iff;
  xt_rsc_5_2_i_qa_d <= xt_rsc_5_2_i_qa_d_1;

  xt_rsc_5_3_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_426_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_5_3_i_qa,
      wea => xt_rsc_5_3_wea,
      da => xt_rsc_5_3_i_da,
      adra => xt_rsc_5_3_i_adra,
      adra_d => xt_rsc_5_3_i_adra_d,
      da_d => xt_rsc_5_3_i_da_d,
      qa_d => xt_rsc_5_3_i_qa_d_1,
      wea_d => xt_rsc_1_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_0_i_wea_d_iff
    );
  xt_rsc_5_3_i_qa <= xt_rsc_5_3_qa;
  xt_rsc_5_3_da <= xt_rsc_5_3_i_da;
  xt_rsc_5_3_adra <= xt_rsc_5_3_i_adra;
  xt_rsc_5_3_i_adra_d <= xt_rsc_0_12_i_adra_d_iff;
  xt_rsc_5_3_i_da_d <= xt_rsc_4_3_i_da_d_iff;
  xt_rsc_5_3_i_qa_d <= xt_rsc_5_3_i_qa_d_1;

  xt_rsc_5_4_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_427_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_5_4_i_qa,
      wea => xt_rsc_5_4_wea,
      da => xt_rsc_5_4_i_da,
      adra => xt_rsc_5_4_i_adra,
      adra_d => xt_rsc_5_4_i_adra_d,
      da_d => xt_rsc_5_4_i_da_d,
      qa_d => xt_rsc_5_4_i_qa_d_1,
      wea_d => xt_rsc_1_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_0_i_wea_d_iff
    );
  xt_rsc_5_4_i_qa <= xt_rsc_5_4_qa;
  xt_rsc_5_4_da <= xt_rsc_5_4_i_da;
  xt_rsc_5_4_adra <= xt_rsc_5_4_i_adra;
  xt_rsc_5_4_i_adra_d <= xt_rsc_0_13_i_adra_d_iff;
  xt_rsc_5_4_i_da_d <= xt_rsc_4_4_i_da_d_iff;
  xt_rsc_5_4_i_qa_d <= xt_rsc_5_4_i_qa_d_1;

  xt_rsc_5_5_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_428_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_5_5_i_qa,
      wea => xt_rsc_5_5_wea,
      da => xt_rsc_5_5_i_da,
      adra => xt_rsc_5_5_i_adra,
      adra_d => xt_rsc_5_5_i_adra_d,
      da_d => xt_rsc_5_5_i_da_d,
      qa_d => xt_rsc_5_5_i_qa_d_1,
      wea_d => xt_rsc_1_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_0_i_wea_d_iff
    );
  xt_rsc_5_5_i_qa <= xt_rsc_5_5_qa;
  xt_rsc_5_5_da <= xt_rsc_5_5_i_da;
  xt_rsc_5_5_adra <= xt_rsc_5_5_i_adra;
  xt_rsc_5_5_i_adra_d <= xt_rsc_0_14_i_adra_d_iff;
  xt_rsc_5_5_i_da_d <= xt_rsc_4_5_i_da_d_iff;
  xt_rsc_5_5_i_qa_d <= xt_rsc_5_5_i_qa_d_1;

  xt_rsc_5_6_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_429_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_5_6_i_qa,
      wea => xt_rsc_5_6_wea,
      da => xt_rsc_5_6_i_da,
      adra => xt_rsc_5_6_i_adra,
      adra_d => xt_rsc_5_6_i_adra_d,
      da_d => xt_rsc_5_6_i_da_d,
      qa_d => xt_rsc_5_6_i_qa_d_1,
      wea_d => xt_rsc_1_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_0_i_wea_d_iff
    );
  xt_rsc_5_6_i_qa <= xt_rsc_5_6_qa;
  xt_rsc_5_6_da <= xt_rsc_5_6_i_da;
  xt_rsc_5_6_adra <= xt_rsc_5_6_i_adra;
  xt_rsc_5_6_i_adra_d <= xt_rsc_0_15_i_adra_d_iff;
  xt_rsc_5_6_i_da_d <= xt_rsc_4_6_i_da_d_iff;
  xt_rsc_5_6_i_qa_d <= xt_rsc_5_6_i_qa_d_1;

  xt_rsc_5_7_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_430_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_5_7_i_qa,
      wea => xt_rsc_5_7_wea,
      da => xt_rsc_5_7_i_da,
      adra => xt_rsc_5_7_i_adra,
      adra_d => xt_rsc_5_7_i_adra_d,
      da_d => xt_rsc_5_7_i_da_d,
      qa_d => xt_rsc_5_7_i_qa_d_1,
      wea_d => xt_rsc_1_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_0_i_wea_d_iff
    );
  xt_rsc_5_7_i_qa <= xt_rsc_5_7_qa;
  xt_rsc_5_7_da <= xt_rsc_5_7_i_da;
  xt_rsc_5_7_adra <= xt_rsc_5_7_i_adra;
  xt_rsc_5_7_i_adra_d <= xt_rsc_0_0_i_adra_d_iff;
  xt_rsc_5_7_i_da_d <= xt_rsc_4_7_i_da_d_iff;
  xt_rsc_5_7_i_qa_d <= xt_rsc_5_7_i_qa_d_1;

  xt_rsc_5_8_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_431_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_5_8_i_qa,
      wea => xt_rsc_5_8_wea,
      da => xt_rsc_5_8_i_da,
      adra => xt_rsc_5_8_i_adra,
      adra_d => xt_rsc_5_8_i_adra_d,
      da_d => xt_rsc_5_8_i_da_d,
      qa_d => xt_rsc_5_8_i_qa_d_1,
      wea_d => xt_rsc_1_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_0_i_wea_d_iff
    );
  xt_rsc_5_8_i_qa <= xt_rsc_5_8_qa;
  xt_rsc_5_8_da <= xt_rsc_5_8_i_da;
  xt_rsc_5_8_adra <= xt_rsc_5_8_i_adra;
  xt_rsc_5_8_i_adra_d <= xt_rsc_0_1_i_adra_d_iff;
  xt_rsc_5_8_i_da_d <= xt_rsc_4_8_i_da_d_iff;
  xt_rsc_5_8_i_qa_d <= xt_rsc_5_8_i_qa_d_1;

  xt_rsc_5_9_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_432_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_5_9_i_qa,
      wea => xt_rsc_5_9_wea,
      da => xt_rsc_5_9_i_da,
      adra => xt_rsc_5_9_i_adra,
      adra_d => xt_rsc_5_9_i_adra_d,
      da_d => xt_rsc_5_9_i_da_d,
      qa_d => xt_rsc_5_9_i_qa_d_1,
      wea_d => xt_rsc_1_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_0_i_wea_d_iff
    );
  xt_rsc_5_9_i_qa <= xt_rsc_5_9_qa;
  xt_rsc_5_9_da <= xt_rsc_5_9_i_da;
  xt_rsc_5_9_adra <= xt_rsc_5_9_i_adra;
  xt_rsc_5_9_i_adra_d <= xt_rsc_4_9_i_adra_d_iff;
  xt_rsc_5_9_i_da_d <= xt_rsc_4_9_i_da_d_iff;
  xt_rsc_5_9_i_qa_d <= xt_rsc_5_9_i_qa_d_1;

  xt_rsc_5_10_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_433_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_5_10_i_qa,
      wea => xt_rsc_5_10_wea,
      da => xt_rsc_5_10_i_da,
      adra => xt_rsc_5_10_i_adra,
      adra_d => xt_rsc_5_10_i_adra_d,
      da_d => xt_rsc_5_10_i_da_d,
      qa_d => xt_rsc_5_10_i_qa_d_1,
      wea_d => xt_rsc_1_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_0_i_wea_d_iff
    );
  xt_rsc_5_10_i_qa <= xt_rsc_5_10_qa;
  xt_rsc_5_10_da <= xt_rsc_5_10_i_da;
  xt_rsc_5_10_adra <= xt_rsc_5_10_i_adra;
  xt_rsc_5_10_i_adra_d <= xt_rsc_4_10_i_adra_d_iff;
  xt_rsc_5_10_i_da_d <= xt_rsc_4_10_i_da_d_iff;
  xt_rsc_5_10_i_qa_d <= xt_rsc_5_10_i_qa_d_1;

  xt_rsc_5_11_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_434_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_5_11_i_qa,
      wea => xt_rsc_5_11_wea,
      da => xt_rsc_5_11_i_da,
      adra => xt_rsc_5_11_i_adra,
      adra_d => xt_rsc_5_11_i_adra_d,
      da_d => xt_rsc_5_11_i_da_d,
      qa_d => xt_rsc_5_11_i_qa_d_1,
      wea_d => xt_rsc_1_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_0_i_wea_d_iff
    );
  xt_rsc_5_11_i_qa <= xt_rsc_5_11_qa;
  xt_rsc_5_11_da <= xt_rsc_5_11_i_da;
  xt_rsc_5_11_adra <= xt_rsc_5_11_i_adra;
  xt_rsc_5_11_i_adra_d <= xt_rsc_0_3_i_adra_d_iff;
  xt_rsc_5_11_i_da_d <= xt_rsc_4_11_i_da_d_iff;
  xt_rsc_5_11_i_qa_d <= xt_rsc_5_11_i_qa_d_1;

  xt_rsc_5_12_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_435_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_5_12_i_qa,
      wea => xt_rsc_5_12_wea,
      da => xt_rsc_5_12_i_da,
      adra => xt_rsc_5_12_i_adra,
      adra_d => xt_rsc_5_12_i_adra_d,
      da_d => xt_rsc_5_12_i_da_d,
      qa_d => xt_rsc_5_12_i_qa_d_1,
      wea_d => xt_rsc_1_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_0_i_wea_d_iff
    );
  xt_rsc_5_12_i_qa <= xt_rsc_5_12_qa;
  xt_rsc_5_12_da <= xt_rsc_5_12_i_da;
  xt_rsc_5_12_adra <= xt_rsc_5_12_i_adra;
  xt_rsc_5_12_i_adra_d <= xt_rsc_0_4_i_adra_d_iff;
  xt_rsc_5_12_i_da_d <= xt_rsc_4_12_i_da_d_iff;
  xt_rsc_5_12_i_qa_d <= xt_rsc_5_12_i_qa_d_1;

  xt_rsc_5_13_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_436_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_5_13_i_qa,
      wea => xt_rsc_5_13_wea,
      da => xt_rsc_5_13_i_da,
      adra => xt_rsc_5_13_i_adra,
      adra_d => xt_rsc_5_13_i_adra_d,
      da_d => xt_rsc_5_13_i_da_d,
      qa_d => xt_rsc_5_13_i_qa_d_1,
      wea_d => xt_rsc_1_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_0_i_wea_d_iff
    );
  xt_rsc_5_13_i_qa <= xt_rsc_5_13_qa;
  xt_rsc_5_13_da <= xt_rsc_5_13_i_da;
  xt_rsc_5_13_adra <= xt_rsc_5_13_i_adra;
  xt_rsc_5_13_i_adra_d <= xt_rsc_0_5_i_adra_d_iff;
  xt_rsc_5_13_i_da_d <= xt_rsc_4_13_i_da_d_iff;
  xt_rsc_5_13_i_qa_d <= xt_rsc_5_13_i_qa_d_1;

  xt_rsc_5_14_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_437_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_5_14_i_qa,
      wea => xt_rsc_5_14_wea,
      da => xt_rsc_5_14_i_da,
      adra => xt_rsc_5_14_i_adra,
      adra_d => xt_rsc_5_14_i_adra_d,
      da_d => xt_rsc_5_14_i_da_d,
      qa_d => xt_rsc_5_14_i_qa_d_1,
      wea_d => xt_rsc_1_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_0_i_wea_d_iff
    );
  xt_rsc_5_14_i_qa <= xt_rsc_5_14_qa;
  xt_rsc_5_14_da <= xt_rsc_5_14_i_da;
  xt_rsc_5_14_adra <= xt_rsc_5_14_i_adra;
  xt_rsc_5_14_i_adra_d <= xt_rsc_0_6_i_adra_d_iff;
  xt_rsc_5_14_i_da_d <= xt_rsc_4_14_i_da_d_iff;
  xt_rsc_5_14_i_qa_d <= xt_rsc_5_14_i_qa_d_1;

  xt_rsc_5_15_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_438_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_5_15_i_qa,
      wea => xt_rsc_5_15_wea,
      da => xt_rsc_5_15_i_da,
      adra => xt_rsc_5_15_i_adra,
      adra_d => xt_rsc_5_15_i_adra_d,
      da_d => xt_rsc_5_15_i_da_d,
      qa_d => xt_rsc_5_15_i_qa_d_1,
      wea_d => xt_rsc_1_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_0_i_wea_d_iff
    );
  xt_rsc_5_15_i_qa <= xt_rsc_5_15_qa;
  xt_rsc_5_15_da <= xt_rsc_5_15_i_da;
  xt_rsc_5_15_adra <= xt_rsc_5_15_i_adra;
  xt_rsc_5_15_i_adra_d <= xt_rsc_0_7_i_adra_d_iff;
  xt_rsc_5_15_i_da_d <= xt_rsc_4_15_i_da_d_iff;
  xt_rsc_5_15_i_qa_d <= xt_rsc_5_15_i_qa_d_1;

  xt_rsc_5_16_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_439_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_5_16_i_qa,
      wea => xt_rsc_5_16_wea,
      da => xt_rsc_5_16_i_da,
      adra => xt_rsc_5_16_i_adra,
      adra_d => xt_rsc_5_16_i_adra_d,
      da_d => xt_rsc_5_16_i_da_d,
      qa_d => xt_rsc_5_16_i_qa_d_1,
      wea_d => xt_rsc_1_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_16_i_wea_d_iff
    );
  xt_rsc_5_16_i_qa <= xt_rsc_5_16_qa;
  xt_rsc_5_16_da <= xt_rsc_5_16_i_da;
  xt_rsc_5_16_adra <= xt_rsc_5_16_i_adra;
  xt_rsc_5_16_i_adra_d <= xt_rsc_0_8_i_adra_d_iff;
  xt_rsc_5_16_i_da_d <= xt_rsc_4_0_i_da_d_iff;
  xt_rsc_5_16_i_qa_d <= xt_rsc_5_16_i_qa_d_1;

  xt_rsc_5_17_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_440_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_5_17_i_qa,
      wea => xt_rsc_5_17_wea,
      da => xt_rsc_5_17_i_da,
      adra => xt_rsc_5_17_i_adra,
      adra_d => xt_rsc_5_17_i_adra_d,
      da_d => xt_rsc_5_17_i_da_d,
      qa_d => xt_rsc_5_17_i_qa_d_1,
      wea_d => xt_rsc_1_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_16_i_wea_d_iff
    );
  xt_rsc_5_17_i_qa <= xt_rsc_5_17_qa;
  xt_rsc_5_17_da <= xt_rsc_5_17_i_da;
  xt_rsc_5_17_adra <= xt_rsc_5_17_i_adra;
  xt_rsc_5_17_i_adra_d <= xt_rsc_4_1_i_adra_d_iff;
  xt_rsc_5_17_i_da_d <= xt_rsc_4_1_i_da_d_iff;
  xt_rsc_5_17_i_qa_d <= xt_rsc_5_17_i_qa_d_1;

  xt_rsc_5_18_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_441_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_5_18_i_qa,
      wea => xt_rsc_5_18_wea,
      da => xt_rsc_5_18_i_da,
      adra => xt_rsc_5_18_i_adra,
      adra_d => xt_rsc_5_18_i_adra_d,
      da_d => xt_rsc_5_18_i_da_d,
      qa_d => xt_rsc_5_18_i_qa_d_1,
      wea_d => xt_rsc_1_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_16_i_wea_d_iff
    );
  xt_rsc_5_18_i_qa <= xt_rsc_5_18_qa;
  xt_rsc_5_18_da <= xt_rsc_5_18_i_da;
  xt_rsc_5_18_adra <= xt_rsc_5_18_i_adra;
  xt_rsc_5_18_i_adra_d <= xt_rsc_4_2_i_adra_d_iff;
  xt_rsc_5_18_i_da_d <= xt_rsc_4_2_i_da_d_iff;
  xt_rsc_5_18_i_qa_d <= xt_rsc_5_18_i_qa_d_1;

  xt_rsc_5_19_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_442_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_5_19_i_qa,
      wea => xt_rsc_5_19_wea,
      da => xt_rsc_5_19_i_da,
      adra => xt_rsc_5_19_i_adra,
      adra_d => xt_rsc_5_19_i_adra_d,
      da_d => xt_rsc_5_19_i_da_d,
      qa_d => xt_rsc_5_19_i_qa_d_1,
      wea_d => xt_rsc_1_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_16_i_wea_d_iff
    );
  xt_rsc_5_19_i_qa <= xt_rsc_5_19_qa;
  xt_rsc_5_19_da <= xt_rsc_5_19_i_da;
  xt_rsc_5_19_adra <= xt_rsc_5_19_i_adra;
  xt_rsc_5_19_i_adra_d <= xt_rsc_0_12_i_adra_d_iff;
  xt_rsc_5_19_i_da_d <= xt_rsc_4_3_i_da_d_iff;
  xt_rsc_5_19_i_qa_d <= xt_rsc_5_19_i_qa_d_1;

  xt_rsc_5_20_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_443_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_5_20_i_qa,
      wea => xt_rsc_5_20_wea,
      da => xt_rsc_5_20_i_da,
      adra => xt_rsc_5_20_i_adra,
      adra_d => xt_rsc_5_20_i_adra_d,
      da_d => xt_rsc_5_20_i_da_d,
      qa_d => xt_rsc_5_20_i_qa_d_1,
      wea_d => xt_rsc_1_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_16_i_wea_d_iff
    );
  xt_rsc_5_20_i_qa <= xt_rsc_5_20_qa;
  xt_rsc_5_20_da <= xt_rsc_5_20_i_da;
  xt_rsc_5_20_adra <= xt_rsc_5_20_i_adra;
  xt_rsc_5_20_i_adra_d <= xt_rsc_0_13_i_adra_d_iff;
  xt_rsc_5_20_i_da_d <= xt_rsc_4_4_i_da_d_iff;
  xt_rsc_5_20_i_qa_d <= xt_rsc_5_20_i_qa_d_1;

  xt_rsc_5_21_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_444_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_5_21_i_qa,
      wea => xt_rsc_5_21_wea,
      da => xt_rsc_5_21_i_da,
      adra => xt_rsc_5_21_i_adra,
      adra_d => xt_rsc_5_21_i_adra_d,
      da_d => xt_rsc_5_21_i_da_d,
      qa_d => xt_rsc_5_21_i_qa_d_1,
      wea_d => xt_rsc_1_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_16_i_wea_d_iff
    );
  xt_rsc_5_21_i_qa <= xt_rsc_5_21_qa;
  xt_rsc_5_21_da <= xt_rsc_5_21_i_da;
  xt_rsc_5_21_adra <= xt_rsc_5_21_i_adra;
  xt_rsc_5_21_i_adra_d <= xt_rsc_0_14_i_adra_d_iff;
  xt_rsc_5_21_i_da_d <= xt_rsc_4_5_i_da_d_iff;
  xt_rsc_5_21_i_qa_d <= xt_rsc_5_21_i_qa_d_1;

  xt_rsc_5_22_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_445_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_5_22_i_qa,
      wea => xt_rsc_5_22_wea,
      da => xt_rsc_5_22_i_da,
      adra => xt_rsc_5_22_i_adra,
      adra_d => xt_rsc_5_22_i_adra_d,
      da_d => xt_rsc_5_22_i_da_d,
      qa_d => xt_rsc_5_22_i_qa_d_1,
      wea_d => xt_rsc_1_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_16_i_wea_d_iff
    );
  xt_rsc_5_22_i_qa <= xt_rsc_5_22_qa;
  xt_rsc_5_22_da <= xt_rsc_5_22_i_da;
  xt_rsc_5_22_adra <= xt_rsc_5_22_i_adra;
  xt_rsc_5_22_i_adra_d <= xt_rsc_0_15_i_adra_d_iff;
  xt_rsc_5_22_i_da_d <= xt_rsc_4_6_i_da_d_iff;
  xt_rsc_5_22_i_qa_d <= xt_rsc_5_22_i_qa_d_1;

  xt_rsc_5_23_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_446_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_5_23_i_qa,
      wea => xt_rsc_5_23_wea,
      da => xt_rsc_5_23_i_da,
      adra => xt_rsc_5_23_i_adra,
      adra_d => xt_rsc_5_23_i_adra_d,
      da_d => xt_rsc_5_23_i_da_d,
      qa_d => xt_rsc_5_23_i_qa_d_1,
      wea_d => xt_rsc_1_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_16_i_wea_d_iff
    );
  xt_rsc_5_23_i_qa <= xt_rsc_5_23_qa;
  xt_rsc_5_23_da <= xt_rsc_5_23_i_da;
  xt_rsc_5_23_adra <= xt_rsc_5_23_i_adra;
  xt_rsc_5_23_i_adra_d <= xt_rsc_0_0_i_adra_d_iff;
  xt_rsc_5_23_i_da_d <= xt_rsc_4_7_i_da_d_iff;
  xt_rsc_5_23_i_qa_d <= xt_rsc_5_23_i_qa_d_1;

  xt_rsc_5_24_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_447_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_5_24_i_qa,
      wea => xt_rsc_5_24_wea,
      da => xt_rsc_5_24_i_da,
      adra => xt_rsc_5_24_i_adra,
      adra_d => xt_rsc_5_24_i_adra_d,
      da_d => xt_rsc_5_24_i_da_d,
      qa_d => xt_rsc_5_24_i_qa_d_1,
      wea_d => xt_rsc_1_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_16_i_wea_d_iff
    );
  xt_rsc_5_24_i_qa <= xt_rsc_5_24_qa;
  xt_rsc_5_24_da <= xt_rsc_5_24_i_da;
  xt_rsc_5_24_adra <= xt_rsc_5_24_i_adra;
  xt_rsc_5_24_i_adra_d <= xt_rsc_0_1_i_adra_d_iff;
  xt_rsc_5_24_i_da_d <= xt_rsc_4_8_i_da_d_iff;
  xt_rsc_5_24_i_qa_d <= xt_rsc_5_24_i_qa_d_1;

  xt_rsc_5_25_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_448_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_5_25_i_qa,
      wea => xt_rsc_5_25_wea,
      da => xt_rsc_5_25_i_da,
      adra => xt_rsc_5_25_i_adra,
      adra_d => xt_rsc_5_25_i_adra_d,
      da_d => xt_rsc_5_25_i_da_d,
      qa_d => xt_rsc_5_25_i_qa_d_1,
      wea_d => xt_rsc_1_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_16_i_wea_d_iff
    );
  xt_rsc_5_25_i_qa <= xt_rsc_5_25_qa;
  xt_rsc_5_25_da <= xt_rsc_5_25_i_da;
  xt_rsc_5_25_adra <= xt_rsc_5_25_i_adra;
  xt_rsc_5_25_i_adra_d <= xt_rsc_4_9_i_adra_d_iff;
  xt_rsc_5_25_i_da_d <= xt_rsc_4_9_i_da_d_iff;
  xt_rsc_5_25_i_qa_d <= xt_rsc_5_25_i_qa_d_1;

  xt_rsc_5_26_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_449_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_5_26_i_qa,
      wea => xt_rsc_5_26_wea,
      da => xt_rsc_5_26_i_da,
      adra => xt_rsc_5_26_i_adra,
      adra_d => xt_rsc_5_26_i_adra_d,
      da_d => xt_rsc_5_26_i_da_d,
      qa_d => xt_rsc_5_26_i_qa_d_1,
      wea_d => xt_rsc_1_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_16_i_wea_d_iff
    );
  xt_rsc_5_26_i_qa <= xt_rsc_5_26_qa;
  xt_rsc_5_26_da <= xt_rsc_5_26_i_da;
  xt_rsc_5_26_adra <= xt_rsc_5_26_i_adra;
  xt_rsc_5_26_i_adra_d <= xt_rsc_4_10_i_adra_d_iff;
  xt_rsc_5_26_i_da_d <= xt_rsc_4_10_i_da_d_iff;
  xt_rsc_5_26_i_qa_d <= xt_rsc_5_26_i_qa_d_1;

  xt_rsc_5_27_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_450_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_5_27_i_qa,
      wea => xt_rsc_5_27_wea,
      da => xt_rsc_5_27_i_da,
      adra => xt_rsc_5_27_i_adra,
      adra_d => xt_rsc_5_27_i_adra_d,
      da_d => xt_rsc_5_27_i_da_d,
      qa_d => xt_rsc_5_27_i_qa_d_1,
      wea_d => xt_rsc_1_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_16_i_wea_d_iff
    );
  xt_rsc_5_27_i_qa <= xt_rsc_5_27_qa;
  xt_rsc_5_27_da <= xt_rsc_5_27_i_da;
  xt_rsc_5_27_adra <= xt_rsc_5_27_i_adra;
  xt_rsc_5_27_i_adra_d <= xt_rsc_0_3_i_adra_d_iff;
  xt_rsc_5_27_i_da_d <= xt_rsc_4_11_i_da_d_iff;
  xt_rsc_5_27_i_qa_d <= xt_rsc_5_27_i_qa_d_1;

  xt_rsc_5_28_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_451_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_5_28_i_qa,
      wea => xt_rsc_5_28_wea,
      da => xt_rsc_5_28_i_da,
      adra => xt_rsc_5_28_i_adra,
      adra_d => xt_rsc_5_28_i_adra_d,
      da_d => xt_rsc_5_28_i_da_d,
      qa_d => xt_rsc_5_28_i_qa_d_1,
      wea_d => xt_rsc_1_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_16_i_wea_d_iff
    );
  xt_rsc_5_28_i_qa <= xt_rsc_5_28_qa;
  xt_rsc_5_28_da <= xt_rsc_5_28_i_da;
  xt_rsc_5_28_adra <= xt_rsc_5_28_i_adra;
  xt_rsc_5_28_i_adra_d <= xt_rsc_0_4_i_adra_d_iff;
  xt_rsc_5_28_i_da_d <= xt_rsc_4_12_i_da_d_iff;
  xt_rsc_5_28_i_qa_d <= xt_rsc_5_28_i_qa_d_1;

  xt_rsc_5_29_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_452_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_5_29_i_qa,
      wea => xt_rsc_5_29_wea,
      da => xt_rsc_5_29_i_da,
      adra => xt_rsc_5_29_i_adra,
      adra_d => xt_rsc_5_29_i_adra_d,
      da_d => xt_rsc_5_29_i_da_d,
      qa_d => xt_rsc_5_29_i_qa_d_1,
      wea_d => xt_rsc_1_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_16_i_wea_d_iff
    );
  xt_rsc_5_29_i_qa <= xt_rsc_5_29_qa;
  xt_rsc_5_29_da <= xt_rsc_5_29_i_da;
  xt_rsc_5_29_adra <= xt_rsc_5_29_i_adra;
  xt_rsc_5_29_i_adra_d <= xt_rsc_0_5_i_adra_d_iff;
  xt_rsc_5_29_i_da_d <= xt_rsc_4_13_i_da_d_iff;
  xt_rsc_5_29_i_qa_d <= xt_rsc_5_29_i_qa_d_1;

  xt_rsc_5_30_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_453_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_5_30_i_qa,
      wea => xt_rsc_5_30_wea,
      da => xt_rsc_5_30_i_da,
      adra => xt_rsc_5_30_i_adra,
      adra_d => xt_rsc_5_30_i_adra_d,
      da_d => xt_rsc_5_30_i_da_d,
      qa_d => xt_rsc_5_30_i_qa_d_1,
      wea_d => xt_rsc_1_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_16_i_wea_d_iff
    );
  xt_rsc_5_30_i_qa <= xt_rsc_5_30_qa;
  xt_rsc_5_30_da <= xt_rsc_5_30_i_da;
  xt_rsc_5_30_adra <= xt_rsc_5_30_i_adra;
  xt_rsc_5_30_i_adra_d <= xt_rsc_0_6_i_adra_d_iff;
  xt_rsc_5_30_i_da_d <= xt_rsc_4_14_i_da_d_iff;
  xt_rsc_5_30_i_qa_d <= xt_rsc_5_30_i_qa_d_1;

  xt_rsc_5_31_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_454_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_5_31_i_qa,
      wea => xt_rsc_5_31_wea,
      da => xt_rsc_5_31_i_da,
      adra => xt_rsc_5_31_i_adra,
      adra_d => xt_rsc_5_31_i_adra_d,
      da_d => xt_rsc_5_31_i_da_d,
      qa_d => xt_rsc_5_31_i_qa_d_1,
      wea_d => xt_rsc_1_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_16_i_wea_d_iff
    );
  xt_rsc_5_31_i_qa <= xt_rsc_5_31_qa;
  xt_rsc_5_31_da <= xt_rsc_5_31_i_da;
  xt_rsc_5_31_adra <= xt_rsc_5_31_i_adra;
  xt_rsc_5_31_i_adra_d <= xt_rsc_0_7_i_adra_d_iff;
  xt_rsc_5_31_i_da_d <= xt_rsc_4_15_i_da_d_iff;
  xt_rsc_5_31_i_qa_d <= xt_rsc_5_31_i_qa_d_1;

  xt_rsc_6_0_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_455_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_6_0_i_qa,
      wea => xt_rsc_6_0_wea,
      da => xt_rsc_6_0_i_da,
      adra => xt_rsc_6_0_i_adra,
      adra_d => xt_rsc_6_0_i_adra_d,
      da_d => xt_rsc_6_0_i_da_d,
      qa_d => xt_rsc_6_0_i_qa_d_1,
      wea_d => xt_rsc_2_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_2_0_i_wea_d_iff
    );
  xt_rsc_6_0_i_qa <= xt_rsc_6_0_qa;
  xt_rsc_6_0_da <= xt_rsc_6_0_i_da;
  xt_rsc_6_0_adra <= xt_rsc_6_0_i_adra;
  xt_rsc_6_0_i_adra_d <= xt_rsc_0_8_i_adra_d_iff;
  xt_rsc_6_0_i_da_d <= xt_rsc_4_0_i_da_d_iff;
  xt_rsc_6_0_i_qa_d <= xt_rsc_6_0_i_qa_d_1;

  xt_rsc_6_1_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_456_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_6_1_i_qa,
      wea => xt_rsc_6_1_wea,
      da => xt_rsc_6_1_i_da,
      adra => xt_rsc_6_1_i_adra,
      adra_d => xt_rsc_6_1_i_adra_d,
      da_d => xt_rsc_6_1_i_da_d,
      qa_d => xt_rsc_6_1_i_qa_d_1,
      wea_d => xt_rsc_2_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_2_0_i_wea_d_iff
    );
  xt_rsc_6_1_i_qa <= xt_rsc_6_1_qa;
  xt_rsc_6_1_da <= xt_rsc_6_1_i_da;
  xt_rsc_6_1_adra <= xt_rsc_6_1_i_adra;
  xt_rsc_6_1_i_adra_d <= xt_rsc_4_1_i_adra_d_iff;
  xt_rsc_6_1_i_da_d <= xt_rsc_4_1_i_da_d_iff;
  xt_rsc_6_1_i_qa_d <= xt_rsc_6_1_i_qa_d_1;

  xt_rsc_6_2_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_457_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_6_2_i_qa,
      wea => xt_rsc_6_2_wea,
      da => xt_rsc_6_2_i_da,
      adra => xt_rsc_6_2_i_adra,
      adra_d => xt_rsc_6_2_i_adra_d,
      da_d => xt_rsc_6_2_i_da_d,
      qa_d => xt_rsc_6_2_i_qa_d_1,
      wea_d => xt_rsc_2_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_2_0_i_wea_d_iff
    );
  xt_rsc_6_2_i_qa <= xt_rsc_6_2_qa;
  xt_rsc_6_2_da <= xt_rsc_6_2_i_da;
  xt_rsc_6_2_adra <= xt_rsc_6_2_i_adra;
  xt_rsc_6_2_i_adra_d <= xt_rsc_4_2_i_adra_d_iff;
  xt_rsc_6_2_i_da_d <= xt_rsc_4_2_i_da_d_iff;
  xt_rsc_6_2_i_qa_d <= xt_rsc_6_2_i_qa_d_1;

  xt_rsc_6_3_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_458_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_6_3_i_qa,
      wea => xt_rsc_6_3_wea,
      da => xt_rsc_6_3_i_da,
      adra => xt_rsc_6_3_i_adra,
      adra_d => xt_rsc_6_3_i_adra_d,
      da_d => xt_rsc_6_3_i_da_d,
      qa_d => xt_rsc_6_3_i_qa_d_1,
      wea_d => xt_rsc_2_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_2_0_i_wea_d_iff
    );
  xt_rsc_6_3_i_qa <= xt_rsc_6_3_qa;
  xt_rsc_6_3_da <= xt_rsc_6_3_i_da;
  xt_rsc_6_3_adra <= xt_rsc_6_3_i_adra;
  xt_rsc_6_3_i_adra_d <= xt_rsc_0_12_i_adra_d_iff;
  xt_rsc_6_3_i_da_d <= xt_rsc_4_3_i_da_d_iff;
  xt_rsc_6_3_i_qa_d <= xt_rsc_6_3_i_qa_d_1;

  xt_rsc_6_4_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_459_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_6_4_i_qa,
      wea => xt_rsc_6_4_wea,
      da => xt_rsc_6_4_i_da,
      adra => xt_rsc_6_4_i_adra,
      adra_d => xt_rsc_6_4_i_adra_d,
      da_d => xt_rsc_6_4_i_da_d,
      qa_d => xt_rsc_6_4_i_qa_d_1,
      wea_d => xt_rsc_2_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_2_0_i_wea_d_iff
    );
  xt_rsc_6_4_i_qa <= xt_rsc_6_4_qa;
  xt_rsc_6_4_da <= xt_rsc_6_4_i_da;
  xt_rsc_6_4_adra <= xt_rsc_6_4_i_adra;
  xt_rsc_6_4_i_adra_d <= xt_rsc_0_13_i_adra_d_iff;
  xt_rsc_6_4_i_da_d <= xt_rsc_4_4_i_da_d_iff;
  xt_rsc_6_4_i_qa_d <= xt_rsc_6_4_i_qa_d_1;

  xt_rsc_6_5_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_460_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_6_5_i_qa,
      wea => xt_rsc_6_5_wea,
      da => xt_rsc_6_5_i_da,
      adra => xt_rsc_6_5_i_adra,
      adra_d => xt_rsc_6_5_i_adra_d,
      da_d => xt_rsc_6_5_i_da_d,
      qa_d => xt_rsc_6_5_i_qa_d_1,
      wea_d => xt_rsc_2_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_2_0_i_wea_d_iff
    );
  xt_rsc_6_5_i_qa <= xt_rsc_6_5_qa;
  xt_rsc_6_5_da <= xt_rsc_6_5_i_da;
  xt_rsc_6_5_adra <= xt_rsc_6_5_i_adra;
  xt_rsc_6_5_i_adra_d <= xt_rsc_0_14_i_adra_d_iff;
  xt_rsc_6_5_i_da_d <= xt_rsc_4_5_i_da_d_iff;
  xt_rsc_6_5_i_qa_d <= xt_rsc_6_5_i_qa_d_1;

  xt_rsc_6_6_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_461_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_6_6_i_qa,
      wea => xt_rsc_6_6_wea,
      da => xt_rsc_6_6_i_da,
      adra => xt_rsc_6_6_i_adra,
      adra_d => xt_rsc_6_6_i_adra_d,
      da_d => xt_rsc_6_6_i_da_d,
      qa_d => xt_rsc_6_6_i_qa_d_1,
      wea_d => xt_rsc_2_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_2_0_i_wea_d_iff
    );
  xt_rsc_6_6_i_qa <= xt_rsc_6_6_qa;
  xt_rsc_6_6_da <= xt_rsc_6_6_i_da;
  xt_rsc_6_6_adra <= xt_rsc_6_6_i_adra;
  xt_rsc_6_6_i_adra_d <= xt_rsc_0_15_i_adra_d_iff;
  xt_rsc_6_6_i_da_d <= xt_rsc_4_6_i_da_d_iff;
  xt_rsc_6_6_i_qa_d <= xt_rsc_6_6_i_qa_d_1;

  xt_rsc_6_7_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_462_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_6_7_i_qa,
      wea => xt_rsc_6_7_wea,
      da => xt_rsc_6_7_i_da,
      adra => xt_rsc_6_7_i_adra,
      adra_d => xt_rsc_6_7_i_adra_d,
      da_d => xt_rsc_6_7_i_da_d,
      qa_d => xt_rsc_6_7_i_qa_d_1,
      wea_d => xt_rsc_2_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_2_0_i_wea_d_iff
    );
  xt_rsc_6_7_i_qa <= xt_rsc_6_7_qa;
  xt_rsc_6_7_da <= xt_rsc_6_7_i_da;
  xt_rsc_6_7_adra <= xt_rsc_6_7_i_adra;
  xt_rsc_6_7_i_adra_d <= xt_rsc_0_0_i_adra_d_iff;
  xt_rsc_6_7_i_da_d <= xt_rsc_4_7_i_da_d_iff;
  xt_rsc_6_7_i_qa_d <= xt_rsc_6_7_i_qa_d_1;

  xt_rsc_6_8_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_463_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_6_8_i_qa,
      wea => xt_rsc_6_8_wea,
      da => xt_rsc_6_8_i_da,
      adra => xt_rsc_6_8_i_adra,
      adra_d => xt_rsc_6_8_i_adra_d,
      da_d => xt_rsc_6_8_i_da_d,
      qa_d => xt_rsc_6_8_i_qa_d_1,
      wea_d => xt_rsc_2_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_2_0_i_wea_d_iff
    );
  xt_rsc_6_8_i_qa <= xt_rsc_6_8_qa;
  xt_rsc_6_8_da <= xt_rsc_6_8_i_da;
  xt_rsc_6_8_adra <= xt_rsc_6_8_i_adra;
  xt_rsc_6_8_i_adra_d <= xt_rsc_0_1_i_adra_d_iff;
  xt_rsc_6_8_i_da_d <= xt_rsc_4_8_i_da_d_iff;
  xt_rsc_6_8_i_qa_d <= xt_rsc_6_8_i_qa_d_1;

  xt_rsc_6_9_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_464_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_6_9_i_qa,
      wea => xt_rsc_6_9_wea,
      da => xt_rsc_6_9_i_da,
      adra => xt_rsc_6_9_i_adra,
      adra_d => xt_rsc_6_9_i_adra_d,
      da_d => xt_rsc_6_9_i_da_d,
      qa_d => xt_rsc_6_9_i_qa_d_1,
      wea_d => xt_rsc_2_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_2_0_i_wea_d_iff
    );
  xt_rsc_6_9_i_qa <= xt_rsc_6_9_qa;
  xt_rsc_6_9_da <= xt_rsc_6_9_i_da;
  xt_rsc_6_9_adra <= xt_rsc_6_9_i_adra;
  xt_rsc_6_9_i_adra_d <= xt_rsc_4_9_i_adra_d_iff;
  xt_rsc_6_9_i_da_d <= xt_rsc_4_9_i_da_d_iff;
  xt_rsc_6_9_i_qa_d <= xt_rsc_6_9_i_qa_d_1;

  xt_rsc_6_10_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_465_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_6_10_i_qa,
      wea => xt_rsc_6_10_wea,
      da => xt_rsc_6_10_i_da,
      adra => xt_rsc_6_10_i_adra,
      adra_d => xt_rsc_6_10_i_adra_d,
      da_d => xt_rsc_6_10_i_da_d,
      qa_d => xt_rsc_6_10_i_qa_d_1,
      wea_d => xt_rsc_2_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_2_0_i_wea_d_iff
    );
  xt_rsc_6_10_i_qa <= xt_rsc_6_10_qa;
  xt_rsc_6_10_da <= xt_rsc_6_10_i_da;
  xt_rsc_6_10_adra <= xt_rsc_6_10_i_adra;
  xt_rsc_6_10_i_adra_d <= xt_rsc_4_10_i_adra_d_iff;
  xt_rsc_6_10_i_da_d <= xt_rsc_4_10_i_da_d_iff;
  xt_rsc_6_10_i_qa_d <= xt_rsc_6_10_i_qa_d_1;

  xt_rsc_6_11_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_466_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_6_11_i_qa,
      wea => xt_rsc_6_11_wea,
      da => xt_rsc_6_11_i_da,
      adra => xt_rsc_6_11_i_adra,
      adra_d => xt_rsc_6_11_i_adra_d,
      da_d => xt_rsc_6_11_i_da_d,
      qa_d => xt_rsc_6_11_i_qa_d_1,
      wea_d => xt_rsc_2_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_2_0_i_wea_d_iff
    );
  xt_rsc_6_11_i_qa <= xt_rsc_6_11_qa;
  xt_rsc_6_11_da <= xt_rsc_6_11_i_da;
  xt_rsc_6_11_adra <= xt_rsc_6_11_i_adra;
  xt_rsc_6_11_i_adra_d <= xt_rsc_0_3_i_adra_d_iff;
  xt_rsc_6_11_i_da_d <= xt_rsc_4_11_i_da_d_iff;
  xt_rsc_6_11_i_qa_d <= xt_rsc_6_11_i_qa_d_1;

  xt_rsc_6_12_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_467_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_6_12_i_qa,
      wea => xt_rsc_6_12_wea,
      da => xt_rsc_6_12_i_da,
      adra => xt_rsc_6_12_i_adra,
      adra_d => xt_rsc_6_12_i_adra_d,
      da_d => xt_rsc_6_12_i_da_d,
      qa_d => xt_rsc_6_12_i_qa_d_1,
      wea_d => xt_rsc_2_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_2_0_i_wea_d_iff
    );
  xt_rsc_6_12_i_qa <= xt_rsc_6_12_qa;
  xt_rsc_6_12_da <= xt_rsc_6_12_i_da;
  xt_rsc_6_12_adra <= xt_rsc_6_12_i_adra;
  xt_rsc_6_12_i_adra_d <= xt_rsc_0_4_i_adra_d_iff;
  xt_rsc_6_12_i_da_d <= xt_rsc_4_12_i_da_d_iff;
  xt_rsc_6_12_i_qa_d <= xt_rsc_6_12_i_qa_d_1;

  xt_rsc_6_13_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_468_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_6_13_i_qa,
      wea => xt_rsc_6_13_wea,
      da => xt_rsc_6_13_i_da,
      adra => xt_rsc_6_13_i_adra,
      adra_d => xt_rsc_6_13_i_adra_d,
      da_d => xt_rsc_6_13_i_da_d,
      qa_d => xt_rsc_6_13_i_qa_d_1,
      wea_d => xt_rsc_2_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_2_0_i_wea_d_iff
    );
  xt_rsc_6_13_i_qa <= xt_rsc_6_13_qa;
  xt_rsc_6_13_da <= xt_rsc_6_13_i_da;
  xt_rsc_6_13_adra <= xt_rsc_6_13_i_adra;
  xt_rsc_6_13_i_adra_d <= xt_rsc_0_5_i_adra_d_iff;
  xt_rsc_6_13_i_da_d <= xt_rsc_4_13_i_da_d_iff;
  xt_rsc_6_13_i_qa_d <= xt_rsc_6_13_i_qa_d_1;

  xt_rsc_6_14_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_469_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_6_14_i_qa,
      wea => xt_rsc_6_14_wea,
      da => xt_rsc_6_14_i_da,
      adra => xt_rsc_6_14_i_adra,
      adra_d => xt_rsc_6_14_i_adra_d,
      da_d => xt_rsc_6_14_i_da_d,
      qa_d => xt_rsc_6_14_i_qa_d_1,
      wea_d => xt_rsc_2_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_2_0_i_wea_d_iff
    );
  xt_rsc_6_14_i_qa <= xt_rsc_6_14_qa;
  xt_rsc_6_14_da <= xt_rsc_6_14_i_da;
  xt_rsc_6_14_adra <= xt_rsc_6_14_i_adra;
  xt_rsc_6_14_i_adra_d <= xt_rsc_0_6_i_adra_d_iff;
  xt_rsc_6_14_i_da_d <= xt_rsc_4_14_i_da_d_iff;
  xt_rsc_6_14_i_qa_d <= xt_rsc_6_14_i_qa_d_1;

  xt_rsc_6_15_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_470_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_6_15_i_qa,
      wea => xt_rsc_6_15_wea,
      da => xt_rsc_6_15_i_da,
      adra => xt_rsc_6_15_i_adra,
      adra_d => xt_rsc_6_15_i_adra_d,
      da_d => xt_rsc_6_15_i_da_d,
      qa_d => xt_rsc_6_15_i_qa_d_1,
      wea_d => xt_rsc_2_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_2_0_i_wea_d_iff
    );
  xt_rsc_6_15_i_qa <= xt_rsc_6_15_qa;
  xt_rsc_6_15_da <= xt_rsc_6_15_i_da;
  xt_rsc_6_15_adra <= xt_rsc_6_15_i_adra;
  xt_rsc_6_15_i_adra_d <= xt_rsc_0_7_i_adra_d_iff;
  xt_rsc_6_15_i_da_d <= xt_rsc_4_15_i_da_d_iff;
  xt_rsc_6_15_i_qa_d <= xt_rsc_6_15_i_qa_d_1;

  xt_rsc_6_16_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_471_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_6_16_i_qa,
      wea => xt_rsc_6_16_wea,
      da => xt_rsc_6_16_i_da,
      adra => xt_rsc_6_16_i_adra,
      adra_d => xt_rsc_6_16_i_adra_d,
      da_d => xt_rsc_6_16_i_da_d,
      qa_d => xt_rsc_6_16_i_qa_d_1,
      wea_d => xt_rsc_2_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_2_16_i_wea_d_iff
    );
  xt_rsc_6_16_i_qa <= xt_rsc_6_16_qa;
  xt_rsc_6_16_da <= xt_rsc_6_16_i_da;
  xt_rsc_6_16_adra <= xt_rsc_6_16_i_adra;
  xt_rsc_6_16_i_adra_d <= xt_rsc_0_8_i_adra_d_iff;
  xt_rsc_6_16_i_da_d <= xt_rsc_4_0_i_da_d_iff;
  xt_rsc_6_16_i_qa_d <= xt_rsc_6_16_i_qa_d_1;

  xt_rsc_6_17_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_472_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_6_17_i_qa,
      wea => xt_rsc_6_17_wea,
      da => xt_rsc_6_17_i_da,
      adra => xt_rsc_6_17_i_adra,
      adra_d => xt_rsc_6_17_i_adra_d,
      da_d => xt_rsc_6_17_i_da_d,
      qa_d => xt_rsc_6_17_i_qa_d_1,
      wea_d => xt_rsc_2_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_2_16_i_wea_d_iff
    );
  xt_rsc_6_17_i_qa <= xt_rsc_6_17_qa;
  xt_rsc_6_17_da <= xt_rsc_6_17_i_da;
  xt_rsc_6_17_adra <= xt_rsc_6_17_i_adra;
  xt_rsc_6_17_i_adra_d <= xt_rsc_4_1_i_adra_d_iff;
  xt_rsc_6_17_i_da_d <= xt_rsc_4_1_i_da_d_iff;
  xt_rsc_6_17_i_qa_d <= xt_rsc_6_17_i_qa_d_1;

  xt_rsc_6_18_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_473_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_6_18_i_qa,
      wea => xt_rsc_6_18_wea,
      da => xt_rsc_6_18_i_da,
      adra => xt_rsc_6_18_i_adra,
      adra_d => xt_rsc_6_18_i_adra_d,
      da_d => xt_rsc_6_18_i_da_d,
      qa_d => xt_rsc_6_18_i_qa_d_1,
      wea_d => xt_rsc_2_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_2_16_i_wea_d_iff
    );
  xt_rsc_6_18_i_qa <= xt_rsc_6_18_qa;
  xt_rsc_6_18_da <= xt_rsc_6_18_i_da;
  xt_rsc_6_18_adra <= xt_rsc_6_18_i_adra;
  xt_rsc_6_18_i_adra_d <= xt_rsc_4_2_i_adra_d_iff;
  xt_rsc_6_18_i_da_d <= xt_rsc_4_2_i_da_d_iff;
  xt_rsc_6_18_i_qa_d <= xt_rsc_6_18_i_qa_d_1;

  xt_rsc_6_19_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_474_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_6_19_i_qa,
      wea => xt_rsc_6_19_wea,
      da => xt_rsc_6_19_i_da,
      adra => xt_rsc_6_19_i_adra,
      adra_d => xt_rsc_6_19_i_adra_d,
      da_d => xt_rsc_6_19_i_da_d,
      qa_d => xt_rsc_6_19_i_qa_d_1,
      wea_d => xt_rsc_2_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_2_16_i_wea_d_iff
    );
  xt_rsc_6_19_i_qa <= xt_rsc_6_19_qa;
  xt_rsc_6_19_da <= xt_rsc_6_19_i_da;
  xt_rsc_6_19_adra <= xt_rsc_6_19_i_adra;
  xt_rsc_6_19_i_adra_d <= xt_rsc_0_12_i_adra_d_iff;
  xt_rsc_6_19_i_da_d <= xt_rsc_4_3_i_da_d_iff;
  xt_rsc_6_19_i_qa_d <= xt_rsc_6_19_i_qa_d_1;

  xt_rsc_6_20_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_475_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_6_20_i_qa,
      wea => xt_rsc_6_20_wea,
      da => xt_rsc_6_20_i_da,
      adra => xt_rsc_6_20_i_adra,
      adra_d => xt_rsc_6_20_i_adra_d,
      da_d => xt_rsc_6_20_i_da_d,
      qa_d => xt_rsc_6_20_i_qa_d_1,
      wea_d => xt_rsc_2_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_2_16_i_wea_d_iff
    );
  xt_rsc_6_20_i_qa <= xt_rsc_6_20_qa;
  xt_rsc_6_20_da <= xt_rsc_6_20_i_da;
  xt_rsc_6_20_adra <= xt_rsc_6_20_i_adra;
  xt_rsc_6_20_i_adra_d <= xt_rsc_0_13_i_adra_d_iff;
  xt_rsc_6_20_i_da_d <= xt_rsc_4_4_i_da_d_iff;
  xt_rsc_6_20_i_qa_d <= xt_rsc_6_20_i_qa_d_1;

  xt_rsc_6_21_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_476_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_6_21_i_qa,
      wea => xt_rsc_6_21_wea,
      da => xt_rsc_6_21_i_da,
      adra => xt_rsc_6_21_i_adra,
      adra_d => xt_rsc_6_21_i_adra_d,
      da_d => xt_rsc_6_21_i_da_d,
      qa_d => xt_rsc_6_21_i_qa_d_1,
      wea_d => xt_rsc_2_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_2_16_i_wea_d_iff
    );
  xt_rsc_6_21_i_qa <= xt_rsc_6_21_qa;
  xt_rsc_6_21_da <= xt_rsc_6_21_i_da;
  xt_rsc_6_21_adra <= xt_rsc_6_21_i_adra;
  xt_rsc_6_21_i_adra_d <= xt_rsc_0_14_i_adra_d_iff;
  xt_rsc_6_21_i_da_d <= xt_rsc_4_5_i_da_d_iff;
  xt_rsc_6_21_i_qa_d <= xt_rsc_6_21_i_qa_d_1;

  xt_rsc_6_22_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_477_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_6_22_i_qa,
      wea => xt_rsc_6_22_wea,
      da => xt_rsc_6_22_i_da,
      adra => xt_rsc_6_22_i_adra,
      adra_d => xt_rsc_6_22_i_adra_d,
      da_d => xt_rsc_6_22_i_da_d,
      qa_d => xt_rsc_6_22_i_qa_d_1,
      wea_d => xt_rsc_2_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_2_16_i_wea_d_iff
    );
  xt_rsc_6_22_i_qa <= xt_rsc_6_22_qa;
  xt_rsc_6_22_da <= xt_rsc_6_22_i_da;
  xt_rsc_6_22_adra <= xt_rsc_6_22_i_adra;
  xt_rsc_6_22_i_adra_d <= xt_rsc_0_15_i_adra_d_iff;
  xt_rsc_6_22_i_da_d <= xt_rsc_4_6_i_da_d_iff;
  xt_rsc_6_22_i_qa_d <= xt_rsc_6_22_i_qa_d_1;

  xt_rsc_6_23_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_478_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_6_23_i_qa,
      wea => xt_rsc_6_23_wea,
      da => xt_rsc_6_23_i_da,
      adra => xt_rsc_6_23_i_adra,
      adra_d => xt_rsc_6_23_i_adra_d,
      da_d => xt_rsc_6_23_i_da_d,
      qa_d => xt_rsc_6_23_i_qa_d_1,
      wea_d => xt_rsc_2_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_2_16_i_wea_d_iff
    );
  xt_rsc_6_23_i_qa <= xt_rsc_6_23_qa;
  xt_rsc_6_23_da <= xt_rsc_6_23_i_da;
  xt_rsc_6_23_adra <= xt_rsc_6_23_i_adra;
  xt_rsc_6_23_i_adra_d <= xt_rsc_0_0_i_adra_d_iff;
  xt_rsc_6_23_i_da_d <= xt_rsc_4_7_i_da_d_iff;
  xt_rsc_6_23_i_qa_d <= xt_rsc_6_23_i_qa_d_1;

  xt_rsc_6_24_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_479_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_6_24_i_qa,
      wea => xt_rsc_6_24_wea,
      da => xt_rsc_6_24_i_da,
      adra => xt_rsc_6_24_i_adra,
      adra_d => xt_rsc_6_24_i_adra_d,
      da_d => xt_rsc_6_24_i_da_d,
      qa_d => xt_rsc_6_24_i_qa_d_1,
      wea_d => xt_rsc_2_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_2_16_i_wea_d_iff
    );
  xt_rsc_6_24_i_qa <= xt_rsc_6_24_qa;
  xt_rsc_6_24_da <= xt_rsc_6_24_i_da;
  xt_rsc_6_24_adra <= xt_rsc_6_24_i_adra;
  xt_rsc_6_24_i_adra_d <= xt_rsc_0_1_i_adra_d_iff;
  xt_rsc_6_24_i_da_d <= xt_rsc_4_8_i_da_d_iff;
  xt_rsc_6_24_i_qa_d <= xt_rsc_6_24_i_qa_d_1;

  xt_rsc_6_25_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_480_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_6_25_i_qa,
      wea => xt_rsc_6_25_wea,
      da => xt_rsc_6_25_i_da,
      adra => xt_rsc_6_25_i_adra,
      adra_d => xt_rsc_6_25_i_adra_d,
      da_d => xt_rsc_6_25_i_da_d,
      qa_d => xt_rsc_6_25_i_qa_d_1,
      wea_d => xt_rsc_2_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_2_16_i_wea_d_iff
    );
  xt_rsc_6_25_i_qa <= xt_rsc_6_25_qa;
  xt_rsc_6_25_da <= xt_rsc_6_25_i_da;
  xt_rsc_6_25_adra <= xt_rsc_6_25_i_adra;
  xt_rsc_6_25_i_adra_d <= xt_rsc_4_9_i_adra_d_iff;
  xt_rsc_6_25_i_da_d <= xt_rsc_4_9_i_da_d_iff;
  xt_rsc_6_25_i_qa_d <= xt_rsc_6_25_i_qa_d_1;

  xt_rsc_6_26_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_481_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_6_26_i_qa,
      wea => xt_rsc_6_26_wea,
      da => xt_rsc_6_26_i_da,
      adra => xt_rsc_6_26_i_adra,
      adra_d => xt_rsc_6_26_i_adra_d,
      da_d => xt_rsc_6_26_i_da_d,
      qa_d => xt_rsc_6_26_i_qa_d_1,
      wea_d => xt_rsc_2_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_2_16_i_wea_d_iff
    );
  xt_rsc_6_26_i_qa <= xt_rsc_6_26_qa;
  xt_rsc_6_26_da <= xt_rsc_6_26_i_da;
  xt_rsc_6_26_adra <= xt_rsc_6_26_i_adra;
  xt_rsc_6_26_i_adra_d <= xt_rsc_4_10_i_adra_d_iff;
  xt_rsc_6_26_i_da_d <= xt_rsc_4_10_i_da_d_iff;
  xt_rsc_6_26_i_qa_d <= xt_rsc_6_26_i_qa_d_1;

  xt_rsc_6_27_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_482_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_6_27_i_qa,
      wea => xt_rsc_6_27_wea,
      da => xt_rsc_6_27_i_da,
      adra => xt_rsc_6_27_i_adra,
      adra_d => xt_rsc_6_27_i_adra_d,
      da_d => xt_rsc_6_27_i_da_d,
      qa_d => xt_rsc_6_27_i_qa_d_1,
      wea_d => xt_rsc_2_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_2_16_i_wea_d_iff
    );
  xt_rsc_6_27_i_qa <= xt_rsc_6_27_qa;
  xt_rsc_6_27_da <= xt_rsc_6_27_i_da;
  xt_rsc_6_27_adra <= xt_rsc_6_27_i_adra;
  xt_rsc_6_27_i_adra_d <= xt_rsc_0_3_i_adra_d_iff;
  xt_rsc_6_27_i_da_d <= xt_rsc_4_11_i_da_d_iff;
  xt_rsc_6_27_i_qa_d <= xt_rsc_6_27_i_qa_d_1;

  xt_rsc_6_28_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_483_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_6_28_i_qa,
      wea => xt_rsc_6_28_wea,
      da => xt_rsc_6_28_i_da,
      adra => xt_rsc_6_28_i_adra,
      adra_d => xt_rsc_6_28_i_adra_d,
      da_d => xt_rsc_6_28_i_da_d,
      qa_d => xt_rsc_6_28_i_qa_d_1,
      wea_d => xt_rsc_2_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_2_16_i_wea_d_iff
    );
  xt_rsc_6_28_i_qa <= xt_rsc_6_28_qa;
  xt_rsc_6_28_da <= xt_rsc_6_28_i_da;
  xt_rsc_6_28_adra <= xt_rsc_6_28_i_adra;
  xt_rsc_6_28_i_adra_d <= xt_rsc_0_4_i_adra_d_iff;
  xt_rsc_6_28_i_da_d <= xt_rsc_4_12_i_da_d_iff;
  xt_rsc_6_28_i_qa_d <= xt_rsc_6_28_i_qa_d_1;

  xt_rsc_6_29_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_484_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_6_29_i_qa,
      wea => xt_rsc_6_29_wea,
      da => xt_rsc_6_29_i_da,
      adra => xt_rsc_6_29_i_adra,
      adra_d => xt_rsc_6_29_i_adra_d,
      da_d => xt_rsc_6_29_i_da_d,
      qa_d => xt_rsc_6_29_i_qa_d_1,
      wea_d => xt_rsc_2_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_2_16_i_wea_d_iff
    );
  xt_rsc_6_29_i_qa <= xt_rsc_6_29_qa;
  xt_rsc_6_29_da <= xt_rsc_6_29_i_da;
  xt_rsc_6_29_adra <= xt_rsc_6_29_i_adra;
  xt_rsc_6_29_i_adra_d <= xt_rsc_0_5_i_adra_d_iff;
  xt_rsc_6_29_i_da_d <= xt_rsc_4_13_i_da_d_iff;
  xt_rsc_6_29_i_qa_d <= xt_rsc_6_29_i_qa_d_1;

  xt_rsc_6_30_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_485_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_6_30_i_qa,
      wea => xt_rsc_6_30_wea,
      da => xt_rsc_6_30_i_da,
      adra => xt_rsc_6_30_i_adra,
      adra_d => xt_rsc_6_30_i_adra_d,
      da_d => xt_rsc_6_30_i_da_d,
      qa_d => xt_rsc_6_30_i_qa_d_1,
      wea_d => xt_rsc_2_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_2_16_i_wea_d_iff
    );
  xt_rsc_6_30_i_qa <= xt_rsc_6_30_qa;
  xt_rsc_6_30_da <= xt_rsc_6_30_i_da;
  xt_rsc_6_30_adra <= xt_rsc_6_30_i_adra;
  xt_rsc_6_30_i_adra_d <= xt_rsc_0_6_i_adra_d_iff;
  xt_rsc_6_30_i_da_d <= xt_rsc_4_14_i_da_d_iff;
  xt_rsc_6_30_i_qa_d <= xt_rsc_6_30_i_qa_d_1;

  xt_rsc_6_31_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_486_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_6_31_i_qa,
      wea => xt_rsc_6_31_wea,
      da => xt_rsc_6_31_i_da,
      adra => xt_rsc_6_31_i_adra,
      adra_d => xt_rsc_6_31_i_adra_d,
      da_d => xt_rsc_6_31_i_da_d,
      qa_d => xt_rsc_6_31_i_qa_d_1,
      wea_d => xt_rsc_2_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_2_16_i_wea_d_iff
    );
  xt_rsc_6_31_i_qa <= xt_rsc_6_31_qa;
  xt_rsc_6_31_da <= xt_rsc_6_31_i_da;
  xt_rsc_6_31_adra <= xt_rsc_6_31_i_adra;
  xt_rsc_6_31_i_adra_d <= xt_rsc_0_7_i_adra_d_iff;
  xt_rsc_6_31_i_da_d <= xt_rsc_4_15_i_da_d_iff;
  xt_rsc_6_31_i_qa_d <= xt_rsc_6_31_i_qa_d_1;

  xt_rsc_7_0_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_487_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_7_0_i_qa,
      wea => xt_rsc_7_0_wea,
      da => xt_rsc_7_0_i_da,
      adra => xt_rsc_7_0_i_adra,
      adra_d => xt_rsc_7_0_i_adra_d,
      da_d => xt_rsc_7_0_i_da_d,
      qa_d => xt_rsc_7_0_i_qa_d_1,
      wea_d => xt_rsc_3_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_3_0_i_wea_d_iff
    );
  xt_rsc_7_0_i_qa <= xt_rsc_7_0_qa;
  xt_rsc_7_0_da <= xt_rsc_7_0_i_da;
  xt_rsc_7_0_adra <= xt_rsc_7_0_i_adra;
  xt_rsc_7_0_i_adra_d <= xt_rsc_0_8_i_adra_d_iff;
  xt_rsc_7_0_i_da_d <= xt_rsc_4_0_i_da_d_iff;
  xt_rsc_7_0_i_qa_d <= xt_rsc_7_0_i_qa_d_1;

  xt_rsc_7_1_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_488_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_7_1_i_qa,
      wea => xt_rsc_7_1_wea,
      da => xt_rsc_7_1_i_da,
      adra => xt_rsc_7_1_i_adra,
      adra_d => xt_rsc_7_1_i_adra_d,
      da_d => xt_rsc_7_1_i_da_d,
      qa_d => xt_rsc_7_1_i_qa_d_1,
      wea_d => xt_rsc_3_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_3_0_i_wea_d_iff
    );
  xt_rsc_7_1_i_qa <= xt_rsc_7_1_qa;
  xt_rsc_7_1_da <= xt_rsc_7_1_i_da;
  xt_rsc_7_1_adra <= xt_rsc_7_1_i_adra;
  xt_rsc_7_1_i_adra_d <= xt_rsc_4_1_i_adra_d_iff;
  xt_rsc_7_1_i_da_d <= xt_rsc_4_1_i_da_d_iff;
  xt_rsc_7_1_i_qa_d <= xt_rsc_7_1_i_qa_d_1;

  xt_rsc_7_2_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_489_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_7_2_i_qa,
      wea => xt_rsc_7_2_wea,
      da => xt_rsc_7_2_i_da,
      adra => xt_rsc_7_2_i_adra,
      adra_d => xt_rsc_7_2_i_adra_d,
      da_d => xt_rsc_7_2_i_da_d,
      qa_d => xt_rsc_7_2_i_qa_d_1,
      wea_d => xt_rsc_3_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_3_0_i_wea_d_iff
    );
  xt_rsc_7_2_i_qa <= xt_rsc_7_2_qa;
  xt_rsc_7_2_da <= xt_rsc_7_2_i_da;
  xt_rsc_7_2_adra <= xt_rsc_7_2_i_adra;
  xt_rsc_7_2_i_adra_d <= xt_rsc_4_2_i_adra_d_iff;
  xt_rsc_7_2_i_da_d <= xt_rsc_4_2_i_da_d_iff;
  xt_rsc_7_2_i_qa_d <= xt_rsc_7_2_i_qa_d_1;

  xt_rsc_7_3_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_490_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_7_3_i_qa,
      wea => xt_rsc_7_3_wea,
      da => xt_rsc_7_3_i_da,
      adra => xt_rsc_7_3_i_adra,
      adra_d => xt_rsc_7_3_i_adra_d,
      da_d => xt_rsc_7_3_i_da_d,
      qa_d => xt_rsc_7_3_i_qa_d_1,
      wea_d => xt_rsc_3_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_3_0_i_wea_d_iff
    );
  xt_rsc_7_3_i_qa <= xt_rsc_7_3_qa;
  xt_rsc_7_3_da <= xt_rsc_7_3_i_da;
  xt_rsc_7_3_adra <= xt_rsc_7_3_i_adra;
  xt_rsc_7_3_i_adra_d <= xt_rsc_0_12_i_adra_d_iff;
  xt_rsc_7_3_i_da_d <= xt_rsc_4_3_i_da_d_iff;
  xt_rsc_7_3_i_qa_d <= xt_rsc_7_3_i_qa_d_1;

  xt_rsc_7_4_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_491_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_7_4_i_qa,
      wea => xt_rsc_7_4_wea,
      da => xt_rsc_7_4_i_da,
      adra => xt_rsc_7_4_i_adra,
      adra_d => xt_rsc_7_4_i_adra_d,
      da_d => xt_rsc_7_4_i_da_d,
      qa_d => xt_rsc_7_4_i_qa_d_1,
      wea_d => xt_rsc_3_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_3_0_i_wea_d_iff
    );
  xt_rsc_7_4_i_qa <= xt_rsc_7_4_qa;
  xt_rsc_7_4_da <= xt_rsc_7_4_i_da;
  xt_rsc_7_4_adra <= xt_rsc_7_4_i_adra;
  xt_rsc_7_4_i_adra_d <= xt_rsc_0_13_i_adra_d_iff;
  xt_rsc_7_4_i_da_d <= xt_rsc_4_4_i_da_d_iff;
  xt_rsc_7_4_i_qa_d <= xt_rsc_7_4_i_qa_d_1;

  xt_rsc_7_5_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_492_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_7_5_i_qa,
      wea => xt_rsc_7_5_wea,
      da => xt_rsc_7_5_i_da,
      adra => xt_rsc_7_5_i_adra,
      adra_d => xt_rsc_7_5_i_adra_d,
      da_d => xt_rsc_7_5_i_da_d,
      qa_d => xt_rsc_7_5_i_qa_d_1,
      wea_d => xt_rsc_3_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_3_0_i_wea_d_iff
    );
  xt_rsc_7_5_i_qa <= xt_rsc_7_5_qa;
  xt_rsc_7_5_da <= xt_rsc_7_5_i_da;
  xt_rsc_7_5_adra <= xt_rsc_7_5_i_adra;
  xt_rsc_7_5_i_adra_d <= xt_rsc_0_14_i_adra_d_iff;
  xt_rsc_7_5_i_da_d <= xt_rsc_4_5_i_da_d_iff;
  xt_rsc_7_5_i_qa_d <= xt_rsc_7_5_i_qa_d_1;

  xt_rsc_7_6_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_493_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_7_6_i_qa,
      wea => xt_rsc_7_6_wea,
      da => xt_rsc_7_6_i_da,
      adra => xt_rsc_7_6_i_adra,
      adra_d => xt_rsc_7_6_i_adra_d,
      da_d => xt_rsc_7_6_i_da_d,
      qa_d => xt_rsc_7_6_i_qa_d_1,
      wea_d => xt_rsc_3_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_3_0_i_wea_d_iff
    );
  xt_rsc_7_6_i_qa <= xt_rsc_7_6_qa;
  xt_rsc_7_6_da <= xt_rsc_7_6_i_da;
  xt_rsc_7_6_adra <= xt_rsc_7_6_i_adra;
  xt_rsc_7_6_i_adra_d <= xt_rsc_0_15_i_adra_d_iff;
  xt_rsc_7_6_i_da_d <= xt_rsc_4_6_i_da_d_iff;
  xt_rsc_7_6_i_qa_d <= xt_rsc_7_6_i_qa_d_1;

  xt_rsc_7_7_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_494_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_7_7_i_qa,
      wea => xt_rsc_7_7_wea,
      da => xt_rsc_7_7_i_da,
      adra => xt_rsc_7_7_i_adra,
      adra_d => xt_rsc_7_7_i_adra_d,
      da_d => xt_rsc_7_7_i_da_d,
      qa_d => xt_rsc_7_7_i_qa_d_1,
      wea_d => xt_rsc_3_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_3_0_i_wea_d_iff
    );
  xt_rsc_7_7_i_qa <= xt_rsc_7_7_qa;
  xt_rsc_7_7_da <= xt_rsc_7_7_i_da;
  xt_rsc_7_7_adra <= xt_rsc_7_7_i_adra;
  xt_rsc_7_7_i_adra_d <= xt_rsc_0_0_i_adra_d_iff;
  xt_rsc_7_7_i_da_d <= xt_rsc_4_7_i_da_d_iff;
  xt_rsc_7_7_i_qa_d <= xt_rsc_7_7_i_qa_d_1;

  xt_rsc_7_8_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_495_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_7_8_i_qa,
      wea => xt_rsc_7_8_wea,
      da => xt_rsc_7_8_i_da,
      adra => xt_rsc_7_8_i_adra,
      adra_d => xt_rsc_7_8_i_adra_d,
      da_d => xt_rsc_7_8_i_da_d,
      qa_d => xt_rsc_7_8_i_qa_d_1,
      wea_d => xt_rsc_3_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_3_0_i_wea_d_iff
    );
  xt_rsc_7_8_i_qa <= xt_rsc_7_8_qa;
  xt_rsc_7_8_da <= xt_rsc_7_8_i_da;
  xt_rsc_7_8_adra <= xt_rsc_7_8_i_adra;
  xt_rsc_7_8_i_adra_d <= xt_rsc_0_1_i_adra_d_iff;
  xt_rsc_7_8_i_da_d <= xt_rsc_4_8_i_da_d_iff;
  xt_rsc_7_8_i_qa_d <= xt_rsc_7_8_i_qa_d_1;

  xt_rsc_7_9_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_496_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_7_9_i_qa,
      wea => xt_rsc_7_9_wea,
      da => xt_rsc_7_9_i_da,
      adra => xt_rsc_7_9_i_adra,
      adra_d => xt_rsc_7_9_i_adra_d,
      da_d => xt_rsc_7_9_i_da_d,
      qa_d => xt_rsc_7_9_i_qa_d_1,
      wea_d => xt_rsc_3_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_3_0_i_wea_d_iff
    );
  xt_rsc_7_9_i_qa <= xt_rsc_7_9_qa;
  xt_rsc_7_9_da <= xt_rsc_7_9_i_da;
  xt_rsc_7_9_adra <= xt_rsc_7_9_i_adra;
  xt_rsc_7_9_i_adra_d <= xt_rsc_4_9_i_adra_d_iff;
  xt_rsc_7_9_i_da_d <= xt_rsc_4_9_i_da_d_iff;
  xt_rsc_7_9_i_qa_d <= xt_rsc_7_9_i_qa_d_1;

  xt_rsc_7_10_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_497_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_7_10_i_qa,
      wea => xt_rsc_7_10_wea,
      da => xt_rsc_7_10_i_da,
      adra => xt_rsc_7_10_i_adra,
      adra_d => xt_rsc_7_10_i_adra_d,
      da_d => xt_rsc_7_10_i_da_d,
      qa_d => xt_rsc_7_10_i_qa_d_1,
      wea_d => xt_rsc_3_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_3_0_i_wea_d_iff
    );
  xt_rsc_7_10_i_qa <= xt_rsc_7_10_qa;
  xt_rsc_7_10_da <= xt_rsc_7_10_i_da;
  xt_rsc_7_10_adra <= xt_rsc_7_10_i_adra;
  xt_rsc_7_10_i_adra_d <= xt_rsc_4_10_i_adra_d_iff;
  xt_rsc_7_10_i_da_d <= xt_rsc_4_10_i_da_d_iff;
  xt_rsc_7_10_i_qa_d <= xt_rsc_7_10_i_qa_d_1;

  xt_rsc_7_11_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_498_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_7_11_i_qa,
      wea => xt_rsc_7_11_wea,
      da => xt_rsc_7_11_i_da,
      adra => xt_rsc_7_11_i_adra,
      adra_d => xt_rsc_7_11_i_adra_d,
      da_d => xt_rsc_7_11_i_da_d,
      qa_d => xt_rsc_7_11_i_qa_d_1,
      wea_d => xt_rsc_3_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_3_0_i_wea_d_iff
    );
  xt_rsc_7_11_i_qa <= xt_rsc_7_11_qa;
  xt_rsc_7_11_da <= xt_rsc_7_11_i_da;
  xt_rsc_7_11_adra <= xt_rsc_7_11_i_adra;
  xt_rsc_7_11_i_adra_d <= xt_rsc_0_3_i_adra_d_iff;
  xt_rsc_7_11_i_da_d <= xt_rsc_4_11_i_da_d_iff;
  xt_rsc_7_11_i_qa_d <= xt_rsc_7_11_i_qa_d_1;

  xt_rsc_7_12_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_499_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_7_12_i_qa,
      wea => xt_rsc_7_12_wea,
      da => xt_rsc_7_12_i_da,
      adra => xt_rsc_7_12_i_adra,
      adra_d => xt_rsc_7_12_i_adra_d,
      da_d => xt_rsc_7_12_i_da_d,
      qa_d => xt_rsc_7_12_i_qa_d_1,
      wea_d => xt_rsc_3_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_3_0_i_wea_d_iff
    );
  xt_rsc_7_12_i_qa <= xt_rsc_7_12_qa;
  xt_rsc_7_12_da <= xt_rsc_7_12_i_da;
  xt_rsc_7_12_adra <= xt_rsc_7_12_i_adra;
  xt_rsc_7_12_i_adra_d <= xt_rsc_0_4_i_adra_d_iff;
  xt_rsc_7_12_i_da_d <= xt_rsc_4_12_i_da_d_iff;
  xt_rsc_7_12_i_qa_d <= xt_rsc_7_12_i_qa_d_1;

  xt_rsc_7_13_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_500_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_7_13_i_qa,
      wea => xt_rsc_7_13_wea,
      da => xt_rsc_7_13_i_da,
      adra => xt_rsc_7_13_i_adra,
      adra_d => xt_rsc_7_13_i_adra_d,
      da_d => xt_rsc_7_13_i_da_d,
      qa_d => xt_rsc_7_13_i_qa_d_1,
      wea_d => xt_rsc_3_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_3_0_i_wea_d_iff
    );
  xt_rsc_7_13_i_qa <= xt_rsc_7_13_qa;
  xt_rsc_7_13_da <= xt_rsc_7_13_i_da;
  xt_rsc_7_13_adra <= xt_rsc_7_13_i_adra;
  xt_rsc_7_13_i_adra_d <= xt_rsc_0_5_i_adra_d_iff;
  xt_rsc_7_13_i_da_d <= xt_rsc_4_13_i_da_d_iff;
  xt_rsc_7_13_i_qa_d <= xt_rsc_7_13_i_qa_d_1;

  xt_rsc_7_14_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_501_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_7_14_i_qa,
      wea => xt_rsc_7_14_wea,
      da => xt_rsc_7_14_i_da,
      adra => xt_rsc_7_14_i_adra,
      adra_d => xt_rsc_7_14_i_adra_d,
      da_d => xt_rsc_7_14_i_da_d,
      qa_d => xt_rsc_7_14_i_qa_d_1,
      wea_d => xt_rsc_3_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_3_0_i_wea_d_iff
    );
  xt_rsc_7_14_i_qa <= xt_rsc_7_14_qa;
  xt_rsc_7_14_da <= xt_rsc_7_14_i_da;
  xt_rsc_7_14_adra <= xt_rsc_7_14_i_adra;
  xt_rsc_7_14_i_adra_d <= xt_rsc_0_6_i_adra_d_iff;
  xt_rsc_7_14_i_da_d <= xt_rsc_4_14_i_da_d_iff;
  xt_rsc_7_14_i_qa_d <= xt_rsc_7_14_i_qa_d_1;

  xt_rsc_7_15_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_502_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_7_15_i_qa,
      wea => xt_rsc_7_15_wea,
      da => xt_rsc_7_15_i_da,
      adra => xt_rsc_7_15_i_adra,
      adra_d => xt_rsc_7_15_i_adra_d,
      da_d => xt_rsc_7_15_i_da_d,
      qa_d => xt_rsc_7_15_i_qa_d_1,
      wea_d => xt_rsc_3_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_3_0_i_wea_d_iff
    );
  xt_rsc_7_15_i_qa <= xt_rsc_7_15_qa;
  xt_rsc_7_15_da <= xt_rsc_7_15_i_da;
  xt_rsc_7_15_adra <= xt_rsc_7_15_i_adra;
  xt_rsc_7_15_i_adra_d <= xt_rsc_0_7_i_adra_d_iff;
  xt_rsc_7_15_i_da_d <= xt_rsc_4_15_i_da_d_iff;
  xt_rsc_7_15_i_qa_d <= xt_rsc_7_15_i_qa_d_1;

  xt_rsc_7_16_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_503_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_7_16_i_qa,
      wea => xt_rsc_7_16_wea,
      da => xt_rsc_7_16_i_da,
      adra => xt_rsc_7_16_i_adra,
      adra_d => xt_rsc_7_16_i_adra_d,
      da_d => xt_rsc_7_16_i_da_d,
      qa_d => xt_rsc_7_16_i_qa_d_1,
      wea_d => xt_rsc_3_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_3_16_i_wea_d_iff
    );
  xt_rsc_7_16_i_qa <= xt_rsc_7_16_qa;
  xt_rsc_7_16_da <= xt_rsc_7_16_i_da;
  xt_rsc_7_16_adra <= xt_rsc_7_16_i_adra;
  xt_rsc_7_16_i_adra_d <= xt_rsc_0_8_i_adra_d_iff;
  xt_rsc_7_16_i_da_d <= xt_rsc_4_0_i_da_d_iff;
  xt_rsc_7_16_i_qa_d <= xt_rsc_7_16_i_qa_d_1;

  xt_rsc_7_17_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_504_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_7_17_i_qa,
      wea => xt_rsc_7_17_wea,
      da => xt_rsc_7_17_i_da,
      adra => xt_rsc_7_17_i_adra,
      adra_d => xt_rsc_7_17_i_adra_d,
      da_d => xt_rsc_7_17_i_da_d,
      qa_d => xt_rsc_7_17_i_qa_d_1,
      wea_d => xt_rsc_3_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_3_16_i_wea_d_iff
    );
  xt_rsc_7_17_i_qa <= xt_rsc_7_17_qa;
  xt_rsc_7_17_da <= xt_rsc_7_17_i_da;
  xt_rsc_7_17_adra <= xt_rsc_7_17_i_adra;
  xt_rsc_7_17_i_adra_d <= xt_rsc_4_1_i_adra_d_iff;
  xt_rsc_7_17_i_da_d <= xt_rsc_4_1_i_da_d_iff;
  xt_rsc_7_17_i_qa_d <= xt_rsc_7_17_i_qa_d_1;

  xt_rsc_7_18_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_505_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_7_18_i_qa,
      wea => xt_rsc_7_18_wea,
      da => xt_rsc_7_18_i_da,
      adra => xt_rsc_7_18_i_adra,
      adra_d => xt_rsc_7_18_i_adra_d,
      da_d => xt_rsc_7_18_i_da_d,
      qa_d => xt_rsc_7_18_i_qa_d_1,
      wea_d => xt_rsc_3_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_3_16_i_wea_d_iff
    );
  xt_rsc_7_18_i_qa <= xt_rsc_7_18_qa;
  xt_rsc_7_18_da <= xt_rsc_7_18_i_da;
  xt_rsc_7_18_adra <= xt_rsc_7_18_i_adra;
  xt_rsc_7_18_i_adra_d <= xt_rsc_4_2_i_adra_d_iff;
  xt_rsc_7_18_i_da_d <= xt_rsc_4_2_i_da_d_iff;
  xt_rsc_7_18_i_qa_d <= xt_rsc_7_18_i_qa_d_1;

  xt_rsc_7_19_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_506_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_7_19_i_qa,
      wea => xt_rsc_7_19_wea,
      da => xt_rsc_7_19_i_da,
      adra => xt_rsc_7_19_i_adra,
      adra_d => xt_rsc_7_19_i_adra_d,
      da_d => xt_rsc_7_19_i_da_d,
      qa_d => xt_rsc_7_19_i_qa_d_1,
      wea_d => xt_rsc_3_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_3_16_i_wea_d_iff
    );
  xt_rsc_7_19_i_qa <= xt_rsc_7_19_qa;
  xt_rsc_7_19_da <= xt_rsc_7_19_i_da;
  xt_rsc_7_19_adra <= xt_rsc_7_19_i_adra;
  xt_rsc_7_19_i_adra_d <= xt_rsc_0_12_i_adra_d_iff;
  xt_rsc_7_19_i_da_d <= xt_rsc_4_3_i_da_d_iff;
  xt_rsc_7_19_i_qa_d <= xt_rsc_7_19_i_qa_d_1;

  xt_rsc_7_20_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_507_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_7_20_i_qa,
      wea => xt_rsc_7_20_wea,
      da => xt_rsc_7_20_i_da,
      adra => xt_rsc_7_20_i_adra,
      adra_d => xt_rsc_7_20_i_adra_d,
      da_d => xt_rsc_7_20_i_da_d,
      qa_d => xt_rsc_7_20_i_qa_d_1,
      wea_d => xt_rsc_3_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_3_16_i_wea_d_iff
    );
  xt_rsc_7_20_i_qa <= xt_rsc_7_20_qa;
  xt_rsc_7_20_da <= xt_rsc_7_20_i_da;
  xt_rsc_7_20_adra <= xt_rsc_7_20_i_adra;
  xt_rsc_7_20_i_adra_d <= xt_rsc_0_13_i_adra_d_iff;
  xt_rsc_7_20_i_da_d <= xt_rsc_4_4_i_da_d_iff;
  xt_rsc_7_20_i_qa_d <= xt_rsc_7_20_i_qa_d_1;

  xt_rsc_7_21_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_508_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_7_21_i_qa,
      wea => xt_rsc_7_21_wea,
      da => xt_rsc_7_21_i_da,
      adra => xt_rsc_7_21_i_adra,
      adra_d => xt_rsc_7_21_i_adra_d,
      da_d => xt_rsc_7_21_i_da_d,
      qa_d => xt_rsc_7_21_i_qa_d_1,
      wea_d => xt_rsc_3_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_3_16_i_wea_d_iff
    );
  xt_rsc_7_21_i_qa <= xt_rsc_7_21_qa;
  xt_rsc_7_21_da <= xt_rsc_7_21_i_da;
  xt_rsc_7_21_adra <= xt_rsc_7_21_i_adra;
  xt_rsc_7_21_i_adra_d <= xt_rsc_0_14_i_adra_d_iff;
  xt_rsc_7_21_i_da_d <= xt_rsc_4_5_i_da_d_iff;
  xt_rsc_7_21_i_qa_d <= xt_rsc_7_21_i_qa_d_1;

  xt_rsc_7_22_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_509_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_7_22_i_qa,
      wea => xt_rsc_7_22_wea,
      da => xt_rsc_7_22_i_da,
      adra => xt_rsc_7_22_i_adra,
      adra_d => xt_rsc_7_22_i_adra_d,
      da_d => xt_rsc_7_22_i_da_d,
      qa_d => xt_rsc_7_22_i_qa_d_1,
      wea_d => xt_rsc_3_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_3_16_i_wea_d_iff
    );
  xt_rsc_7_22_i_qa <= xt_rsc_7_22_qa;
  xt_rsc_7_22_da <= xt_rsc_7_22_i_da;
  xt_rsc_7_22_adra <= xt_rsc_7_22_i_adra;
  xt_rsc_7_22_i_adra_d <= xt_rsc_0_15_i_adra_d_iff;
  xt_rsc_7_22_i_da_d <= xt_rsc_4_6_i_da_d_iff;
  xt_rsc_7_22_i_qa_d <= xt_rsc_7_22_i_qa_d_1;

  xt_rsc_7_23_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_510_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_7_23_i_qa,
      wea => xt_rsc_7_23_wea,
      da => xt_rsc_7_23_i_da,
      adra => xt_rsc_7_23_i_adra,
      adra_d => xt_rsc_7_23_i_adra_d,
      da_d => xt_rsc_7_23_i_da_d,
      qa_d => xt_rsc_7_23_i_qa_d_1,
      wea_d => xt_rsc_3_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_3_16_i_wea_d_iff
    );
  xt_rsc_7_23_i_qa <= xt_rsc_7_23_qa;
  xt_rsc_7_23_da <= xt_rsc_7_23_i_da;
  xt_rsc_7_23_adra <= xt_rsc_7_23_i_adra;
  xt_rsc_7_23_i_adra_d <= xt_rsc_0_0_i_adra_d_iff;
  xt_rsc_7_23_i_da_d <= xt_rsc_4_7_i_da_d_iff;
  xt_rsc_7_23_i_qa_d <= xt_rsc_7_23_i_qa_d_1;

  xt_rsc_7_24_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_511_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_7_24_i_qa,
      wea => xt_rsc_7_24_wea,
      da => xt_rsc_7_24_i_da,
      adra => xt_rsc_7_24_i_adra,
      adra_d => xt_rsc_7_24_i_adra_d,
      da_d => xt_rsc_7_24_i_da_d,
      qa_d => xt_rsc_7_24_i_qa_d_1,
      wea_d => xt_rsc_3_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_3_16_i_wea_d_iff
    );
  xt_rsc_7_24_i_qa <= xt_rsc_7_24_qa;
  xt_rsc_7_24_da <= xt_rsc_7_24_i_da;
  xt_rsc_7_24_adra <= xt_rsc_7_24_i_adra;
  xt_rsc_7_24_i_adra_d <= xt_rsc_0_1_i_adra_d_iff;
  xt_rsc_7_24_i_da_d <= xt_rsc_4_8_i_da_d_iff;
  xt_rsc_7_24_i_qa_d <= xt_rsc_7_24_i_qa_d_1;

  xt_rsc_7_25_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_512_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_7_25_i_qa,
      wea => xt_rsc_7_25_wea,
      da => xt_rsc_7_25_i_da,
      adra => xt_rsc_7_25_i_adra,
      adra_d => xt_rsc_7_25_i_adra_d,
      da_d => xt_rsc_7_25_i_da_d,
      qa_d => xt_rsc_7_25_i_qa_d_1,
      wea_d => xt_rsc_3_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_3_16_i_wea_d_iff
    );
  xt_rsc_7_25_i_qa <= xt_rsc_7_25_qa;
  xt_rsc_7_25_da <= xt_rsc_7_25_i_da;
  xt_rsc_7_25_adra <= xt_rsc_7_25_i_adra;
  xt_rsc_7_25_i_adra_d <= xt_rsc_4_9_i_adra_d_iff;
  xt_rsc_7_25_i_da_d <= xt_rsc_4_9_i_da_d_iff;
  xt_rsc_7_25_i_qa_d <= xt_rsc_7_25_i_qa_d_1;

  xt_rsc_7_26_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_513_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_7_26_i_qa,
      wea => xt_rsc_7_26_wea,
      da => xt_rsc_7_26_i_da,
      adra => xt_rsc_7_26_i_adra,
      adra_d => xt_rsc_7_26_i_adra_d,
      da_d => xt_rsc_7_26_i_da_d,
      qa_d => xt_rsc_7_26_i_qa_d_1,
      wea_d => xt_rsc_3_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_3_16_i_wea_d_iff
    );
  xt_rsc_7_26_i_qa <= xt_rsc_7_26_qa;
  xt_rsc_7_26_da <= xt_rsc_7_26_i_da;
  xt_rsc_7_26_adra <= xt_rsc_7_26_i_adra;
  xt_rsc_7_26_i_adra_d <= xt_rsc_4_10_i_adra_d_iff;
  xt_rsc_7_26_i_da_d <= xt_rsc_4_10_i_da_d_iff;
  xt_rsc_7_26_i_qa_d <= xt_rsc_7_26_i_qa_d_1;

  xt_rsc_7_27_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_514_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_7_27_i_qa,
      wea => xt_rsc_7_27_wea,
      da => xt_rsc_7_27_i_da,
      adra => xt_rsc_7_27_i_adra,
      adra_d => xt_rsc_7_27_i_adra_d,
      da_d => xt_rsc_7_27_i_da_d,
      qa_d => xt_rsc_7_27_i_qa_d_1,
      wea_d => xt_rsc_3_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_3_16_i_wea_d_iff
    );
  xt_rsc_7_27_i_qa <= xt_rsc_7_27_qa;
  xt_rsc_7_27_da <= xt_rsc_7_27_i_da;
  xt_rsc_7_27_adra <= xt_rsc_7_27_i_adra;
  xt_rsc_7_27_i_adra_d <= xt_rsc_0_3_i_adra_d_iff;
  xt_rsc_7_27_i_da_d <= xt_rsc_4_11_i_da_d_iff;
  xt_rsc_7_27_i_qa_d <= xt_rsc_7_27_i_qa_d_1;

  xt_rsc_7_28_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_515_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_7_28_i_qa,
      wea => xt_rsc_7_28_wea,
      da => xt_rsc_7_28_i_da,
      adra => xt_rsc_7_28_i_adra,
      adra_d => xt_rsc_7_28_i_adra_d,
      da_d => xt_rsc_7_28_i_da_d,
      qa_d => xt_rsc_7_28_i_qa_d_1,
      wea_d => xt_rsc_3_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_3_16_i_wea_d_iff
    );
  xt_rsc_7_28_i_qa <= xt_rsc_7_28_qa;
  xt_rsc_7_28_da <= xt_rsc_7_28_i_da;
  xt_rsc_7_28_adra <= xt_rsc_7_28_i_adra;
  xt_rsc_7_28_i_adra_d <= xt_rsc_0_4_i_adra_d_iff;
  xt_rsc_7_28_i_da_d <= xt_rsc_4_12_i_da_d_iff;
  xt_rsc_7_28_i_qa_d <= xt_rsc_7_28_i_qa_d_1;

  xt_rsc_7_29_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_516_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_7_29_i_qa,
      wea => xt_rsc_7_29_wea,
      da => xt_rsc_7_29_i_da,
      adra => xt_rsc_7_29_i_adra,
      adra_d => xt_rsc_7_29_i_adra_d,
      da_d => xt_rsc_7_29_i_da_d,
      qa_d => xt_rsc_7_29_i_qa_d_1,
      wea_d => xt_rsc_3_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_3_16_i_wea_d_iff
    );
  xt_rsc_7_29_i_qa <= xt_rsc_7_29_qa;
  xt_rsc_7_29_da <= xt_rsc_7_29_i_da;
  xt_rsc_7_29_adra <= xt_rsc_7_29_i_adra;
  xt_rsc_7_29_i_adra_d <= xt_rsc_0_5_i_adra_d_iff;
  xt_rsc_7_29_i_da_d <= xt_rsc_4_13_i_da_d_iff;
  xt_rsc_7_29_i_qa_d <= xt_rsc_7_29_i_qa_d_1;

  xt_rsc_7_30_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_517_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_7_30_i_qa,
      wea => xt_rsc_7_30_wea,
      da => xt_rsc_7_30_i_da,
      adra => xt_rsc_7_30_i_adra,
      adra_d => xt_rsc_7_30_i_adra_d,
      da_d => xt_rsc_7_30_i_da_d,
      qa_d => xt_rsc_7_30_i_qa_d_1,
      wea_d => xt_rsc_3_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_3_16_i_wea_d_iff
    );
  xt_rsc_7_30_i_qa <= xt_rsc_7_30_qa;
  xt_rsc_7_30_da <= xt_rsc_7_30_i_da;
  xt_rsc_7_30_adra <= xt_rsc_7_30_i_adra;
  xt_rsc_7_30_i_adra_d <= xt_rsc_0_6_i_adra_d_iff;
  xt_rsc_7_30_i_da_d <= xt_rsc_4_14_i_da_d_iff;
  xt_rsc_7_30_i_qa_d <= xt_rsc_7_30_i_qa_d_1;

  xt_rsc_7_31_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_518_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_7_31_i_qa,
      wea => xt_rsc_7_31_wea,
      da => xt_rsc_7_31_i_da,
      adra => xt_rsc_7_31_i_adra,
      adra_d => xt_rsc_7_31_i_adra_d,
      da_d => xt_rsc_7_31_i_da_d,
      qa_d => xt_rsc_7_31_i_qa_d_1,
      wea_d => xt_rsc_3_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_3_16_i_wea_d_iff
    );
  xt_rsc_7_31_i_qa <= xt_rsc_7_31_qa;
  xt_rsc_7_31_da <= xt_rsc_7_31_i_da;
  xt_rsc_7_31_adra <= xt_rsc_7_31_i_adra;
  xt_rsc_7_31_i_adra_d <= xt_rsc_0_7_i_adra_d_iff;
  xt_rsc_7_31_i_da_d <= xt_rsc_4_15_i_da_d_iff;
  xt_rsc_7_31_i_qa_d <= xt_rsc_7_31_i_qa_d_1;

  twiddle_rsc_0_0_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_519_8_32_256_256_32_1_gen
    PORT MAP(
      qb => twiddle_rsc_0_0_i_qb,
      web => twiddle_rsc_0_0_web,
      db => twiddle_rsc_0_0_i_db,
      adrb => twiddle_rsc_0_0_i_adrb,
      qa => twiddle_rsc_0_0_i_qa,
      wea => twiddle_rsc_0_0_wea,
      da => twiddle_rsc_0_0_i_da,
      adra => twiddle_rsc_0_0_i_adra,
      adra_d => twiddle_rsc_0_0_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => twiddle_rsc_0_0_i_da_d,
      qa_d => twiddle_rsc_0_0_i_qa_d_1,
      wea_d => twiddle_rsc_0_0_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => twiddle_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  twiddle_rsc_0_0_i_qb <= twiddle_rsc_0_0_qb;
  twiddle_rsc_0_0_db <= twiddle_rsc_0_0_i_db;
  twiddle_rsc_0_0_adrb <= twiddle_rsc_0_0_i_adrb;
  twiddle_rsc_0_0_i_qa <= twiddle_rsc_0_0_qa;
  twiddle_rsc_0_0_da <= twiddle_rsc_0_0_i_da;
  twiddle_rsc_0_0_adra <= twiddle_rsc_0_0_i_adra;
  twiddle_rsc_0_0_i_adra_d_1 <= STD_LOGIC_VECTOR'( "00000000") & twiddle_rsc_0_0_i_adra_d;
  twiddle_rsc_0_0_i_da_d <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
  twiddle_rsc_0_0_i_qa_d <= twiddle_rsc_0_0_i_qa_d_1;
  twiddle_rsc_0_0_i_wea_d <= STD_LOGIC_VECTOR'( "00");
  twiddle_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= twiddle_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( "00");

  twiddle_rsc_0_1_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_520_8_32_256_256_32_1_gen
    PORT MAP(
      qb => twiddle_rsc_0_1_i_qb,
      web => twiddle_rsc_0_1_web,
      db => twiddle_rsc_0_1_i_db,
      adrb => twiddle_rsc_0_1_i_adrb,
      qa => twiddle_rsc_0_1_i_qa,
      wea => twiddle_rsc_0_1_wea,
      da => twiddle_rsc_0_1_i_da,
      adra => twiddle_rsc_0_1_i_adra,
      adra_d => twiddle_rsc_0_1_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => twiddle_rsc_0_1_i_da_d,
      qa_d => twiddle_rsc_0_1_i_qa_d_1,
      wea_d => twiddle_rsc_0_1_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => twiddle_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  twiddle_rsc_0_1_i_qb <= twiddle_rsc_0_1_qb;
  twiddle_rsc_0_1_db <= twiddle_rsc_0_1_i_db;
  twiddle_rsc_0_1_adrb <= twiddle_rsc_0_1_i_adrb;
  twiddle_rsc_0_1_i_qa <= twiddle_rsc_0_1_qa;
  twiddle_rsc_0_1_da <= twiddle_rsc_0_1_i_da;
  twiddle_rsc_0_1_adra <= twiddle_rsc_0_1_i_adra;
  twiddle_rsc_0_1_i_adra_d_1 <= STD_LOGIC_VECTOR'( "00000000") & twiddle_rsc_0_1_i_adra_d;
  twiddle_rsc_0_1_i_da_d <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
  twiddle_rsc_0_1_i_qa_d <= twiddle_rsc_0_1_i_qa_d_1;
  twiddle_rsc_0_1_i_wea_d <= STD_LOGIC_VECTOR'( "00");
  twiddle_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= twiddle_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( "00");

  twiddle_rsc_0_2_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_521_8_32_256_256_32_1_gen
    PORT MAP(
      qb => twiddle_rsc_0_2_i_qb,
      web => twiddle_rsc_0_2_web,
      db => twiddle_rsc_0_2_i_db,
      adrb => twiddle_rsc_0_2_i_adrb,
      qa => twiddle_rsc_0_2_i_qa,
      wea => twiddle_rsc_0_2_wea,
      da => twiddle_rsc_0_2_i_da,
      adra => twiddle_rsc_0_2_i_adra,
      adra_d => twiddle_rsc_0_2_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => twiddle_rsc_0_2_i_da_d,
      qa_d => twiddle_rsc_0_2_i_qa_d_1,
      wea_d => twiddle_rsc_0_2_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => twiddle_rsc_0_2_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  twiddle_rsc_0_2_i_qb <= twiddle_rsc_0_2_qb;
  twiddle_rsc_0_2_db <= twiddle_rsc_0_2_i_db;
  twiddle_rsc_0_2_adrb <= twiddle_rsc_0_2_i_adrb;
  twiddle_rsc_0_2_i_qa <= twiddle_rsc_0_2_qa;
  twiddle_rsc_0_2_da <= twiddle_rsc_0_2_i_da;
  twiddle_rsc_0_2_adra <= twiddle_rsc_0_2_i_adra;
  twiddle_rsc_0_2_i_adra_d_1 <= STD_LOGIC_VECTOR'( "00000000") & twiddle_rsc_0_2_i_adra_d;
  twiddle_rsc_0_2_i_da_d <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
  twiddle_rsc_0_2_i_qa_d <= twiddle_rsc_0_2_i_qa_d_1;
  twiddle_rsc_0_2_i_wea_d <= STD_LOGIC_VECTOR'( "00");
  twiddle_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= twiddle_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_rsc_0_2_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( "00");

  twiddle_rsc_0_3_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_522_8_32_256_256_32_1_gen
    PORT MAP(
      qb => twiddle_rsc_0_3_i_qb,
      web => twiddle_rsc_0_3_web,
      db => twiddle_rsc_0_3_i_db,
      adrb => twiddle_rsc_0_3_i_adrb,
      qa => twiddle_rsc_0_3_i_qa,
      wea => twiddle_rsc_0_3_wea,
      da => twiddle_rsc_0_3_i_da,
      adra => twiddle_rsc_0_3_i_adra,
      adra_d => twiddle_rsc_0_3_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => twiddle_rsc_0_3_i_da_d,
      qa_d => twiddle_rsc_0_3_i_qa_d_1,
      wea_d => twiddle_rsc_0_3_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => twiddle_rsc_0_3_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  twiddle_rsc_0_3_i_qb <= twiddle_rsc_0_3_qb;
  twiddle_rsc_0_3_db <= twiddle_rsc_0_3_i_db;
  twiddle_rsc_0_3_adrb <= twiddle_rsc_0_3_i_adrb;
  twiddle_rsc_0_3_i_qa <= twiddle_rsc_0_3_qa;
  twiddle_rsc_0_3_da <= twiddle_rsc_0_3_i_da;
  twiddle_rsc_0_3_adra <= twiddle_rsc_0_3_i_adra;
  twiddle_rsc_0_3_i_adra_d_1 <= STD_LOGIC_VECTOR'( "00000000") & twiddle_rsc_0_3_i_adra_d;
  twiddle_rsc_0_3_i_da_d <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
  twiddle_rsc_0_3_i_qa_d <= twiddle_rsc_0_3_i_qa_d_1;
  twiddle_rsc_0_3_i_wea_d <= STD_LOGIC_VECTOR'( "00");
  twiddle_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= twiddle_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_rsc_0_3_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( "00");

  twiddle_rsc_0_4_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_523_8_32_256_256_32_1_gen
    PORT MAP(
      qb => twiddle_rsc_0_4_i_qb,
      web => twiddle_rsc_0_4_web,
      db => twiddle_rsc_0_4_i_db,
      adrb => twiddle_rsc_0_4_i_adrb,
      qa => twiddle_rsc_0_4_i_qa,
      wea => twiddle_rsc_0_4_wea,
      da => twiddle_rsc_0_4_i_da,
      adra => twiddle_rsc_0_4_i_adra,
      adra_d => twiddle_rsc_0_4_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => twiddle_rsc_0_4_i_da_d,
      qa_d => twiddle_rsc_0_4_i_qa_d_1,
      wea_d => twiddle_rsc_0_4_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => twiddle_rsc_0_4_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  twiddle_rsc_0_4_i_qb <= twiddle_rsc_0_4_qb;
  twiddle_rsc_0_4_db <= twiddle_rsc_0_4_i_db;
  twiddle_rsc_0_4_adrb <= twiddle_rsc_0_4_i_adrb;
  twiddle_rsc_0_4_i_qa <= twiddle_rsc_0_4_qa;
  twiddle_rsc_0_4_da <= twiddle_rsc_0_4_i_da;
  twiddle_rsc_0_4_adra <= twiddle_rsc_0_4_i_adra;
  twiddle_rsc_0_4_i_adra_d_1 <= STD_LOGIC_VECTOR'( "00000000") & twiddle_rsc_0_4_i_adra_d;
  twiddle_rsc_0_4_i_da_d <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
  twiddle_rsc_0_4_i_qa_d <= twiddle_rsc_0_4_i_qa_d_1;
  twiddle_rsc_0_4_i_wea_d <= STD_LOGIC_VECTOR'( "00");
  twiddle_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= twiddle_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_rsc_0_4_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( "00");

  twiddle_rsc_0_5_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_524_8_32_256_256_32_1_gen
    PORT MAP(
      qb => twiddle_rsc_0_5_i_qb,
      web => twiddle_rsc_0_5_web,
      db => twiddle_rsc_0_5_i_db,
      adrb => twiddle_rsc_0_5_i_adrb,
      qa => twiddle_rsc_0_5_i_qa,
      wea => twiddle_rsc_0_5_wea,
      da => twiddle_rsc_0_5_i_da,
      adra => twiddle_rsc_0_5_i_adra,
      adra_d => twiddle_rsc_0_5_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => twiddle_rsc_0_5_i_da_d,
      qa_d => twiddle_rsc_0_5_i_qa_d_1,
      wea_d => twiddle_rsc_0_5_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => twiddle_rsc_0_5_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  twiddle_rsc_0_5_i_qb <= twiddle_rsc_0_5_qb;
  twiddle_rsc_0_5_db <= twiddle_rsc_0_5_i_db;
  twiddle_rsc_0_5_adrb <= twiddle_rsc_0_5_i_adrb;
  twiddle_rsc_0_5_i_qa <= twiddle_rsc_0_5_qa;
  twiddle_rsc_0_5_da <= twiddle_rsc_0_5_i_da;
  twiddle_rsc_0_5_adra <= twiddle_rsc_0_5_i_adra;
  twiddle_rsc_0_5_i_adra_d_1 <= STD_LOGIC_VECTOR'( "00000000") & twiddle_rsc_0_5_i_adra_d;
  twiddle_rsc_0_5_i_da_d <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
  twiddle_rsc_0_5_i_qa_d <= twiddle_rsc_0_5_i_qa_d_1;
  twiddle_rsc_0_5_i_wea_d <= STD_LOGIC_VECTOR'( "00");
  twiddle_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= twiddle_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_rsc_0_5_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( "00");

  twiddle_rsc_0_6_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_525_8_32_256_256_32_1_gen
    PORT MAP(
      qb => twiddle_rsc_0_6_i_qb,
      web => twiddle_rsc_0_6_web,
      db => twiddle_rsc_0_6_i_db,
      adrb => twiddle_rsc_0_6_i_adrb,
      qa => twiddle_rsc_0_6_i_qa,
      wea => twiddle_rsc_0_6_wea,
      da => twiddle_rsc_0_6_i_da,
      adra => twiddle_rsc_0_6_i_adra,
      adra_d => twiddle_rsc_0_6_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => twiddle_rsc_0_6_i_da_d,
      qa_d => twiddle_rsc_0_6_i_qa_d_1,
      wea_d => twiddle_rsc_0_6_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => twiddle_rsc_0_6_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  twiddle_rsc_0_6_i_qb <= twiddle_rsc_0_6_qb;
  twiddle_rsc_0_6_db <= twiddle_rsc_0_6_i_db;
  twiddle_rsc_0_6_adrb <= twiddle_rsc_0_6_i_adrb;
  twiddle_rsc_0_6_i_qa <= twiddle_rsc_0_6_qa;
  twiddle_rsc_0_6_da <= twiddle_rsc_0_6_i_da;
  twiddle_rsc_0_6_adra <= twiddle_rsc_0_6_i_adra;
  twiddle_rsc_0_6_i_adra_d_1 <= STD_LOGIC_VECTOR'( "00000000") & twiddle_rsc_0_6_i_adra_d;
  twiddle_rsc_0_6_i_da_d <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
  twiddle_rsc_0_6_i_qa_d <= twiddle_rsc_0_6_i_qa_d_1;
  twiddle_rsc_0_6_i_wea_d <= STD_LOGIC_VECTOR'( "00");
  twiddle_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= twiddle_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_rsc_0_6_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( "00");

  twiddle_rsc_0_7_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_526_8_32_256_256_32_1_gen
    PORT MAP(
      qb => twiddle_rsc_0_7_i_qb,
      web => twiddle_rsc_0_7_web,
      db => twiddle_rsc_0_7_i_db,
      adrb => twiddle_rsc_0_7_i_adrb,
      qa => twiddle_rsc_0_7_i_qa,
      wea => twiddle_rsc_0_7_wea,
      da => twiddle_rsc_0_7_i_da,
      adra => twiddle_rsc_0_7_i_adra,
      adra_d => twiddle_rsc_0_7_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => twiddle_rsc_0_7_i_da_d,
      qa_d => twiddle_rsc_0_7_i_qa_d_1,
      wea_d => twiddle_rsc_0_7_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => twiddle_rsc_0_7_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  twiddle_rsc_0_7_i_qb <= twiddle_rsc_0_7_qb;
  twiddle_rsc_0_7_db <= twiddle_rsc_0_7_i_db;
  twiddle_rsc_0_7_adrb <= twiddle_rsc_0_7_i_adrb;
  twiddle_rsc_0_7_i_qa <= twiddle_rsc_0_7_qa;
  twiddle_rsc_0_7_da <= twiddle_rsc_0_7_i_da;
  twiddle_rsc_0_7_adra <= twiddle_rsc_0_7_i_adra;
  twiddle_rsc_0_7_i_adra_d_1 <= STD_LOGIC_VECTOR'( "00000000") & twiddle_rsc_0_7_i_adra_d;
  twiddle_rsc_0_7_i_da_d <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
  twiddle_rsc_0_7_i_qa_d <= twiddle_rsc_0_7_i_qa_d_1;
  twiddle_rsc_0_7_i_wea_d <= STD_LOGIC_VECTOR'( "00");
  twiddle_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= twiddle_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_rsc_0_7_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( "00");

  twiddle_rsc_0_8_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_527_8_32_256_256_32_1_gen
    PORT MAP(
      qb => twiddle_rsc_0_8_i_qb,
      web => twiddle_rsc_0_8_web,
      db => twiddle_rsc_0_8_i_db,
      adrb => twiddle_rsc_0_8_i_adrb,
      qa => twiddle_rsc_0_8_i_qa,
      wea => twiddle_rsc_0_8_wea,
      da => twiddle_rsc_0_8_i_da,
      adra => twiddle_rsc_0_8_i_adra,
      adra_d => twiddle_rsc_0_8_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => twiddle_rsc_0_8_i_da_d,
      qa_d => twiddle_rsc_0_8_i_qa_d_1,
      wea_d => twiddle_rsc_0_8_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => twiddle_rsc_0_8_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  twiddle_rsc_0_8_i_qb <= twiddle_rsc_0_8_qb;
  twiddle_rsc_0_8_db <= twiddle_rsc_0_8_i_db;
  twiddle_rsc_0_8_adrb <= twiddle_rsc_0_8_i_adrb;
  twiddle_rsc_0_8_i_qa <= twiddle_rsc_0_8_qa;
  twiddle_rsc_0_8_da <= twiddle_rsc_0_8_i_da;
  twiddle_rsc_0_8_adra <= twiddle_rsc_0_8_i_adra;
  twiddle_rsc_0_8_i_adra_d_1 <= STD_LOGIC_VECTOR'( "00000000") & twiddle_rsc_0_8_i_adra_d;
  twiddle_rsc_0_8_i_da_d <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
  twiddle_rsc_0_8_i_qa_d <= twiddle_rsc_0_8_i_qa_d_1;
  twiddle_rsc_0_8_i_wea_d <= STD_LOGIC_VECTOR'( "00");
  twiddle_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= twiddle_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_rsc_0_8_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( "00");

  twiddle_rsc_0_9_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_528_8_32_256_256_32_1_gen
    PORT MAP(
      qb => twiddle_rsc_0_9_i_qb,
      web => twiddle_rsc_0_9_web,
      db => twiddle_rsc_0_9_i_db,
      adrb => twiddle_rsc_0_9_i_adrb,
      qa => twiddle_rsc_0_9_i_qa,
      wea => twiddle_rsc_0_9_wea,
      da => twiddle_rsc_0_9_i_da,
      adra => twiddle_rsc_0_9_i_adra,
      adra_d => twiddle_rsc_0_9_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => twiddle_rsc_0_9_i_da_d,
      qa_d => twiddle_rsc_0_9_i_qa_d_1,
      wea_d => twiddle_rsc_0_9_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => twiddle_rsc_0_9_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  twiddle_rsc_0_9_i_qb <= twiddle_rsc_0_9_qb;
  twiddle_rsc_0_9_db <= twiddle_rsc_0_9_i_db;
  twiddle_rsc_0_9_adrb <= twiddle_rsc_0_9_i_adrb;
  twiddle_rsc_0_9_i_qa <= twiddle_rsc_0_9_qa;
  twiddle_rsc_0_9_da <= twiddle_rsc_0_9_i_da;
  twiddle_rsc_0_9_adra <= twiddle_rsc_0_9_i_adra;
  twiddle_rsc_0_9_i_adra_d_1 <= STD_LOGIC_VECTOR'( "00000000") & twiddle_rsc_0_9_i_adra_d;
  twiddle_rsc_0_9_i_da_d <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
  twiddle_rsc_0_9_i_qa_d <= twiddle_rsc_0_9_i_qa_d_1;
  twiddle_rsc_0_9_i_wea_d <= STD_LOGIC_VECTOR'( "00");
  twiddle_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= twiddle_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_rsc_0_9_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( "00");

  twiddle_rsc_0_10_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_529_8_32_256_256_32_1_gen
    PORT MAP(
      qb => twiddle_rsc_0_10_i_qb,
      web => twiddle_rsc_0_10_web,
      db => twiddle_rsc_0_10_i_db,
      adrb => twiddle_rsc_0_10_i_adrb,
      qa => twiddle_rsc_0_10_i_qa,
      wea => twiddle_rsc_0_10_wea,
      da => twiddle_rsc_0_10_i_da,
      adra => twiddle_rsc_0_10_i_adra,
      adra_d => twiddle_rsc_0_10_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => twiddle_rsc_0_10_i_da_d,
      qa_d => twiddle_rsc_0_10_i_qa_d_1,
      wea_d => twiddle_rsc_0_10_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => twiddle_rsc_0_10_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  twiddle_rsc_0_10_i_qb <= twiddle_rsc_0_10_qb;
  twiddle_rsc_0_10_db <= twiddle_rsc_0_10_i_db;
  twiddle_rsc_0_10_adrb <= twiddle_rsc_0_10_i_adrb;
  twiddle_rsc_0_10_i_qa <= twiddle_rsc_0_10_qa;
  twiddle_rsc_0_10_da <= twiddle_rsc_0_10_i_da;
  twiddle_rsc_0_10_adra <= twiddle_rsc_0_10_i_adra;
  twiddle_rsc_0_10_i_adra_d_1 <= STD_LOGIC_VECTOR'( "00000000") & twiddle_rsc_0_10_i_adra_d;
  twiddle_rsc_0_10_i_da_d <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
  twiddle_rsc_0_10_i_qa_d <= twiddle_rsc_0_10_i_qa_d_1;
  twiddle_rsc_0_10_i_wea_d <= STD_LOGIC_VECTOR'( "00");
  twiddle_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= twiddle_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_rsc_0_10_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( "00");

  twiddle_rsc_0_11_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_530_8_32_256_256_32_1_gen
    PORT MAP(
      qb => twiddle_rsc_0_11_i_qb,
      web => twiddle_rsc_0_11_web,
      db => twiddle_rsc_0_11_i_db,
      adrb => twiddle_rsc_0_11_i_adrb,
      qa => twiddle_rsc_0_11_i_qa,
      wea => twiddle_rsc_0_11_wea,
      da => twiddle_rsc_0_11_i_da,
      adra => twiddle_rsc_0_11_i_adra,
      adra_d => twiddle_rsc_0_11_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => twiddle_rsc_0_11_i_da_d,
      qa_d => twiddle_rsc_0_11_i_qa_d_1,
      wea_d => twiddle_rsc_0_11_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => twiddle_rsc_0_11_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  twiddle_rsc_0_11_i_qb <= twiddle_rsc_0_11_qb;
  twiddle_rsc_0_11_db <= twiddle_rsc_0_11_i_db;
  twiddle_rsc_0_11_adrb <= twiddle_rsc_0_11_i_adrb;
  twiddle_rsc_0_11_i_qa <= twiddle_rsc_0_11_qa;
  twiddle_rsc_0_11_da <= twiddle_rsc_0_11_i_da;
  twiddle_rsc_0_11_adra <= twiddle_rsc_0_11_i_adra;
  twiddle_rsc_0_11_i_adra_d_1 <= STD_LOGIC_VECTOR'( "00000000") & twiddle_rsc_0_11_i_adra_d;
  twiddle_rsc_0_11_i_da_d <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
  twiddle_rsc_0_11_i_qa_d <= twiddle_rsc_0_11_i_qa_d_1;
  twiddle_rsc_0_11_i_wea_d <= STD_LOGIC_VECTOR'( "00");
  twiddle_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= twiddle_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_rsc_0_11_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( "00");

  twiddle_rsc_0_12_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_531_8_32_256_256_32_1_gen
    PORT MAP(
      qb => twiddle_rsc_0_12_i_qb,
      web => twiddle_rsc_0_12_web,
      db => twiddle_rsc_0_12_i_db,
      adrb => twiddle_rsc_0_12_i_adrb,
      qa => twiddle_rsc_0_12_i_qa,
      wea => twiddle_rsc_0_12_wea,
      da => twiddle_rsc_0_12_i_da,
      adra => twiddle_rsc_0_12_i_adra,
      adra_d => twiddle_rsc_0_12_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => twiddle_rsc_0_12_i_da_d,
      qa_d => twiddle_rsc_0_12_i_qa_d_1,
      wea_d => twiddle_rsc_0_12_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => twiddle_rsc_0_12_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  twiddle_rsc_0_12_i_qb <= twiddle_rsc_0_12_qb;
  twiddle_rsc_0_12_db <= twiddle_rsc_0_12_i_db;
  twiddle_rsc_0_12_adrb <= twiddle_rsc_0_12_i_adrb;
  twiddle_rsc_0_12_i_qa <= twiddle_rsc_0_12_qa;
  twiddle_rsc_0_12_da <= twiddle_rsc_0_12_i_da;
  twiddle_rsc_0_12_adra <= twiddle_rsc_0_12_i_adra;
  twiddle_rsc_0_12_i_adra_d_1 <= STD_LOGIC_VECTOR'( "00000000") & twiddle_rsc_0_12_i_adra_d;
  twiddle_rsc_0_12_i_da_d <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
  twiddle_rsc_0_12_i_qa_d <= twiddle_rsc_0_12_i_qa_d_1;
  twiddle_rsc_0_12_i_wea_d <= STD_LOGIC_VECTOR'( "00");
  twiddle_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= twiddle_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_rsc_0_12_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( "00");

  twiddle_rsc_0_13_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_532_8_32_256_256_32_1_gen
    PORT MAP(
      qb => twiddle_rsc_0_13_i_qb,
      web => twiddle_rsc_0_13_web,
      db => twiddle_rsc_0_13_i_db,
      adrb => twiddle_rsc_0_13_i_adrb,
      qa => twiddle_rsc_0_13_i_qa,
      wea => twiddle_rsc_0_13_wea,
      da => twiddle_rsc_0_13_i_da,
      adra => twiddle_rsc_0_13_i_adra,
      adra_d => twiddle_rsc_0_13_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => twiddle_rsc_0_13_i_da_d,
      qa_d => twiddle_rsc_0_13_i_qa_d_1,
      wea_d => twiddle_rsc_0_13_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => twiddle_rsc_0_13_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  twiddle_rsc_0_13_i_qb <= twiddle_rsc_0_13_qb;
  twiddle_rsc_0_13_db <= twiddle_rsc_0_13_i_db;
  twiddle_rsc_0_13_adrb <= twiddle_rsc_0_13_i_adrb;
  twiddle_rsc_0_13_i_qa <= twiddle_rsc_0_13_qa;
  twiddle_rsc_0_13_da <= twiddle_rsc_0_13_i_da;
  twiddle_rsc_0_13_adra <= twiddle_rsc_0_13_i_adra;
  twiddle_rsc_0_13_i_adra_d_1 <= STD_LOGIC_VECTOR'( "00000000") & twiddle_rsc_0_13_i_adra_d;
  twiddle_rsc_0_13_i_da_d <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
  twiddle_rsc_0_13_i_qa_d <= twiddle_rsc_0_13_i_qa_d_1;
  twiddle_rsc_0_13_i_wea_d <= STD_LOGIC_VECTOR'( "00");
  twiddle_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= twiddle_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_rsc_0_13_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( "00");

  twiddle_rsc_0_14_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_533_8_32_256_256_32_1_gen
    PORT MAP(
      qb => twiddle_rsc_0_14_i_qb,
      web => twiddle_rsc_0_14_web,
      db => twiddle_rsc_0_14_i_db,
      adrb => twiddle_rsc_0_14_i_adrb,
      qa => twiddle_rsc_0_14_i_qa,
      wea => twiddle_rsc_0_14_wea,
      da => twiddle_rsc_0_14_i_da,
      adra => twiddle_rsc_0_14_i_adra,
      adra_d => twiddle_rsc_0_14_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => twiddle_rsc_0_14_i_da_d,
      qa_d => twiddle_rsc_0_14_i_qa_d_1,
      wea_d => twiddle_rsc_0_14_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => twiddle_rsc_0_14_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  twiddle_rsc_0_14_i_qb <= twiddle_rsc_0_14_qb;
  twiddle_rsc_0_14_db <= twiddle_rsc_0_14_i_db;
  twiddle_rsc_0_14_adrb <= twiddle_rsc_0_14_i_adrb;
  twiddle_rsc_0_14_i_qa <= twiddle_rsc_0_14_qa;
  twiddle_rsc_0_14_da <= twiddle_rsc_0_14_i_da;
  twiddle_rsc_0_14_adra <= twiddle_rsc_0_14_i_adra;
  twiddle_rsc_0_14_i_adra_d_1 <= STD_LOGIC_VECTOR'( "00000000") & twiddle_rsc_0_14_i_adra_d;
  twiddle_rsc_0_14_i_da_d <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
  twiddle_rsc_0_14_i_qa_d <= twiddle_rsc_0_14_i_qa_d_1;
  twiddle_rsc_0_14_i_wea_d <= STD_LOGIC_VECTOR'( "00");
  twiddle_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= twiddle_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_rsc_0_14_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( "00");

  twiddle_rsc_0_15_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_534_8_32_256_256_32_1_gen
    PORT MAP(
      qb => twiddle_rsc_0_15_i_qb,
      web => twiddle_rsc_0_15_web,
      db => twiddle_rsc_0_15_i_db,
      adrb => twiddle_rsc_0_15_i_adrb,
      qa => twiddle_rsc_0_15_i_qa,
      wea => twiddle_rsc_0_15_wea,
      da => twiddle_rsc_0_15_i_da,
      adra => twiddle_rsc_0_15_i_adra,
      adra_d => twiddle_rsc_0_15_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => twiddle_rsc_0_15_i_da_d,
      qa_d => twiddle_rsc_0_15_i_qa_d_1,
      wea_d => twiddle_rsc_0_15_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => twiddle_rsc_0_15_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  twiddle_rsc_0_15_i_qb <= twiddle_rsc_0_15_qb;
  twiddle_rsc_0_15_db <= twiddle_rsc_0_15_i_db;
  twiddle_rsc_0_15_adrb <= twiddle_rsc_0_15_i_adrb;
  twiddle_rsc_0_15_i_qa <= twiddle_rsc_0_15_qa;
  twiddle_rsc_0_15_da <= twiddle_rsc_0_15_i_da;
  twiddle_rsc_0_15_adra <= twiddle_rsc_0_15_i_adra;
  twiddle_rsc_0_15_i_adra_d_1 <= STD_LOGIC_VECTOR'( "00000000") & twiddle_rsc_0_15_i_adra_d;
  twiddle_rsc_0_15_i_da_d <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
  twiddle_rsc_0_15_i_qa_d <= twiddle_rsc_0_15_i_qa_d_1;
  twiddle_rsc_0_15_i_wea_d <= STD_LOGIC_VECTOR'( "00");
  twiddle_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= twiddle_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_rsc_0_15_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( "00");

  twiddle_h_rsc_0_0_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_535_8_32_256_256_32_1_gen
    PORT MAP(
      qb => twiddle_h_rsc_0_0_i_qb,
      web => twiddle_h_rsc_0_0_web,
      db => twiddle_h_rsc_0_0_i_db,
      adrb => twiddle_h_rsc_0_0_i_adrb,
      qa => twiddle_h_rsc_0_0_i_qa,
      wea => twiddle_h_rsc_0_0_wea,
      da => twiddle_h_rsc_0_0_i_da,
      adra => twiddle_h_rsc_0_0_i_adra,
      adra_d => twiddle_h_rsc_0_0_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => twiddle_h_rsc_0_0_i_da_d,
      qa_d => twiddle_h_rsc_0_0_i_qa_d_1,
      wea_d => twiddle_h_rsc_0_0_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => twiddle_h_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  twiddle_h_rsc_0_0_i_qb <= twiddle_h_rsc_0_0_qb;
  twiddle_h_rsc_0_0_db <= twiddle_h_rsc_0_0_i_db;
  twiddle_h_rsc_0_0_adrb <= twiddle_h_rsc_0_0_i_adrb;
  twiddle_h_rsc_0_0_i_qa <= twiddle_h_rsc_0_0_qa;
  twiddle_h_rsc_0_0_da <= twiddle_h_rsc_0_0_i_da;
  twiddle_h_rsc_0_0_adra <= twiddle_h_rsc_0_0_i_adra;
  twiddle_h_rsc_0_0_i_adra_d_1 <= STD_LOGIC_VECTOR'( "00000000") & twiddle_h_rsc_0_0_i_adra_d;
  twiddle_h_rsc_0_0_i_da_d <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
  twiddle_h_rsc_0_0_i_qa_d <= twiddle_h_rsc_0_0_i_qa_d_1;
  twiddle_h_rsc_0_0_i_wea_d <= STD_LOGIC_VECTOR'( "00");
  twiddle_h_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= twiddle_h_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_h_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( "00");

  twiddle_h_rsc_0_1_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_536_8_32_256_256_32_1_gen
    PORT MAP(
      qb => twiddle_h_rsc_0_1_i_qb,
      web => twiddle_h_rsc_0_1_web,
      db => twiddle_h_rsc_0_1_i_db,
      adrb => twiddle_h_rsc_0_1_i_adrb,
      qa => twiddle_h_rsc_0_1_i_qa,
      wea => twiddle_h_rsc_0_1_wea,
      da => twiddle_h_rsc_0_1_i_da,
      adra => twiddle_h_rsc_0_1_i_adra,
      adra_d => twiddle_h_rsc_0_1_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => twiddle_h_rsc_0_1_i_da_d,
      qa_d => twiddle_h_rsc_0_1_i_qa_d_1,
      wea_d => twiddle_h_rsc_0_1_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => twiddle_h_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  twiddle_h_rsc_0_1_i_qb <= twiddle_h_rsc_0_1_qb;
  twiddle_h_rsc_0_1_db <= twiddle_h_rsc_0_1_i_db;
  twiddle_h_rsc_0_1_adrb <= twiddle_h_rsc_0_1_i_adrb;
  twiddle_h_rsc_0_1_i_qa <= twiddle_h_rsc_0_1_qa;
  twiddle_h_rsc_0_1_da <= twiddle_h_rsc_0_1_i_da;
  twiddle_h_rsc_0_1_adra <= twiddle_h_rsc_0_1_i_adra;
  twiddle_h_rsc_0_1_i_adra_d_1 <= STD_LOGIC_VECTOR'( "00000000") & twiddle_h_rsc_0_1_i_adra_d;
  twiddle_h_rsc_0_1_i_da_d <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
  twiddle_h_rsc_0_1_i_qa_d <= twiddle_h_rsc_0_1_i_qa_d_1;
  twiddle_h_rsc_0_1_i_wea_d <= STD_LOGIC_VECTOR'( "00");
  twiddle_h_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= twiddle_h_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_h_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( "00");

  twiddle_h_rsc_0_2_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_537_8_32_256_256_32_1_gen
    PORT MAP(
      qb => twiddle_h_rsc_0_2_i_qb,
      web => twiddle_h_rsc_0_2_web,
      db => twiddle_h_rsc_0_2_i_db,
      adrb => twiddle_h_rsc_0_2_i_adrb,
      qa => twiddle_h_rsc_0_2_i_qa,
      wea => twiddle_h_rsc_0_2_wea,
      da => twiddle_h_rsc_0_2_i_da,
      adra => twiddle_h_rsc_0_2_i_adra,
      adra_d => twiddle_h_rsc_0_2_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => twiddle_h_rsc_0_2_i_da_d,
      qa_d => twiddle_h_rsc_0_2_i_qa_d_1,
      wea_d => twiddle_h_rsc_0_2_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => twiddle_h_rsc_0_2_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  twiddle_h_rsc_0_2_i_qb <= twiddle_h_rsc_0_2_qb;
  twiddle_h_rsc_0_2_db <= twiddle_h_rsc_0_2_i_db;
  twiddle_h_rsc_0_2_adrb <= twiddle_h_rsc_0_2_i_adrb;
  twiddle_h_rsc_0_2_i_qa <= twiddle_h_rsc_0_2_qa;
  twiddle_h_rsc_0_2_da <= twiddle_h_rsc_0_2_i_da;
  twiddle_h_rsc_0_2_adra <= twiddle_h_rsc_0_2_i_adra;
  twiddle_h_rsc_0_2_i_adra_d_1 <= STD_LOGIC_VECTOR'( "00000000") & twiddle_h_rsc_0_2_i_adra_d;
  twiddle_h_rsc_0_2_i_da_d <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
  twiddle_h_rsc_0_2_i_qa_d <= twiddle_h_rsc_0_2_i_qa_d_1;
  twiddle_h_rsc_0_2_i_wea_d <= STD_LOGIC_VECTOR'( "00");
  twiddle_h_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= twiddle_h_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_h_rsc_0_2_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( "00");

  twiddle_h_rsc_0_3_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_538_8_32_256_256_32_1_gen
    PORT MAP(
      qb => twiddle_h_rsc_0_3_i_qb,
      web => twiddle_h_rsc_0_3_web,
      db => twiddle_h_rsc_0_3_i_db,
      adrb => twiddle_h_rsc_0_3_i_adrb,
      qa => twiddle_h_rsc_0_3_i_qa,
      wea => twiddle_h_rsc_0_3_wea,
      da => twiddle_h_rsc_0_3_i_da,
      adra => twiddle_h_rsc_0_3_i_adra,
      adra_d => twiddle_h_rsc_0_3_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => twiddle_h_rsc_0_3_i_da_d,
      qa_d => twiddle_h_rsc_0_3_i_qa_d_1,
      wea_d => twiddle_h_rsc_0_3_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => twiddle_h_rsc_0_3_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  twiddle_h_rsc_0_3_i_qb <= twiddle_h_rsc_0_3_qb;
  twiddle_h_rsc_0_3_db <= twiddle_h_rsc_0_3_i_db;
  twiddle_h_rsc_0_3_adrb <= twiddle_h_rsc_0_3_i_adrb;
  twiddle_h_rsc_0_3_i_qa <= twiddle_h_rsc_0_3_qa;
  twiddle_h_rsc_0_3_da <= twiddle_h_rsc_0_3_i_da;
  twiddle_h_rsc_0_3_adra <= twiddle_h_rsc_0_3_i_adra;
  twiddle_h_rsc_0_3_i_adra_d_1 <= STD_LOGIC_VECTOR'( "00000000") & twiddle_h_rsc_0_3_i_adra_d;
  twiddle_h_rsc_0_3_i_da_d <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
  twiddle_h_rsc_0_3_i_qa_d <= twiddle_h_rsc_0_3_i_qa_d_1;
  twiddle_h_rsc_0_3_i_wea_d <= STD_LOGIC_VECTOR'( "00");
  twiddle_h_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= twiddle_h_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_h_rsc_0_3_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( "00");

  twiddle_h_rsc_0_4_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_539_8_32_256_256_32_1_gen
    PORT MAP(
      qb => twiddle_h_rsc_0_4_i_qb,
      web => twiddle_h_rsc_0_4_web,
      db => twiddle_h_rsc_0_4_i_db,
      adrb => twiddle_h_rsc_0_4_i_adrb,
      qa => twiddle_h_rsc_0_4_i_qa,
      wea => twiddle_h_rsc_0_4_wea,
      da => twiddle_h_rsc_0_4_i_da,
      adra => twiddle_h_rsc_0_4_i_adra,
      adra_d => twiddle_h_rsc_0_4_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => twiddle_h_rsc_0_4_i_da_d,
      qa_d => twiddle_h_rsc_0_4_i_qa_d_1,
      wea_d => twiddle_h_rsc_0_4_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => twiddle_h_rsc_0_4_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  twiddle_h_rsc_0_4_i_qb <= twiddle_h_rsc_0_4_qb;
  twiddle_h_rsc_0_4_db <= twiddle_h_rsc_0_4_i_db;
  twiddle_h_rsc_0_4_adrb <= twiddle_h_rsc_0_4_i_adrb;
  twiddle_h_rsc_0_4_i_qa <= twiddle_h_rsc_0_4_qa;
  twiddle_h_rsc_0_4_da <= twiddle_h_rsc_0_4_i_da;
  twiddle_h_rsc_0_4_adra <= twiddle_h_rsc_0_4_i_adra;
  twiddle_h_rsc_0_4_i_adra_d_1 <= STD_LOGIC_VECTOR'( "00000000") & twiddle_h_rsc_0_4_i_adra_d;
  twiddle_h_rsc_0_4_i_da_d <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
  twiddle_h_rsc_0_4_i_qa_d <= twiddle_h_rsc_0_4_i_qa_d_1;
  twiddle_h_rsc_0_4_i_wea_d <= STD_LOGIC_VECTOR'( "00");
  twiddle_h_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= twiddle_h_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_h_rsc_0_4_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( "00");

  twiddle_h_rsc_0_5_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_540_8_32_256_256_32_1_gen
    PORT MAP(
      qb => twiddle_h_rsc_0_5_i_qb,
      web => twiddle_h_rsc_0_5_web,
      db => twiddle_h_rsc_0_5_i_db,
      adrb => twiddle_h_rsc_0_5_i_adrb,
      qa => twiddle_h_rsc_0_5_i_qa,
      wea => twiddle_h_rsc_0_5_wea,
      da => twiddle_h_rsc_0_5_i_da,
      adra => twiddle_h_rsc_0_5_i_adra,
      adra_d => twiddle_h_rsc_0_5_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => twiddle_h_rsc_0_5_i_da_d,
      qa_d => twiddle_h_rsc_0_5_i_qa_d_1,
      wea_d => twiddle_h_rsc_0_5_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => twiddle_h_rsc_0_5_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  twiddle_h_rsc_0_5_i_qb <= twiddle_h_rsc_0_5_qb;
  twiddle_h_rsc_0_5_db <= twiddle_h_rsc_0_5_i_db;
  twiddle_h_rsc_0_5_adrb <= twiddle_h_rsc_0_5_i_adrb;
  twiddle_h_rsc_0_5_i_qa <= twiddle_h_rsc_0_5_qa;
  twiddle_h_rsc_0_5_da <= twiddle_h_rsc_0_5_i_da;
  twiddle_h_rsc_0_5_adra <= twiddle_h_rsc_0_5_i_adra;
  twiddle_h_rsc_0_5_i_adra_d_1 <= STD_LOGIC_VECTOR'( "00000000") & twiddle_h_rsc_0_5_i_adra_d;
  twiddle_h_rsc_0_5_i_da_d <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
  twiddle_h_rsc_0_5_i_qa_d <= twiddle_h_rsc_0_5_i_qa_d_1;
  twiddle_h_rsc_0_5_i_wea_d <= STD_LOGIC_VECTOR'( "00");
  twiddle_h_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= twiddle_h_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_h_rsc_0_5_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( "00");

  twiddle_h_rsc_0_6_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_541_8_32_256_256_32_1_gen
    PORT MAP(
      qb => twiddle_h_rsc_0_6_i_qb,
      web => twiddle_h_rsc_0_6_web,
      db => twiddle_h_rsc_0_6_i_db,
      adrb => twiddle_h_rsc_0_6_i_adrb,
      qa => twiddle_h_rsc_0_6_i_qa,
      wea => twiddle_h_rsc_0_6_wea,
      da => twiddle_h_rsc_0_6_i_da,
      adra => twiddle_h_rsc_0_6_i_adra,
      adra_d => twiddle_h_rsc_0_6_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => twiddle_h_rsc_0_6_i_da_d,
      qa_d => twiddle_h_rsc_0_6_i_qa_d_1,
      wea_d => twiddle_h_rsc_0_6_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => twiddle_h_rsc_0_6_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  twiddle_h_rsc_0_6_i_qb <= twiddle_h_rsc_0_6_qb;
  twiddle_h_rsc_0_6_db <= twiddle_h_rsc_0_6_i_db;
  twiddle_h_rsc_0_6_adrb <= twiddle_h_rsc_0_6_i_adrb;
  twiddle_h_rsc_0_6_i_qa <= twiddle_h_rsc_0_6_qa;
  twiddle_h_rsc_0_6_da <= twiddle_h_rsc_0_6_i_da;
  twiddle_h_rsc_0_6_adra <= twiddle_h_rsc_0_6_i_adra;
  twiddle_h_rsc_0_6_i_adra_d_1 <= STD_LOGIC_VECTOR'( "00000000") & twiddle_h_rsc_0_6_i_adra_d;
  twiddle_h_rsc_0_6_i_da_d <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
  twiddle_h_rsc_0_6_i_qa_d <= twiddle_h_rsc_0_6_i_qa_d_1;
  twiddle_h_rsc_0_6_i_wea_d <= STD_LOGIC_VECTOR'( "00");
  twiddle_h_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= twiddle_h_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_h_rsc_0_6_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( "00");

  twiddle_h_rsc_0_7_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_542_8_32_256_256_32_1_gen
    PORT MAP(
      qb => twiddle_h_rsc_0_7_i_qb,
      web => twiddle_h_rsc_0_7_web,
      db => twiddle_h_rsc_0_7_i_db,
      adrb => twiddle_h_rsc_0_7_i_adrb,
      qa => twiddle_h_rsc_0_7_i_qa,
      wea => twiddle_h_rsc_0_7_wea,
      da => twiddle_h_rsc_0_7_i_da,
      adra => twiddle_h_rsc_0_7_i_adra,
      adra_d => twiddle_h_rsc_0_7_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => twiddle_h_rsc_0_7_i_da_d,
      qa_d => twiddle_h_rsc_0_7_i_qa_d_1,
      wea_d => twiddle_h_rsc_0_7_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => twiddle_h_rsc_0_7_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  twiddle_h_rsc_0_7_i_qb <= twiddle_h_rsc_0_7_qb;
  twiddle_h_rsc_0_7_db <= twiddle_h_rsc_0_7_i_db;
  twiddle_h_rsc_0_7_adrb <= twiddle_h_rsc_0_7_i_adrb;
  twiddle_h_rsc_0_7_i_qa <= twiddle_h_rsc_0_7_qa;
  twiddle_h_rsc_0_7_da <= twiddle_h_rsc_0_7_i_da;
  twiddle_h_rsc_0_7_adra <= twiddle_h_rsc_0_7_i_adra;
  twiddle_h_rsc_0_7_i_adra_d_1 <= STD_LOGIC_VECTOR'( "00000000") & twiddle_h_rsc_0_7_i_adra_d;
  twiddle_h_rsc_0_7_i_da_d <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
  twiddle_h_rsc_0_7_i_qa_d <= twiddle_h_rsc_0_7_i_qa_d_1;
  twiddle_h_rsc_0_7_i_wea_d <= STD_LOGIC_VECTOR'( "00");
  twiddle_h_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= twiddle_h_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_h_rsc_0_7_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( "00");

  twiddle_h_rsc_0_8_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_543_8_32_256_256_32_1_gen
    PORT MAP(
      qb => twiddle_h_rsc_0_8_i_qb,
      web => twiddle_h_rsc_0_8_web,
      db => twiddle_h_rsc_0_8_i_db,
      adrb => twiddle_h_rsc_0_8_i_adrb,
      qa => twiddle_h_rsc_0_8_i_qa,
      wea => twiddle_h_rsc_0_8_wea,
      da => twiddle_h_rsc_0_8_i_da,
      adra => twiddle_h_rsc_0_8_i_adra,
      adra_d => twiddle_h_rsc_0_8_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => twiddle_h_rsc_0_8_i_da_d,
      qa_d => twiddle_h_rsc_0_8_i_qa_d_1,
      wea_d => twiddle_h_rsc_0_8_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => twiddle_h_rsc_0_8_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  twiddle_h_rsc_0_8_i_qb <= twiddle_h_rsc_0_8_qb;
  twiddle_h_rsc_0_8_db <= twiddle_h_rsc_0_8_i_db;
  twiddle_h_rsc_0_8_adrb <= twiddle_h_rsc_0_8_i_adrb;
  twiddle_h_rsc_0_8_i_qa <= twiddle_h_rsc_0_8_qa;
  twiddle_h_rsc_0_8_da <= twiddle_h_rsc_0_8_i_da;
  twiddle_h_rsc_0_8_adra <= twiddle_h_rsc_0_8_i_adra;
  twiddle_h_rsc_0_8_i_adra_d_1 <= STD_LOGIC_VECTOR'( "00000000") & twiddle_h_rsc_0_8_i_adra_d;
  twiddle_h_rsc_0_8_i_da_d <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
  twiddle_h_rsc_0_8_i_qa_d <= twiddle_h_rsc_0_8_i_qa_d_1;
  twiddle_h_rsc_0_8_i_wea_d <= STD_LOGIC_VECTOR'( "00");
  twiddle_h_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= twiddle_h_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_h_rsc_0_8_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( "00");

  twiddle_h_rsc_0_9_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_544_8_32_256_256_32_1_gen
    PORT MAP(
      qb => twiddle_h_rsc_0_9_i_qb,
      web => twiddle_h_rsc_0_9_web,
      db => twiddle_h_rsc_0_9_i_db,
      adrb => twiddle_h_rsc_0_9_i_adrb,
      qa => twiddle_h_rsc_0_9_i_qa,
      wea => twiddle_h_rsc_0_9_wea,
      da => twiddle_h_rsc_0_9_i_da,
      adra => twiddle_h_rsc_0_9_i_adra,
      adra_d => twiddle_h_rsc_0_9_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => twiddle_h_rsc_0_9_i_da_d,
      qa_d => twiddle_h_rsc_0_9_i_qa_d_1,
      wea_d => twiddle_h_rsc_0_9_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => twiddle_h_rsc_0_9_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  twiddle_h_rsc_0_9_i_qb <= twiddle_h_rsc_0_9_qb;
  twiddle_h_rsc_0_9_db <= twiddle_h_rsc_0_9_i_db;
  twiddle_h_rsc_0_9_adrb <= twiddle_h_rsc_0_9_i_adrb;
  twiddle_h_rsc_0_9_i_qa <= twiddle_h_rsc_0_9_qa;
  twiddle_h_rsc_0_9_da <= twiddle_h_rsc_0_9_i_da;
  twiddle_h_rsc_0_9_adra <= twiddle_h_rsc_0_9_i_adra;
  twiddle_h_rsc_0_9_i_adra_d_1 <= STD_LOGIC_VECTOR'( "00000000") & twiddle_h_rsc_0_9_i_adra_d;
  twiddle_h_rsc_0_9_i_da_d <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
  twiddle_h_rsc_0_9_i_qa_d <= twiddle_h_rsc_0_9_i_qa_d_1;
  twiddle_h_rsc_0_9_i_wea_d <= STD_LOGIC_VECTOR'( "00");
  twiddle_h_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= twiddle_h_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_h_rsc_0_9_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( "00");

  twiddle_h_rsc_0_10_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_545_8_32_256_256_32_1_gen
    PORT MAP(
      qb => twiddle_h_rsc_0_10_i_qb,
      web => twiddle_h_rsc_0_10_web,
      db => twiddle_h_rsc_0_10_i_db,
      adrb => twiddle_h_rsc_0_10_i_adrb,
      qa => twiddle_h_rsc_0_10_i_qa,
      wea => twiddle_h_rsc_0_10_wea,
      da => twiddle_h_rsc_0_10_i_da,
      adra => twiddle_h_rsc_0_10_i_adra,
      adra_d => twiddle_h_rsc_0_10_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => twiddle_h_rsc_0_10_i_da_d,
      qa_d => twiddle_h_rsc_0_10_i_qa_d_1,
      wea_d => twiddle_h_rsc_0_10_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => twiddle_h_rsc_0_10_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  twiddle_h_rsc_0_10_i_qb <= twiddle_h_rsc_0_10_qb;
  twiddle_h_rsc_0_10_db <= twiddle_h_rsc_0_10_i_db;
  twiddle_h_rsc_0_10_adrb <= twiddle_h_rsc_0_10_i_adrb;
  twiddle_h_rsc_0_10_i_qa <= twiddle_h_rsc_0_10_qa;
  twiddle_h_rsc_0_10_da <= twiddle_h_rsc_0_10_i_da;
  twiddle_h_rsc_0_10_adra <= twiddle_h_rsc_0_10_i_adra;
  twiddle_h_rsc_0_10_i_adra_d_1 <= STD_LOGIC_VECTOR'( "00000000") & twiddle_h_rsc_0_10_i_adra_d;
  twiddle_h_rsc_0_10_i_da_d <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
  twiddle_h_rsc_0_10_i_qa_d <= twiddle_h_rsc_0_10_i_qa_d_1;
  twiddle_h_rsc_0_10_i_wea_d <= STD_LOGIC_VECTOR'( "00");
  twiddle_h_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= twiddle_h_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_h_rsc_0_10_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( "00");

  twiddle_h_rsc_0_11_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_546_8_32_256_256_32_1_gen
    PORT MAP(
      qb => twiddle_h_rsc_0_11_i_qb,
      web => twiddle_h_rsc_0_11_web,
      db => twiddle_h_rsc_0_11_i_db,
      adrb => twiddle_h_rsc_0_11_i_adrb,
      qa => twiddle_h_rsc_0_11_i_qa,
      wea => twiddle_h_rsc_0_11_wea,
      da => twiddle_h_rsc_0_11_i_da,
      adra => twiddle_h_rsc_0_11_i_adra,
      adra_d => twiddle_h_rsc_0_11_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => twiddle_h_rsc_0_11_i_da_d,
      qa_d => twiddle_h_rsc_0_11_i_qa_d_1,
      wea_d => twiddle_h_rsc_0_11_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => twiddle_h_rsc_0_11_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  twiddle_h_rsc_0_11_i_qb <= twiddle_h_rsc_0_11_qb;
  twiddle_h_rsc_0_11_db <= twiddle_h_rsc_0_11_i_db;
  twiddle_h_rsc_0_11_adrb <= twiddle_h_rsc_0_11_i_adrb;
  twiddle_h_rsc_0_11_i_qa <= twiddle_h_rsc_0_11_qa;
  twiddle_h_rsc_0_11_da <= twiddle_h_rsc_0_11_i_da;
  twiddle_h_rsc_0_11_adra <= twiddle_h_rsc_0_11_i_adra;
  twiddle_h_rsc_0_11_i_adra_d_1 <= STD_LOGIC_VECTOR'( "00000000") & twiddle_h_rsc_0_11_i_adra_d;
  twiddle_h_rsc_0_11_i_da_d <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
  twiddle_h_rsc_0_11_i_qa_d <= twiddle_h_rsc_0_11_i_qa_d_1;
  twiddle_h_rsc_0_11_i_wea_d <= STD_LOGIC_VECTOR'( "00");
  twiddle_h_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= twiddle_h_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_h_rsc_0_11_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( "00");

  twiddle_h_rsc_0_12_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_547_8_32_256_256_32_1_gen
    PORT MAP(
      qb => twiddle_h_rsc_0_12_i_qb,
      web => twiddle_h_rsc_0_12_web,
      db => twiddle_h_rsc_0_12_i_db,
      adrb => twiddle_h_rsc_0_12_i_adrb,
      qa => twiddle_h_rsc_0_12_i_qa,
      wea => twiddle_h_rsc_0_12_wea,
      da => twiddle_h_rsc_0_12_i_da,
      adra => twiddle_h_rsc_0_12_i_adra,
      adra_d => twiddle_h_rsc_0_12_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => twiddle_h_rsc_0_12_i_da_d,
      qa_d => twiddle_h_rsc_0_12_i_qa_d_1,
      wea_d => twiddle_h_rsc_0_12_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => twiddle_h_rsc_0_12_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  twiddle_h_rsc_0_12_i_qb <= twiddle_h_rsc_0_12_qb;
  twiddle_h_rsc_0_12_db <= twiddle_h_rsc_0_12_i_db;
  twiddle_h_rsc_0_12_adrb <= twiddle_h_rsc_0_12_i_adrb;
  twiddle_h_rsc_0_12_i_qa <= twiddle_h_rsc_0_12_qa;
  twiddle_h_rsc_0_12_da <= twiddle_h_rsc_0_12_i_da;
  twiddle_h_rsc_0_12_adra <= twiddle_h_rsc_0_12_i_adra;
  twiddle_h_rsc_0_12_i_adra_d_1 <= STD_LOGIC_VECTOR'( "00000000") & twiddle_h_rsc_0_12_i_adra_d;
  twiddle_h_rsc_0_12_i_da_d <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
  twiddle_h_rsc_0_12_i_qa_d <= twiddle_h_rsc_0_12_i_qa_d_1;
  twiddle_h_rsc_0_12_i_wea_d <= STD_LOGIC_VECTOR'( "00");
  twiddle_h_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= twiddle_h_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_h_rsc_0_12_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( "00");

  twiddle_h_rsc_0_13_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_548_8_32_256_256_32_1_gen
    PORT MAP(
      qb => twiddle_h_rsc_0_13_i_qb,
      web => twiddle_h_rsc_0_13_web,
      db => twiddle_h_rsc_0_13_i_db,
      adrb => twiddle_h_rsc_0_13_i_adrb,
      qa => twiddle_h_rsc_0_13_i_qa,
      wea => twiddle_h_rsc_0_13_wea,
      da => twiddle_h_rsc_0_13_i_da,
      adra => twiddle_h_rsc_0_13_i_adra,
      adra_d => twiddle_h_rsc_0_13_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => twiddle_h_rsc_0_13_i_da_d,
      qa_d => twiddle_h_rsc_0_13_i_qa_d_1,
      wea_d => twiddle_h_rsc_0_13_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => twiddle_h_rsc_0_13_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  twiddle_h_rsc_0_13_i_qb <= twiddle_h_rsc_0_13_qb;
  twiddle_h_rsc_0_13_db <= twiddle_h_rsc_0_13_i_db;
  twiddle_h_rsc_0_13_adrb <= twiddle_h_rsc_0_13_i_adrb;
  twiddle_h_rsc_0_13_i_qa <= twiddle_h_rsc_0_13_qa;
  twiddle_h_rsc_0_13_da <= twiddle_h_rsc_0_13_i_da;
  twiddle_h_rsc_0_13_adra <= twiddle_h_rsc_0_13_i_adra;
  twiddle_h_rsc_0_13_i_adra_d_1 <= STD_LOGIC_VECTOR'( "00000000") & twiddle_h_rsc_0_13_i_adra_d;
  twiddle_h_rsc_0_13_i_da_d <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
  twiddle_h_rsc_0_13_i_qa_d <= twiddle_h_rsc_0_13_i_qa_d_1;
  twiddle_h_rsc_0_13_i_wea_d <= STD_LOGIC_VECTOR'( "00");
  twiddle_h_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= twiddle_h_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_h_rsc_0_13_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( "00");

  twiddle_h_rsc_0_14_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_549_8_32_256_256_32_1_gen
    PORT MAP(
      qb => twiddle_h_rsc_0_14_i_qb,
      web => twiddle_h_rsc_0_14_web,
      db => twiddle_h_rsc_0_14_i_db,
      adrb => twiddle_h_rsc_0_14_i_adrb,
      qa => twiddle_h_rsc_0_14_i_qa,
      wea => twiddle_h_rsc_0_14_wea,
      da => twiddle_h_rsc_0_14_i_da,
      adra => twiddle_h_rsc_0_14_i_adra,
      adra_d => twiddle_h_rsc_0_14_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => twiddle_h_rsc_0_14_i_da_d,
      qa_d => twiddle_h_rsc_0_14_i_qa_d_1,
      wea_d => twiddle_h_rsc_0_14_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => twiddle_h_rsc_0_14_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  twiddle_h_rsc_0_14_i_qb <= twiddle_h_rsc_0_14_qb;
  twiddle_h_rsc_0_14_db <= twiddle_h_rsc_0_14_i_db;
  twiddle_h_rsc_0_14_adrb <= twiddle_h_rsc_0_14_i_adrb;
  twiddle_h_rsc_0_14_i_qa <= twiddle_h_rsc_0_14_qa;
  twiddle_h_rsc_0_14_da <= twiddle_h_rsc_0_14_i_da;
  twiddle_h_rsc_0_14_adra <= twiddle_h_rsc_0_14_i_adra;
  twiddle_h_rsc_0_14_i_adra_d_1 <= STD_LOGIC_VECTOR'( "00000000") & twiddle_h_rsc_0_14_i_adra_d;
  twiddle_h_rsc_0_14_i_da_d <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
  twiddle_h_rsc_0_14_i_qa_d <= twiddle_h_rsc_0_14_i_qa_d_1;
  twiddle_h_rsc_0_14_i_wea_d <= STD_LOGIC_VECTOR'( "00");
  twiddle_h_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= twiddle_h_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_h_rsc_0_14_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( "00");

  twiddle_h_rsc_0_15_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_550_8_32_256_256_32_1_gen
    PORT MAP(
      qb => twiddle_h_rsc_0_15_i_qb,
      web => twiddle_h_rsc_0_15_web,
      db => twiddle_h_rsc_0_15_i_db,
      adrb => twiddle_h_rsc_0_15_i_adrb,
      qa => twiddle_h_rsc_0_15_i_qa,
      wea => twiddle_h_rsc_0_15_wea,
      da => twiddle_h_rsc_0_15_i_da,
      adra => twiddle_h_rsc_0_15_i_adra,
      adra_d => twiddle_h_rsc_0_15_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => twiddle_h_rsc_0_15_i_da_d,
      qa_d => twiddle_h_rsc_0_15_i_qa_d_1,
      wea_d => twiddle_h_rsc_0_15_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => twiddle_h_rsc_0_15_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  twiddle_h_rsc_0_15_i_qb <= twiddle_h_rsc_0_15_qb;
  twiddle_h_rsc_0_15_db <= twiddle_h_rsc_0_15_i_db;
  twiddle_h_rsc_0_15_adrb <= twiddle_h_rsc_0_15_i_adrb;
  twiddle_h_rsc_0_15_i_qa <= twiddle_h_rsc_0_15_qa;
  twiddle_h_rsc_0_15_da <= twiddle_h_rsc_0_15_i_da;
  twiddle_h_rsc_0_15_adra <= twiddle_h_rsc_0_15_i_adra;
  twiddle_h_rsc_0_15_i_adra_d_1 <= STD_LOGIC_VECTOR'( "00000000") & twiddle_h_rsc_0_15_i_adra_d;
  twiddle_h_rsc_0_15_i_da_d <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
  twiddle_h_rsc_0_15_i_qa_d <= twiddle_h_rsc_0_15_i_qa_d_1;
  twiddle_h_rsc_0_15_i_wea_d <= STD_LOGIC_VECTOR'( "00");
  twiddle_h_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= twiddle_h_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_h_rsc_0_15_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( "00");

  peaseNTT_core_inst : peaseNTT_core
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_triosy_0_0_lz => xt_rsc_triosy_0_0_lz,
      xt_rsc_triosy_0_1_lz => xt_rsc_triosy_0_1_lz,
      xt_rsc_triosy_0_2_lz => xt_rsc_triosy_0_2_lz,
      xt_rsc_triosy_0_3_lz => xt_rsc_triosy_0_3_lz,
      xt_rsc_triosy_0_4_lz => xt_rsc_triosy_0_4_lz,
      xt_rsc_triosy_0_5_lz => xt_rsc_triosy_0_5_lz,
      xt_rsc_triosy_0_6_lz => xt_rsc_triosy_0_6_lz,
      xt_rsc_triosy_0_7_lz => xt_rsc_triosy_0_7_lz,
      xt_rsc_triosy_0_8_lz => xt_rsc_triosy_0_8_lz,
      xt_rsc_triosy_0_9_lz => xt_rsc_triosy_0_9_lz,
      xt_rsc_triosy_0_10_lz => xt_rsc_triosy_0_10_lz,
      xt_rsc_triosy_0_11_lz => xt_rsc_triosy_0_11_lz,
      xt_rsc_triosy_0_12_lz => xt_rsc_triosy_0_12_lz,
      xt_rsc_triosy_0_13_lz => xt_rsc_triosy_0_13_lz,
      xt_rsc_triosy_0_14_lz => xt_rsc_triosy_0_14_lz,
      xt_rsc_triosy_0_15_lz => xt_rsc_triosy_0_15_lz,
      xt_rsc_triosy_0_16_lz => xt_rsc_triosy_0_16_lz,
      xt_rsc_triosy_0_17_lz => xt_rsc_triosy_0_17_lz,
      xt_rsc_triosy_0_18_lz => xt_rsc_triosy_0_18_lz,
      xt_rsc_triosy_0_19_lz => xt_rsc_triosy_0_19_lz,
      xt_rsc_triosy_0_20_lz => xt_rsc_triosy_0_20_lz,
      xt_rsc_triosy_0_21_lz => xt_rsc_triosy_0_21_lz,
      xt_rsc_triosy_0_22_lz => xt_rsc_triosy_0_22_lz,
      xt_rsc_triosy_0_23_lz => xt_rsc_triosy_0_23_lz,
      xt_rsc_triosy_0_24_lz => xt_rsc_triosy_0_24_lz,
      xt_rsc_triosy_0_25_lz => xt_rsc_triosy_0_25_lz,
      xt_rsc_triosy_0_26_lz => xt_rsc_triosy_0_26_lz,
      xt_rsc_triosy_0_27_lz => xt_rsc_triosy_0_27_lz,
      xt_rsc_triosy_0_28_lz => xt_rsc_triosy_0_28_lz,
      xt_rsc_triosy_0_29_lz => xt_rsc_triosy_0_29_lz,
      xt_rsc_triosy_0_30_lz => xt_rsc_triosy_0_30_lz,
      xt_rsc_triosy_0_31_lz => xt_rsc_triosy_0_31_lz,
      xt_rsc_triosy_1_0_lz => xt_rsc_triosy_1_0_lz,
      xt_rsc_triosy_1_1_lz => xt_rsc_triosy_1_1_lz,
      xt_rsc_triosy_1_2_lz => xt_rsc_triosy_1_2_lz,
      xt_rsc_triosy_1_3_lz => xt_rsc_triosy_1_3_lz,
      xt_rsc_triosy_1_4_lz => xt_rsc_triosy_1_4_lz,
      xt_rsc_triosy_1_5_lz => xt_rsc_triosy_1_5_lz,
      xt_rsc_triosy_1_6_lz => xt_rsc_triosy_1_6_lz,
      xt_rsc_triosy_1_7_lz => xt_rsc_triosy_1_7_lz,
      xt_rsc_triosy_1_8_lz => xt_rsc_triosy_1_8_lz,
      xt_rsc_triosy_1_9_lz => xt_rsc_triosy_1_9_lz,
      xt_rsc_triosy_1_10_lz => xt_rsc_triosy_1_10_lz,
      xt_rsc_triosy_1_11_lz => xt_rsc_triosy_1_11_lz,
      xt_rsc_triosy_1_12_lz => xt_rsc_triosy_1_12_lz,
      xt_rsc_triosy_1_13_lz => xt_rsc_triosy_1_13_lz,
      xt_rsc_triosy_1_14_lz => xt_rsc_triosy_1_14_lz,
      xt_rsc_triosy_1_15_lz => xt_rsc_triosy_1_15_lz,
      xt_rsc_triosy_1_16_lz => xt_rsc_triosy_1_16_lz,
      xt_rsc_triosy_1_17_lz => xt_rsc_triosy_1_17_lz,
      xt_rsc_triosy_1_18_lz => xt_rsc_triosy_1_18_lz,
      xt_rsc_triosy_1_19_lz => xt_rsc_triosy_1_19_lz,
      xt_rsc_triosy_1_20_lz => xt_rsc_triosy_1_20_lz,
      xt_rsc_triosy_1_21_lz => xt_rsc_triosy_1_21_lz,
      xt_rsc_triosy_1_22_lz => xt_rsc_triosy_1_22_lz,
      xt_rsc_triosy_1_23_lz => xt_rsc_triosy_1_23_lz,
      xt_rsc_triosy_1_24_lz => xt_rsc_triosy_1_24_lz,
      xt_rsc_triosy_1_25_lz => xt_rsc_triosy_1_25_lz,
      xt_rsc_triosy_1_26_lz => xt_rsc_triosy_1_26_lz,
      xt_rsc_triosy_1_27_lz => xt_rsc_triosy_1_27_lz,
      xt_rsc_triosy_1_28_lz => xt_rsc_triosy_1_28_lz,
      xt_rsc_triosy_1_29_lz => xt_rsc_triosy_1_29_lz,
      xt_rsc_triosy_1_30_lz => xt_rsc_triosy_1_30_lz,
      xt_rsc_triosy_1_31_lz => xt_rsc_triosy_1_31_lz,
      xt_rsc_triosy_2_0_lz => xt_rsc_triosy_2_0_lz,
      xt_rsc_triosy_2_1_lz => xt_rsc_triosy_2_1_lz,
      xt_rsc_triosy_2_2_lz => xt_rsc_triosy_2_2_lz,
      xt_rsc_triosy_2_3_lz => xt_rsc_triosy_2_3_lz,
      xt_rsc_triosy_2_4_lz => xt_rsc_triosy_2_4_lz,
      xt_rsc_triosy_2_5_lz => xt_rsc_triosy_2_5_lz,
      xt_rsc_triosy_2_6_lz => xt_rsc_triosy_2_6_lz,
      xt_rsc_triosy_2_7_lz => xt_rsc_triosy_2_7_lz,
      xt_rsc_triosy_2_8_lz => xt_rsc_triosy_2_8_lz,
      xt_rsc_triosy_2_9_lz => xt_rsc_triosy_2_9_lz,
      xt_rsc_triosy_2_10_lz => xt_rsc_triosy_2_10_lz,
      xt_rsc_triosy_2_11_lz => xt_rsc_triosy_2_11_lz,
      xt_rsc_triosy_2_12_lz => xt_rsc_triosy_2_12_lz,
      xt_rsc_triosy_2_13_lz => xt_rsc_triosy_2_13_lz,
      xt_rsc_triosy_2_14_lz => xt_rsc_triosy_2_14_lz,
      xt_rsc_triosy_2_15_lz => xt_rsc_triosy_2_15_lz,
      xt_rsc_triosy_2_16_lz => xt_rsc_triosy_2_16_lz,
      xt_rsc_triosy_2_17_lz => xt_rsc_triosy_2_17_lz,
      xt_rsc_triosy_2_18_lz => xt_rsc_triosy_2_18_lz,
      xt_rsc_triosy_2_19_lz => xt_rsc_triosy_2_19_lz,
      xt_rsc_triosy_2_20_lz => xt_rsc_triosy_2_20_lz,
      xt_rsc_triosy_2_21_lz => xt_rsc_triosy_2_21_lz,
      xt_rsc_triosy_2_22_lz => xt_rsc_triosy_2_22_lz,
      xt_rsc_triosy_2_23_lz => xt_rsc_triosy_2_23_lz,
      xt_rsc_triosy_2_24_lz => xt_rsc_triosy_2_24_lz,
      xt_rsc_triosy_2_25_lz => xt_rsc_triosy_2_25_lz,
      xt_rsc_triosy_2_26_lz => xt_rsc_triosy_2_26_lz,
      xt_rsc_triosy_2_27_lz => xt_rsc_triosy_2_27_lz,
      xt_rsc_triosy_2_28_lz => xt_rsc_triosy_2_28_lz,
      xt_rsc_triosy_2_29_lz => xt_rsc_triosy_2_29_lz,
      xt_rsc_triosy_2_30_lz => xt_rsc_triosy_2_30_lz,
      xt_rsc_triosy_2_31_lz => xt_rsc_triosy_2_31_lz,
      xt_rsc_triosy_3_0_lz => xt_rsc_triosy_3_0_lz,
      xt_rsc_triosy_3_1_lz => xt_rsc_triosy_3_1_lz,
      xt_rsc_triosy_3_2_lz => xt_rsc_triosy_3_2_lz,
      xt_rsc_triosy_3_3_lz => xt_rsc_triosy_3_3_lz,
      xt_rsc_triosy_3_4_lz => xt_rsc_triosy_3_4_lz,
      xt_rsc_triosy_3_5_lz => xt_rsc_triosy_3_5_lz,
      xt_rsc_triosy_3_6_lz => xt_rsc_triosy_3_6_lz,
      xt_rsc_triosy_3_7_lz => xt_rsc_triosy_3_7_lz,
      xt_rsc_triosy_3_8_lz => xt_rsc_triosy_3_8_lz,
      xt_rsc_triosy_3_9_lz => xt_rsc_triosy_3_9_lz,
      xt_rsc_triosy_3_10_lz => xt_rsc_triosy_3_10_lz,
      xt_rsc_triosy_3_11_lz => xt_rsc_triosy_3_11_lz,
      xt_rsc_triosy_3_12_lz => xt_rsc_triosy_3_12_lz,
      xt_rsc_triosy_3_13_lz => xt_rsc_triosy_3_13_lz,
      xt_rsc_triosy_3_14_lz => xt_rsc_triosy_3_14_lz,
      xt_rsc_triosy_3_15_lz => xt_rsc_triosy_3_15_lz,
      xt_rsc_triosy_3_16_lz => xt_rsc_triosy_3_16_lz,
      xt_rsc_triosy_3_17_lz => xt_rsc_triosy_3_17_lz,
      xt_rsc_triosy_3_18_lz => xt_rsc_triosy_3_18_lz,
      xt_rsc_triosy_3_19_lz => xt_rsc_triosy_3_19_lz,
      xt_rsc_triosy_3_20_lz => xt_rsc_triosy_3_20_lz,
      xt_rsc_triosy_3_21_lz => xt_rsc_triosy_3_21_lz,
      xt_rsc_triosy_3_22_lz => xt_rsc_triosy_3_22_lz,
      xt_rsc_triosy_3_23_lz => xt_rsc_triosy_3_23_lz,
      xt_rsc_triosy_3_24_lz => xt_rsc_triosy_3_24_lz,
      xt_rsc_triosy_3_25_lz => xt_rsc_triosy_3_25_lz,
      xt_rsc_triosy_3_26_lz => xt_rsc_triosy_3_26_lz,
      xt_rsc_triosy_3_27_lz => xt_rsc_triosy_3_27_lz,
      xt_rsc_triosy_3_28_lz => xt_rsc_triosy_3_28_lz,
      xt_rsc_triosy_3_29_lz => xt_rsc_triosy_3_29_lz,
      xt_rsc_triosy_3_30_lz => xt_rsc_triosy_3_30_lz,
      xt_rsc_triosy_3_31_lz => xt_rsc_triosy_3_31_lz,
      xt_rsc_triosy_4_0_lz => xt_rsc_triosy_4_0_lz,
      xt_rsc_triosy_4_1_lz => xt_rsc_triosy_4_1_lz,
      xt_rsc_triosy_4_2_lz => xt_rsc_triosy_4_2_lz,
      xt_rsc_triosy_4_3_lz => xt_rsc_triosy_4_3_lz,
      xt_rsc_triosy_4_4_lz => xt_rsc_triosy_4_4_lz,
      xt_rsc_triosy_4_5_lz => xt_rsc_triosy_4_5_lz,
      xt_rsc_triosy_4_6_lz => xt_rsc_triosy_4_6_lz,
      xt_rsc_triosy_4_7_lz => xt_rsc_triosy_4_7_lz,
      xt_rsc_triosy_4_8_lz => xt_rsc_triosy_4_8_lz,
      xt_rsc_triosy_4_9_lz => xt_rsc_triosy_4_9_lz,
      xt_rsc_triosy_4_10_lz => xt_rsc_triosy_4_10_lz,
      xt_rsc_triosy_4_11_lz => xt_rsc_triosy_4_11_lz,
      xt_rsc_triosy_4_12_lz => xt_rsc_triosy_4_12_lz,
      xt_rsc_triosy_4_13_lz => xt_rsc_triosy_4_13_lz,
      xt_rsc_triosy_4_14_lz => xt_rsc_triosy_4_14_lz,
      xt_rsc_triosy_4_15_lz => xt_rsc_triosy_4_15_lz,
      xt_rsc_triosy_4_16_lz => xt_rsc_triosy_4_16_lz,
      xt_rsc_triosy_4_17_lz => xt_rsc_triosy_4_17_lz,
      xt_rsc_triosy_4_18_lz => xt_rsc_triosy_4_18_lz,
      xt_rsc_triosy_4_19_lz => xt_rsc_triosy_4_19_lz,
      xt_rsc_triosy_4_20_lz => xt_rsc_triosy_4_20_lz,
      xt_rsc_triosy_4_21_lz => xt_rsc_triosy_4_21_lz,
      xt_rsc_triosy_4_22_lz => xt_rsc_triosy_4_22_lz,
      xt_rsc_triosy_4_23_lz => xt_rsc_triosy_4_23_lz,
      xt_rsc_triosy_4_24_lz => xt_rsc_triosy_4_24_lz,
      xt_rsc_triosy_4_25_lz => xt_rsc_triosy_4_25_lz,
      xt_rsc_triosy_4_26_lz => xt_rsc_triosy_4_26_lz,
      xt_rsc_triosy_4_27_lz => xt_rsc_triosy_4_27_lz,
      xt_rsc_triosy_4_28_lz => xt_rsc_triosy_4_28_lz,
      xt_rsc_triosy_4_29_lz => xt_rsc_triosy_4_29_lz,
      xt_rsc_triosy_4_30_lz => xt_rsc_triosy_4_30_lz,
      xt_rsc_triosy_4_31_lz => xt_rsc_triosy_4_31_lz,
      xt_rsc_triosy_5_0_lz => xt_rsc_triosy_5_0_lz,
      xt_rsc_triosy_5_1_lz => xt_rsc_triosy_5_1_lz,
      xt_rsc_triosy_5_2_lz => xt_rsc_triosy_5_2_lz,
      xt_rsc_triosy_5_3_lz => xt_rsc_triosy_5_3_lz,
      xt_rsc_triosy_5_4_lz => xt_rsc_triosy_5_4_lz,
      xt_rsc_triosy_5_5_lz => xt_rsc_triosy_5_5_lz,
      xt_rsc_triosy_5_6_lz => xt_rsc_triosy_5_6_lz,
      xt_rsc_triosy_5_7_lz => xt_rsc_triosy_5_7_lz,
      xt_rsc_triosy_5_8_lz => xt_rsc_triosy_5_8_lz,
      xt_rsc_triosy_5_9_lz => xt_rsc_triosy_5_9_lz,
      xt_rsc_triosy_5_10_lz => xt_rsc_triosy_5_10_lz,
      xt_rsc_triosy_5_11_lz => xt_rsc_triosy_5_11_lz,
      xt_rsc_triosy_5_12_lz => xt_rsc_triosy_5_12_lz,
      xt_rsc_triosy_5_13_lz => xt_rsc_triosy_5_13_lz,
      xt_rsc_triosy_5_14_lz => xt_rsc_triosy_5_14_lz,
      xt_rsc_triosy_5_15_lz => xt_rsc_triosy_5_15_lz,
      xt_rsc_triosy_5_16_lz => xt_rsc_triosy_5_16_lz,
      xt_rsc_triosy_5_17_lz => xt_rsc_triosy_5_17_lz,
      xt_rsc_triosy_5_18_lz => xt_rsc_triosy_5_18_lz,
      xt_rsc_triosy_5_19_lz => xt_rsc_triosy_5_19_lz,
      xt_rsc_triosy_5_20_lz => xt_rsc_triosy_5_20_lz,
      xt_rsc_triosy_5_21_lz => xt_rsc_triosy_5_21_lz,
      xt_rsc_triosy_5_22_lz => xt_rsc_triosy_5_22_lz,
      xt_rsc_triosy_5_23_lz => xt_rsc_triosy_5_23_lz,
      xt_rsc_triosy_5_24_lz => xt_rsc_triosy_5_24_lz,
      xt_rsc_triosy_5_25_lz => xt_rsc_triosy_5_25_lz,
      xt_rsc_triosy_5_26_lz => xt_rsc_triosy_5_26_lz,
      xt_rsc_triosy_5_27_lz => xt_rsc_triosy_5_27_lz,
      xt_rsc_triosy_5_28_lz => xt_rsc_triosy_5_28_lz,
      xt_rsc_triosy_5_29_lz => xt_rsc_triosy_5_29_lz,
      xt_rsc_triosy_5_30_lz => xt_rsc_triosy_5_30_lz,
      xt_rsc_triosy_5_31_lz => xt_rsc_triosy_5_31_lz,
      xt_rsc_triosy_6_0_lz => xt_rsc_triosy_6_0_lz,
      xt_rsc_triosy_6_1_lz => xt_rsc_triosy_6_1_lz,
      xt_rsc_triosy_6_2_lz => xt_rsc_triosy_6_2_lz,
      xt_rsc_triosy_6_3_lz => xt_rsc_triosy_6_3_lz,
      xt_rsc_triosy_6_4_lz => xt_rsc_triosy_6_4_lz,
      xt_rsc_triosy_6_5_lz => xt_rsc_triosy_6_5_lz,
      xt_rsc_triosy_6_6_lz => xt_rsc_triosy_6_6_lz,
      xt_rsc_triosy_6_7_lz => xt_rsc_triosy_6_7_lz,
      xt_rsc_triosy_6_8_lz => xt_rsc_triosy_6_8_lz,
      xt_rsc_triosy_6_9_lz => xt_rsc_triosy_6_9_lz,
      xt_rsc_triosy_6_10_lz => xt_rsc_triosy_6_10_lz,
      xt_rsc_triosy_6_11_lz => xt_rsc_triosy_6_11_lz,
      xt_rsc_triosy_6_12_lz => xt_rsc_triosy_6_12_lz,
      xt_rsc_triosy_6_13_lz => xt_rsc_triosy_6_13_lz,
      xt_rsc_triosy_6_14_lz => xt_rsc_triosy_6_14_lz,
      xt_rsc_triosy_6_15_lz => xt_rsc_triosy_6_15_lz,
      xt_rsc_triosy_6_16_lz => xt_rsc_triosy_6_16_lz,
      xt_rsc_triosy_6_17_lz => xt_rsc_triosy_6_17_lz,
      xt_rsc_triosy_6_18_lz => xt_rsc_triosy_6_18_lz,
      xt_rsc_triosy_6_19_lz => xt_rsc_triosy_6_19_lz,
      xt_rsc_triosy_6_20_lz => xt_rsc_triosy_6_20_lz,
      xt_rsc_triosy_6_21_lz => xt_rsc_triosy_6_21_lz,
      xt_rsc_triosy_6_22_lz => xt_rsc_triosy_6_22_lz,
      xt_rsc_triosy_6_23_lz => xt_rsc_triosy_6_23_lz,
      xt_rsc_triosy_6_24_lz => xt_rsc_triosy_6_24_lz,
      xt_rsc_triosy_6_25_lz => xt_rsc_triosy_6_25_lz,
      xt_rsc_triosy_6_26_lz => xt_rsc_triosy_6_26_lz,
      xt_rsc_triosy_6_27_lz => xt_rsc_triosy_6_27_lz,
      xt_rsc_triosy_6_28_lz => xt_rsc_triosy_6_28_lz,
      xt_rsc_triosy_6_29_lz => xt_rsc_triosy_6_29_lz,
      xt_rsc_triosy_6_30_lz => xt_rsc_triosy_6_30_lz,
      xt_rsc_triosy_6_31_lz => xt_rsc_triosy_6_31_lz,
      xt_rsc_triosy_7_0_lz => xt_rsc_triosy_7_0_lz,
      xt_rsc_triosy_7_1_lz => xt_rsc_triosy_7_1_lz,
      xt_rsc_triosy_7_2_lz => xt_rsc_triosy_7_2_lz,
      xt_rsc_triosy_7_3_lz => xt_rsc_triosy_7_3_lz,
      xt_rsc_triosy_7_4_lz => xt_rsc_triosy_7_4_lz,
      xt_rsc_triosy_7_5_lz => xt_rsc_triosy_7_5_lz,
      xt_rsc_triosy_7_6_lz => xt_rsc_triosy_7_6_lz,
      xt_rsc_triosy_7_7_lz => xt_rsc_triosy_7_7_lz,
      xt_rsc_triosy_7_8_lz => xt_rsc_triosy_7_8_lz,
      xt_rsc_triosy_7_9_lz => xt_rsc_triosy_7_9_lz,
      xt_rsc_triosy_7_10_lz => xt_rsc_triosy_7_10_lz,
      xt_rsc_triosy_7_11_lz => xt_rsc_triosy_7_11_lz,
      xt_rsc_triosy_7_12_lz => xt_rsc_triosy_7_12_lz,
      xt_rsc_triosy_7_13_lz => xt_rsc_triosy_7_13_lz,
      xt_rsc_triosy_7_14_lz => xt_rsc_triosy_7_14_lz,
      xt_rsc_triosy_7_15_lz => xt_rsc_triosy_7_15_lz,
      xt_rsc_triosy_7_16_lz => xt_rsc_triosy_7_16_lz,
      xt_rsc_triosy_7_17_lz => xt_rsc_triosy_7_17_lz,
      xt_rsc_triosy_7_18_lz => xt_rsc_triosy_7_18_lz,
      xt_rsc_triosy_7_19_lz => xt_rsc_triosy_7_19_lz,
      xt_rsc_triosy_7_20_lz => xt_rsc_triosy_7_20_lz,
      xt_rsc_triosy_7_21_lz => xt_rsc_triosy_7_21_lz,
      xt_rsc_triosy_7_22_lz => xt_rsc_triosy_7_22_lz,
      xt_rsc_triosy_7_23_lz => xt_rsc_triosy_7_23_lz,
      xt_rsc_triosy_7_24_lz => xt_rsc_triosy_7_24_lz,
      xt_rsc_triosy_7_25_lz => xt_rsc_triosy_7_25_lz,
      xt_rsc_triosy_7_26_lz => xt_rsc_triosy_7_26_lz,
      xt_rsc_triosy_7_27_lz => xt_rsc_triosy_7_27_lz,
      xt_rsc_triosy_7_28_lz => xt_rsc_triosy_7_28_lz,
      xt_rsc_triosy_7_29_lz => xt_rsc_triosy_7_29_lz,
      xt_rsc_triosy_7_30_lz => xt_rsc_triosy_7_30_lz,
      xt_rsc_triosy_7_31_lz => xt_rsc_triosy_7_31_lz,
      p_rsc_dat => peaseNTT_core_inst_p_rsc_dat,
      p_rsc_triosy_lz => p_rsc_triosy_lz,
      r_rsc_triosy_lz => r_rsc_triosy_lz,
      twiddle_rsc_triosy_0_0_lz => twiddle_rsc_triosy_0_0_lz,
      twiddle_rsc_triosy_0_1_lz => twiddle_rsc_triosy_0_1_lz,
      twiddle_rsc_triosy_0_2_lz => twiddle_rsc_triosy_0_2_lz,
      twiddle_rsc_triosy_0_3_lz => twiddle_rsc_triosy_0_3_lz,
      twiddle_rsc_triosy_0_4_lz => twiddle_rsc_triosy_0_4_lz,
      twiddle_rsc_triosy_0_5_lz => twiddle_rsc_triosy_0_5_lz,
      twiddle_rsc_triosy_0_6_lz => twiddle_rsc_triosy_0_6_lz,
      twiddle_rsc_triosy_0_7_lz => twiddle_rsc_triosy_0_7_lz,
      twiddle_rsc_triosy_0_8_lz => twiddle_rsc_triosy_0_8_lz,
      twiddle_rsc_triosy_0_9_lz => twiddle_rsc_triosy_0_9_lz,
      twiddle_rsc_triosy_0_10_lz => twiddle_rsc_triosy_0_10_lz,
      twiddle_rsc_triosy_0_11_lz => twiddle_rsc_triosy_0_11_lz,
      twiddle_rsc_triosy_0_12_lz => twiddle_rsc_triosy_0_12_lz,
      twiddle_rsc_triosy_0_13_lz => twiddle_rsc_triosy_0_13_lz,
      twiddle_rsc_triosy_0_14_lz => twiddle_rsc_triosy_0_14_lz,
      twiddle_rsc_triosy_0_15_lz => twiddle_rsc_triosy_0_15_lz,
      twiddle_h_rsc_triosy_0_0_lz => twiddle_h_rsc_triosy_0_0_lz,
      twiddle_h_rsc_triosy_0_1_lz => twiddle_h_rsc_triosy_0_1_lz,
      twiddle_h_rsc_triosy_0_2_lz => twiddle_h_rsc_triosy_0_2_lz,
      twiddle_h_rsc_triosy_0_3_lz => twiddle_h_rsc_triosy_0_3_lz,
      twiddle_h_rsc_triosy_0_4_lz => twiddle_h_rsc_triosy_0_4_lz,
      twiddle_h_rsc_triosy_0_5_lz => twiddle_h_rsc_triosy_0_5_lz,
      twiddle_h_rsc_triosy_0_6_lz => twiddle_h_rsc_triosy_0_6_lz,
      twiddle_h_rsc_triosy_0_7_lz => twiddle_h_rsc_triosy_0_7_lz,
      twiddle_h_rsc_triosy_0_8_lz => twiddle_h_rsc_triosy_0_8_lz,
      twiddle_h_rsc_triosy_0_9_lz => twiddle_h_rsc_triosy_0_9_lz,
      twiddle_h_rsc_triosy_0_10_lz => twiddle_h_rsc_triosy_0_10_lz,
      twiddle_h_rsc_triosy_0_11_lz => twiddle_h_rsc_triosy_0_11_lz,
      twiddle_h_rsc_triosy_0_12_lz => twiddle_h_rsc_triosy_0_12_lz,
      twiddle_h_rsc_triosy_0_13_lz => twiddle_h_rsc_triosy_0_13_lz,
      twiddle_h_rsc_triosy_0_14_lz => twiddle_h_rsc_triosy_0_14_lz,
      twiddle_h_rsc_triosy_0_15_lz => twiddle_h_rsc_triosy_0_15_lz,
      yt_rsc_0_0_i_clkr_en_d => yt_rsc_0_0_i_clkr_en_d,
      yt_rsc_0_0_i_q_d => peaseNTT_core_inst_yt_rsc_0_0_i_q_d,
      yt_rsc_0_1_i_q_d => peaseNTT_core_inst_yt_rsc_0_1_i_q_d,
      yt_rsc_0_2_i_q_d => peaseNTT_core_inst_yt_rsc_0_2_i_q_d,
      yt_rsc_0_3_i_q_d => peaseNTT_core_inst_yt_rsc_0_3_i_q_d,
      yt_rsc_0_4_i_q_d => peaseNTT_core_inst_yt_rsc_0_4_i_q_d,
      yt_rsc_0_5_i_q_d => peaseNTT_core_inst_yt_rsc_0_5_i_q_d,
      yt_rsc_0_6_i_q_d => peaseNTT_core_inst_yt_rsc_0_6_i_q_d,
      yt_rsc_0_7_i_q_d => peaseNTT_core_inst_yt_rsc_0_7_i_q_d,
      yt_rsc_0_8_i_q_d => peaseNTT_core_inst_yt_rsc_0_8_i_q_d,
      yt_rsc_0_9_i_q_d => peaseNTT_core_inst_yt_rsc_0_9_i_q_d,
      yt_rsc_0_10_i_q_d => peaseNTT_core_inst_yt_rsc_0_10_i_q_d,
      yt_rsc_0_11_i_q_d => peaseNTT_core_inst_yt_rsc_0_11_i_q_d,
      yt_rsc_0_12_i_q_d => peaseNTT_core_inst_yt_rsc_0_12_i_q_d,
      yt_rsc_0_13_i_q_d => peaseNTT_core_inst_yt_rsc_0_13_i_q_d,
      yt_rsc_0_14_i_q_d => peaseNTT_core_inst_yt_rsc_0_14_i_q_d,
      yt_rsc_0_15_i_q_d => peaseNTT_core_inst_yt_rsc_0_15_i_q_d,
      yt_rsc_0_16_i_clkr_en_d => yt_rsc_0_16_i_clkr_en_d,
      yt_rsc_0_16_i_q_d => peaseNTT_core_inst_yt_rsc_0_16_i_q_d,
      yt_rsc_0_17_i_q_d => peaseNTT_core_inst_yt_rsc_0_17_i_q_d,
      yt_rsc_0_18_i_q_d => peaseNTT_core_inst_yt_rsc_0_18_i_q_d,
      yt_rsc_0_19_i_q_d => peaseNTT_core_inst_yt_rsc_0_19_i_q_d,
      yt_rsc_0_20_i_q_d => peaseNTT_core_inst_yt_rsc_0_20_i_q_d,
      yt_rsc_0_21_i_q_d => peaseNTT_core_inst_yt_rsc_0_21_i_q_d,
      yt_rsc_0_22_i_q_d => peaseNTT_core_inst_yt_rsc_0_22_i_q_d,
      yt_rsc_0_23_i_q_d => peaseNTT_core_inst_yt_rsc_0_23_i_q_d,
      yt_rsc_0_24_i_q_d => peaseNTT_core_inst_yt_rsc_0_24_i_q_d,
      yt_rsc_0_25_i_q_d => peaseNTT_core_inst_yt_rsc_0_25_i_q_d,
      yt_rsc_0_26_i_q_d => peaseNTT_core_inst_yt_rsc_0_26_i_q_d,
      yt_rsc_0_27_i_q_d => peaseNTT_core_inst_yt_rsc_0_27_i_q_d,
      yt_rsc_0_28_i_q_d => peaseNTT_core_inst_yt_rsc_0_28_i_q_d,
      yt_rsc_0_29_i_q_d => peaseNTT_core_inst_yt_rsc_0_29_i_q_d,
      yt_rsc_0_30_i_q_d => peaseNTT_core_inst_yt_rsc_0_30_i_q_d,
      yt_rsc_0_31_i_q_d => peaseNTT_core_inst_yt_rsc_0_31_i_q_d,
      yt_rsc_1_0_i_clkr_en_d => yt_rsc_1_0_i_clkr_en_d,
      yt_rsc_1_0_i_q_d => peaseNTT_core_inst_yt_rsc_1_0_i_q_d,
      yt_rsc_1_1_i_q_d => peaseNTT_core_inst_yt_rsc_1_1_i_q_d,
      yt_rsc_1_2_i_q_d => peaseNTT_core_inst_yt_rsc_1_2_i_q_d,
      yt_rsc_1_3_i_q_d => peaseNTT_core_inst_yt_rsc_1_3_i_q_d,
      yt_rsc_1_4_i_q_d => peaseNTT_core_inst_yt_rsc_1_4_i_q_d,
      yt_rsc_1_5_i_q_d => peaseNTT_core_inst_yt_rsc_1_5_i_q_d,
      yt_rsc_1_6_i_q_d => peaseNTT_core_inst_yt_rsc_1_6_i_q_d,
      yt_rsc_1_7_i_q_d => peaseNTT_core_inst_yt_rsc_1_7_i_q_d,
      yt_rsc_1_8_i_q_d => peaseNTT_core_inst_yt_rsc_1_8_i_q_d,
      yt_rsc_1_9_i_q_d => peaseNTT_core_inst_yt_rsc_1_9_i_q_d,
      yt_rsc_1_10_i_q_d => peaseNTT_core_inst_yt_rsc_1_10_i_q_d,
      yt_rsc_1_11_i_q_d => peaseNTT_core_inst_yt_rsc_1_11_i_q_d,
      yt_rsc_1_12_i_q_d => peaseNTT_core_inst_yt_rsc_1_12_i_q_d,
      yt_rsc_1_13_i_q_d => peaseNTT_core_inst_yt_rsc_1_13_i_q_d,
      yt_rsc_1_14_i_q_d => peaseNTT_core_inst_yt_rsc_1_14_i_q_d,
      yt_rsc_1_15_i_q_d => peaseNTT_core_inst_yt_rsc_1_15_i_q_d,
      yt_rsc_1_16_i_clkr_en_d => yt_rsc_1_16_i_clkr_en_d,
      yt_rsc_1_16_i_q_d => peaseNTT_core_inst_yt_rsc_1_16_i_q_d,
      yt_rsc_1_17_i_q_d => peaseNTT_core_inst_yt_rsc_1_17_i_q_d,
      yt_rsc_1_18_i_q_d => peaseNTT_core_inst_yt_rsc_1_18_i_q_d,
      yt_rsc_1_19_i_q_d => peaseNTT_core_inst_yt_rsc_1_19_i_q_d,
      yt_rsc_1_20_i_q_d => peaseNTT_core_inst_yt_rsc_1_20_i_q_d,
      yt_rsc_1_21_i_q_d => peaseNTT_core_inst_yt_rsc_1_21_i_q_d,
      yt_rsc_1_22_i_q_d => peaseNTT_core_inst_yt_rsc_1_22_i_q_d,
      yt_rsc_1_23_i_q_d => peaseNTT_core_inst_yt_rsc_1_23_i_q_d,
      yt_rsc_1_24_i_q_d => peaseNTT_core_inst_yt_rsc_1_24_i_q_d,
      yt_rsc_1_25_i_q_d => peaseNTT_core_inst_yt_rsc_1_25_i_q_d,
      yt_rsc_1_26_i_q_d => peaseNTT_core_inst_yt_rsc_1_26_i_q_d,
      yt_rsc_1_27_i_q_d => peaseNTT_core_inst_yt_rsc_1_27_i_q_d,
      yt_rsc_1_28_i_q_d => peaseNTT_core_inst_yt_rsc_1_28_i_q_d,
      yt_rsc_1_29_i_q_d => peaseNTT_core_inst_yt_rsc_1_29_i_q_d,
      yt_rsc_1_30_i_q_d => peaseNTT_core_inst_yt_rsc_1_30_i_q_d,
      yt_rsc_1_31_i_q_d => peaseNTT_core_inst_yt_rsc_1_31_i_q_d,
      yt_rsc_2_0_i_clkr_en_d => yt_rsc_2_0_i_clkr_en_d,
      yt_rsc_2_0_i_q_d => peaseNTT_core_inst_yt_rsc_2_0_i_q_d,
      yt_rsc_2_1_i_q_d => peaseNTT_core_inst_yt_rsc_2_1_i_q_d,
      yt_rsc_2_2_i_q_d => peaseNTT_core_inst_yt_rsc_2_2_i_q_d,
      yt_rsc_2_3_i_q_d => peaseNTT_core_inst_yt_rsc_2_3_i_q_d,
      yt_rsc_2_4_i_q_d => peaseNTT_core_inst_yt_rsc_2_4_i_q_d,
      yt_rsc_2_5_i_q_d => peaseNTT_core_inst_yt_rsc_2_5_i_q_d,
      yt_rsc_2_6_i_q_d => peaseNTT_core_inst_yt_rsc_2_6_i_q_d,
      yt_rsc_2_7_i_q_d => peaseNTT_core_inst_yt_rsc_2_7_i_q_d,
      yt_rsc_2_8_i_q_d => peaseNTT_core_inst_yt_rsc_2_8_i_q_d,
      yt_rsc_2_9_i_q_d => peaseNTT_core_inst_yt_rsc_2_9_i_q_d,
      yt_rsc_2_10_i_q_d => peaseNTT_core_inst_yt_rsc_2_10_i_q_d,
      yt_rsc_2_11_i_q_d => peaseNTT_core_inst_yt_rsc_2_11_i_q_d,
      yt_rsc_2_12_i_q_d => peaseNTT_core_inst_yt_rsc_2_12_i_q_d,
      yt_rsc_2_13_i_q_d => peaseNTT_core_inst_yt_rsc_2_13_i_q_d,
      yt_rsc_2_14_i_q_d => peaseNTT_core_inst_yt_rsc_2_14_i_q_d,
      yt_rsc_2_15_i_q_d => peaseNTT_core_inst_yt_rsc_2_15_i_q_d,
      yt_rsc_2_16_i_clkr_en_d => yt_rsc_2_16_i_clkr_en_d,
      yt_rsc_2_16_i_q_d => peaseNTT_core_inst_yt_rsc_2_16_i_q_d,
      yt_rsc_2_17_i_q_d => peaseNTT_core_inst_yt_rsc_2_17_i_q_d,
      yt_rsc_2_18_i_q_d => peaseNTT_core_inst_yt_rsc_2_18_i_q_d,
      yt_rsc_2_19_i_q_d => peaseNTT_core_inst_yt_rsc_2_19_i_q_d,
      yt_rsc_2_20_i_q_d => peaseNTT_core_inst_yt_rsc_2_20_i_q_d,
      yt_rsc_2_21_i_q_d => peaseNTT_core_inst_yt_rsc_2_21_i_q_d,
      yt_rsc_2_22_i_q_d => peaseNTT_core_inst_yt_rsc_2_22_i_q_d,
      yt_rsc_2_23_i_q_d => peaseNTT_core_inst_yt_rsc_2_23_i_q_d,
      yt_rsc_2_24_i_q_d => peaseNTT_core_inst_yt_rsc_2_24_i_q_d,
      yt_rsc_2_25_i_q_d => peaseNTT_core_inst_yt_rsc_2_25_i_q_d,
      yt_rsc_2_26_i_q_d => peaseNTT_core_inst_yt_rsc_2_26_i_q_d,
      yt_rsc_2_27_i_q_d => peaseNTT_core_inst_yt_rsc_2_27_i_q_d,
      yt_rsc_2_28_i_q_d => peaseNTT_core_inst_yt_rsc_2_28_i_q_d,
      yt_rsc_2_29_i_q_d => peaseNTT_core_inst_yt_rsc_2_29_i_q_d,
      yt_rsc_2_30_i_q_d => peaseNTT_core_inst_yt_rsc_2_30_i_q_d,
      yt_rsc_2_31_i_q_d => peaseNTT_core_inst_yt_rsc_2_31_i_q_d,
      yt_rsc_3_0_i_clkr_en_d => yt_rsc_3_0_i_clkr_en_d,
      yt_rsc_3_0_i_q_d => peaseNTT_core_inst_yt_rsc_3_0_i_q_d,
      yt_rsc_3_1_i_q_d => peaseNTT_core_inst_yt_rsc_3_1_i_q_d,
      yt_rsc_3_2_i_q_d => peaseNTT_core_inst_yt_rsc_3_2_i_q_d,
      yt_rsc_3_3_i_q_d => peaseNTT_core_inst_yt_rsc_3_3_i_q_d,
      yt_rsc_3_4_i_q_d => peaseNTT_core_inst_yt_rsc_3_4_i_q_d,
      yt_rsc_3_5_i_q_d => peaseNTT_core_inst_yt_rsc_3_5_i_q_d,
      yt_rsc_3_6_i_q_d => peaseNTT_core_inst_yt_rsc_3_6_i_q_d,
      yt_rsc_3_7_i_q_d => peaseNTT_core_inst_yt_rsc_3_7_i_q_d,
      yt_rsc_3_8_i_q_d => peaseNTT_core_inst_yt_rsc_3_8_i_q_d,
      yt_rsc_3_9_i_q_d => peaseNTT_core_inst_yt_rsc_3_9_i_q_d,
      yt_rsc_3_10_i_q_d => peaseNTT_core_inst_yt_rsc_3_10_i_q_d,
      yt_rsc_3_11_i_q_d => peaseNTT_core_inst_yt_rsc_3_11_i_q_d,
      yt_rsc_3_12_i_q_d => peaseNTT_core_inst_yt_rsc_3_12_i_q_d,
      yt_rsc_3_13_i_q_d => peaseNTT_core_inst_yt_rsc_3_13_i_q_d,
      yt_rsc_3_14_i_q_d => peaseNTT_core_inst_yt_rsc_3_14_i_q_d,
      yt_rsc_3_15_i_q_d => peaseNTT_core_inst_yt_rsc_3_15_i_q_d,
      yt_rsc_3_16_i_clkr_en_d => yt_rsc_3_16_i_clkr_en_d,
      yt_rsc_3_16_i_q_d => peaseNTT_core_inst_yt_rsc_3_16_i_q_d,
      yt_rsc_3_17_i_q_d => peaseNTT_core_inst_yt_rsc_3_17_i_q_d,
      yt_rsc_3_18_i_q_d => peaseNTT_core_inst_yt_rsc_3_18_i_q_d,
      yt_rsc_3_19_i_q_d => peaseNTT_core_inst_yt_rsc_3_19_i_q_d,
      yt_rsc_3_20_i_q_d => peaseNTT_core_inst_yt_rsc_3_20_i_q_d,
      yt_rsc_3_21_i_q_d => peaseNTT_core_inst_yt_rsc_3_21_i_q_d,
      yt_rsc_3_22_i_q_d => peaseNTT_core_inst_yt_rsc_3_22_i_q_d,
      yt_rsc_3_23_i_q_d => peaseNTT_core_inst_yt_rsc_3_23_i_q_d,
      yt_rsc_3_24_i_q_d => peaseNTT_core_inst_yt_rsc_3_24_i_q_d,
      yt_rsc_3_25_i_q_d => peaseNTT_core_inst_yt_rsc_3_25_i_q_d,
      yt_rsc_3_26_i_q_d => peaseNTT_core_inst_yt_rsc_3_26_i_q_d,
      yt_rsc_3_27_i_q_d => peaseNTT_core_inst_yt_rsc_3_27_i_q_d,
      yt_rsc_3_28_i_q_d => peaseNTT_core_inst_yt_rsc_3_28_i_q_d,
      yt_rsc_3_29_i_q_d => peaseNTT_core_inst_yt_rsc_3_29_i_q_d,
      yt_rsc_3_30_i_q_d => peaseNTT_core_inst_yt_rsc_3_30_i_q_d,
      yt_rsc_3_31_i_q_d => peaseNTT_core_inst_yt_rsc_3_31_i_q_d,
      yt_rsc_4_0_i_clkr_en_d => yt_rsc_4_0_i_clkr_en_d,
      yt_rsc_4_0_i_q_d => peaseNTT_core_inst_yt_rsc_4_0_i_q_d,
      yt_rsc_4_1_i_q_d => peaseNTT_core_inst_yt_rsc_4_1_i_q_d,
      yt_rsc_4_2_i_q_d => peaseNTT_core_inst_yt_rsc_4_2_i_q_d,
      yt_rsc_4_3_i_q_d => peaseNTT_core_inst_yt_rsc_4_3_i_q_d,
      yt_rsc_4_4_i_q_d => peaseNTT_core_inst_yt_rsc_4_4_i_q_d,
      yt_rsc_4_5_i_q_d => peaseNTT_core_inst_yt_rsc_4_5_i_q_d,
      yt_rsc_4_6_i_q_d => peaseNTT_core_inst_yt_rsc_4_6_i_q_d,
      yt_rsc_4_7_i_q_d => peaseNTT_core_inst_yt_rsc_4_7_i_q_d,
      yt_rsc_4_8_i_q_d => peaseNTT_core_inst_yt_rsc_4_8_i_q_d,
      yt_rsc_4_9_i_q_d => peaseNTT_core_inst_yt_rsc_4_9_i_q_d,
      yt_rsc_4_10_i_q_d => peaseNTT_core_inst_yt_rsc_4_10_i_q_d,
      yt_rsc_4_11_i_q_d => peaseNTT_core_inst_yt_rsc_4_11_i_q_d,
      yt_rsc_4_12_i_q_d => peaseNTT_core_inst_yt_rsc_4_12_i_q_d,
      yt_rsc_4_13_i_q_d => peaseNTT_core_inst_yt_rsc_4_13_i_q_d,
      yt_rsc_4_14_i_q_d => peaseNTT_core_inst_yt_rsc_4_14_i_q_d,
      yt_rsc_4_15_i_q_d => peaseNTT_core_inst_yt_rsc_4_15_i_q_d,
      yt_rsc_4_16_i_clkr_en_d => yt_rsc_4_16_i_clkr_en_d,
      yt_rsc_4_16_i_q_d => peaseNTT_core_inst_yt_rsc_4_16_i_q_d,
      yt_rsc_4_17_i_q_d => peaseNTT_core_inst_yt_rsc_4_17_i_q_d,
      yt_rsc_4_18_i_q_d => peaseNTT_core_inst_yt_rsc_4_18_i_q_d,
      yt_rsc_4_19_i_q_d => peaseNTT_core_inst_yt_rsc_4_19_i_q_d,
      yt_rsc_4_20_i_q_d => peaseNTT_core_inst_yt_rsc_4_20_i_q_d,
      yt_rsc_4_21_i_q_d => peaseNTT_core_inst_yt_rsc_4_21_i_q_d,
      yt_rsc_4_22_i_q_d => peaseNTT_core_inst_yt_rsc_4_22_i_q_d,
      yt_rsc_4_23_i_q_d => peaseNTT_core_inst_yt_rsc_4_23_i_q_d,
      yt_rsc_4_24_i_q_d => peaseNTT_core_inst_yt_rsc_4_24_i_q_d,
      yt_rsc_4_25_i_q_d => peaseNTT_core_inst_yt_rsc_4_25_i_q_d,
      yt_rsc_4_26_i_q_d => peaseNTT_core_inst_yt_rsc_4_26_i_q_d,
      yt_rsc_4_27_i_q_d => peaseNTT_core_inst_yt_rsc_4_27_i_q_d,
      yt_rsc_4_28_i_q_d => peaseNTT_core_inst_yt_rsc_4_28_i_q_d,
      yt_rsc_4_29_i_q_d => peaseNTT_core_inst_yt_rsc_4_29_i_q_d,
      yt_rsc_4_30_i_q_d => peaseNTT_core_inst_yt_rsc_4_30_i_q_d,
      yt_rsc_4_31_i_q_d => peaseNTT_core_inst_yt_rsc_4_31_i_q_d,
      yt_rsc_5_0_i_clkr_en_d => yt_rsc_5_0_i_clkr_en_d,
      yt_rsc_5_0_i_q_d => peaseNTT_core_inst_yt_rsc_5_0_i_q_d,
      yt_rsc_5_1_i_q_d => peaseNTT_core_inst_yt_rsc_5_1_i_q_d,
      yt_rsc_5_2_i_q_d => peaseNTT_core_inst_yt_rsc_5_2_i_q_d,
      yt_rsc_5_3_i_q_d => peaseNTT_core_inst_yt_rsc_5_3_i_q_d,
      yt_rsc_5_4_i_q_d => peaseNTT_core_inst_yt_rsc_5_4_i_q_d,
      yt_rsc_5_5_i_q_d => peaseNTT_core_inst_yt_rsc_5_5_i_q_d,
      yt_rsc_5_6_i_q_d => peaseNTT_core_inst_yt_rsc_5_6_i_q_d,
      yt_rsc_5_7_i_q_d => peaseNTT_core_inst_yt_rsc_5_7_i_q_d,
      yt_rsc_5_8_i_q_d => peaseNTT_core_inst_yt_rsc_5_8_i_q_d,
      yt_rsc_5_9_i_q_d => peaseNTT_core_inst_yt_rsc_5_9_i_q_d,
      yt_rsc_5_10_i_q_d => peaseNTT_core_inst_yt_rsc_5_10_i_q_d,
      yt_rsc_5_11_i_q_d => peaseNTT_core_inst_yt_rsc_5_11_i_q_d,
      yt_rsc_5_12_i_q_d => peaseNTT_core_inst_yt_rsc_5_12_i_q_d,
      yt_rsc_5_13_i_q_d => peaseNTT_core_inst_yt_rsc_5_13_i_q_d,
      yt_rsc_5_14_i_q_d => peaseNTT_core_inst_yt_rsc_5_14_i_q_d,
      yt_rsc_5_15_i_q_d => peaseNTT_core_inst_yt_rsc_5_15_i_q_d,
      yt_rsc_5_16_i_clkr_en_d => yt_rsc_5_16_i_clkr_en_d,
      yt_rsc_5_16_i_q_d => peaseNTT_core_inst_yt_rsc_5_16_i_q_d,
      yt_rsc_5_17_i_q_d => peaseNTT_core_inst_yt_rsc_5_17_i_q_d,
      yt_rsc_5_18_i_q_d => peaseNTT_core_inst_yt_rsc_5_18_i_q_d,
      yt_rsc_5_19_i_q_d => peaseNTT_core_inst_yt_rsc_5_19_i_q_d,
      yt_rsc_5_20_i_q_d => peaseNTT_core_inst_yt_rsc_5_20_i_q_d,
      yt_rsc_5_21_i_q_d => peaseNTT_core_inst_yt_rsc_5_21_i_q_d,
      yt_rsc_5_22_i_q_d => peaseNTT_core_inst_yt_rsc_5_22_i_q_d,
      yt_rsc_5_23_i_q_d => peaseNTT_core_inst_yt_rsc_5_23_i_q_d,
      yt_rsc_5_24_i_q_d => peaseNTT_core_inst_yt_rsc_5_24_i_q_d,
      yt_rsc_5_25_i_q_d => peaseNTT_core_inst_yt_rsc_5_25_i_q_d,
      yt_rsc_5_26_i_q_d => peaseNTT_core_inst_yt_rsc_5_26_i_q_d,
      yt_rsc_5_27_i_q_d => peaseNTT_core_inst_yt_rsc_5_27_i_q_d,
      yt_rsc_5_28_i_q_d => peaseNTT_core_inst_yt_rsc_5_28_i_q_d,
      yt_rsc_5_29_i_q_d => peaseNTT_core_inst_yt_rsc_5_29_i_q_d,
      yt_rsc_5_30_i_q_d => peaseNTT_core_inst_yt_rsc_5_30_i_q_d,
      yt_rsc_5_31_i_q_d => peaseNTT_core_inst_yt_rsc_5_31_i_q_d,
      yt_rsc_6_0_i_clkr_en_d => yt_rsc_6_0_i_clkr_en_d,
      yt_rsc_6_0_i_q_d => peaseNTT_core_inst_yt_rsc_6_0_i_q_d,
      yt_rsc_6_1_i_q_d => peaseNTT_core_inst_yt_rsc_6_1_i_q_d,
      yt_rsc_6_2_i_q_d => peaseNTT_core_inst_yt_rsc_6_2_i_q_d,
      yt_rsc_6_3_i_q_d => peaseNTT_core_inst_yt_rsc_6_3_i_q_d,
      yt_rsc_6_4_i_q_d => peaseNTT_core_inst_yt_rsc_6_4_i_q_d,
      yt_rsc_6_5_i_q_d => peaseNTT_core_inst_yt_rsc_6_5_i_q_d,
      yt_rsc_6_6_i_q_d => peaseNTT_core_inst_yt_rsc_6_6_i_q_d,
      yt_rsc_6_7_i_q_d => peaseNTT_core_inst_yt_rsc_6_7_i_q_d,
      yt_rsc_6_8_i_q_d => peaseNTT_core_inst_yt_rsc_6_8_i_q_d,
      yt_rsc_6_9_i_q_d => peaseNTT_core_inst_yt_rsc_6_9_i_q_d,
      yt_rsc_6_10_i_q_d => peaseNTT_core_inst_yt_rsc_6_10_i_q_d,
      yt_rsc_6_11_i_q_d => peaseNTT_core_inst_yt_rsc_6_11_i_q_d,
      yt_rsc_6_12_i_q_d => peaseNTT_core_inst_yt_rsc_6_12_i_q_d,
      yt_rsc_6_13_i_q_d => peaseNTT_core_inst_yt_rsc_6_13_i_q_d,
      yt_rsc_6_14_i_q_d => peaseNTT_core_inst_yt_rsc_6_14_i_q_d,
      yt_rsc_6_15_i_q_d => peaseNTT_core_inst_yt_rsc_6_15_i_q_d,
      yt_rsc_6_16_i_clkr_en_d => yt_rsc_6_16_i_clkr_en_d,
      yt_rsc_6_16_i_q_d => peaseNTT_core_inst_yt_rsc_6_16_i_q_d,
      yt_rsc_6_17_i_q_d => peaseNTT_core_inst_yt_rsc_6_17_i_q_d,
      yt_rsc_6_18_i_q_d => peaseNTT_core_inst_yt_rsc_6_18_i_q_d,
      yt_rsc_6_19_i_q_d => peaseNTT_core_inst_yt_rsc_6_19_i_q_d,
      yt_rsc_6_20_i_q_d => peaseNTT_core_inst_yt_rsc_6_20_i_q_d,
      yt_rsc_6_21_i_q_d => peaseNTT_core_inst_yt_rsc_6_21_i_q_d,
      yt_rsc_6_22_i_q_d => peaseNTT_core_inst_yt_rsc_6_22_i_q_d,
      yt_rsc_6_23_i_q_d => peaseNTT_core_inst_yt_rsc_6_23_i_q_d,
      yt_rsc_6_24_i_q_d => peaseNTT_core_inst_yt_rsc_6_24_i_q_d,
      yt_rsc_6_25_i_q_d => peaseNTT_core_inst_yt_rsc_6_25_i_q_d,
      yt_rsc_6_26_i_q_d => peaseNTT_core_inst_yt_rsc_6_26_i_q_d,
      yt_rsc_6_27_i_q_d => peaseNTT_core_inst_yt_rsc_6_27_i_q_d,
      yt_rsc_6_28_i_q_d => peaseNTT_core_inst_yt_rsc_6_28_i_q_d,
      yt_rsc_6_29_i_q_d => peaseNTT_core_inst_yt_rsc_6_29_i_q_d,
      yt_rsc_6_30_i_q_d => peaseNTT_core_inst_yt_rsc_6_30_i_q_d,
      yt_rsc_6_31_i_q_d => peaseNTT_core_inst_yt_rsc_6_31_i_q_d,
      yt_rsc_7_0_i_clkr_en_d => yt_rsc_7_0_i_clkr_en_d,
      yt_rsc_7_0_i_q_d => peaseNTT_core_inst_yt_rsc_7_0_i_q_d,
      yt_rsc_7_1_i_q_d => peaseNTT_core_inst_yt_rsc_7_1_i_q_d,
      yt_rsc_7_2_i_q_d => peaseNTT_core_inst_yt_rsc_7_2_i_q_d,
      yt_rsc_7_3_i_q_d => peaseNTT_core_inst_yt_rsc_7_3_i_q_d,
      yt_rsc_7_4_i_q_d => peaseNTT_core_inst_yt_rsc_7_4_i_q_d,
      yt_rsc_7_5_i_q_d => peaseNTT_core_inst_yt_rsc_7_5_i_q_d,
      yt_rsc_7_6_i_q_d => peaseNTT_core_inst_yt_rsc_7_6_i_q_d,
      yt_rsc_7_7_i_q_d => peaseNTT_core_inst_yt_rsc_7_7_i_q_d,
      yt_rsc_7_8_i_q_d => peaseNTT_core_inst_yt_rsc_7_8_i_q_d,
      yt_rsc_7_9_i_q_d => peaseNTT_core_inst_yt_rsc_7_9_i_q_d,
      yt_rsc_7_10_i_q_d => peaseNTT_core_inst_yt_rsc_7_10_i_q_d,
      yt_rsc_7_11_i_q_d => peaseNTT_core_inst_yt_rsc_7_11_i_q_d,
      yt_rsc_7_12_i_q_d => peaseNTT_core_inst_yt_rsc_7_12_i_q_d,
      yt_rsc_7_13_i_q_d => peaseNTT_core_inst_yt_rsc_7_13_i_q_d,
      yt_rsc_7_14_i_q_d => peaseNTT_core_inst_yt_rsc_7_14_i_q_d,
      yt_rsc_7_15_i_q_d => peaseNTT_core_inst_yt_rsc_7_15_i_q_d,
      yt_rsc_7_16_i_clkr_en_d => yt_rsc_7_16_i_clkr_en_d,
      yt_rsc_7_16_i_q_d => peaseNTT_core_inst_yt_rsc_7_16_i_q_d,
      yt_rsc_7_17_i_q_d => peaseNTT_core_inst_yt_rsc_7_17_i_q_d,
      yt_rsc_7_18_i_q_d => peaseNTT_core_inst_yt_rsc_7_18_i_q_d,
      yt_rsc_7_19_i_q_d => peaseNTT_core_inst_yt_rsc_7_19_i_q_d,
      yt_rsc_7_20_i_q_d => peaseNTT_core_inst_yt_rsc_7_20_i_q_d,
      yt_rsc_7_21_i_q_d => peaseNTT_core_inst_yt_rsc_7_21_i_q_d,
      yt_rsc_7_22_i_q_d => peaseNTT_core_inst_yt_rsc_7_22_i_q_d,
      yt_rsc_7_23_i_q_d => peaseNTT_core_inst_yt_rsc_7_23_i_q_d,
      yt_rsc_7_24_i_q_d => peaseNTT_core_inst_yt_rsc_7_24_i_q_d,
      yt_rsc_7_25_i_q_d => peaseNTT_core_inst_yt_rsc_7_25_i_q_d,
      yt_rsc_7_26_i_q_d => peaseNTT_core_inst_yt_rsc_7_26_i_q_d,
      yt_rsc_7_27_i_q_d => peaseNTT_core_inst_yt_rsc_7_27_i_q_d,
      yt_rsc_7_28_i_q_d => peaseNTT_core_inst_yt_rsc_7_28_i_q_d,
      yt_rsc_7_29_i_q_d => peaseNTT_core_inst_yt_rsc_7_29_i_q_d,
      yt_rsc_7_30_i_q_d => peaseNTT_core_inst_yt_rsc_7_30_i_q_d,
      yt_rsc_7_31_i_q_d => peaseNTT_core_inst_yt_rsc_7_31_i_q_d,
      xt_rsc_0_0_i_qa_d => peaseNTT_core_inst_xt_rsc_0_0_i_qa_d,
      xt_rsc_0_1_i_qa_d => peaseNTT_core_inst_xt_rsc_0_1_i_qa_d,
      xt_rsc_0_2_i_qa_d => peaseNTT_core_inst_xt_rsc_0_2_i_qa_d,
      xt_rsc_0_3_i_qa_d => peaseNTT_core_inst_xt_rsc_0_3_i_qa_d,
      xt_rsc_0_4_i_qa_d => peaseNTT_core_inst_xt_rsc_0_4_i_qa_d,
      xt_rsc_0_5_i_qa_d => peaseNTT_core_inst_xt_rsc_0_5_i_qa_d,
      xt_rsc_0_6_i_qa_d => peaseNTT_core_inst_xt_rsc_0_6_i_qa_d,
      xt_rsc_0_7_i_qa_d => peaseNTT_core_inst_xt_rsc_0_7_i_qa_d,
      xt_rsc_0_8_i_qa_d => peaseNTT_core_inst_xt_rsc_0_8_i_qa_d,
      xt_rsc_0_9_i_qa_d => peaseNTT_core_inst_xt_rsc_0_9_i_qa_d,
      xt_rsc_0_10_i_qa_d => peaseNTT_core_inst_xt_rsc_0_10_i_qa_d,
      xt_rsc_0_11_i_qa_d => peaseNTT_core_inst_xt_rsc_0_11_i_qa_d,
      xt_rsc_0_12_i_qa_d => peaseNTT_core_inst_xt_rsc_0_12_i_qa_d,
      xt_rsc_0_13_i_qa_d => peaseNTT_core_inst_xt_rsc_0_13_i_qa_d,
      xt_rsc_0_14_i_qa_d => peaseNTT_core_inst_xt_rsc_0_14_i_qa_d,
      xt_rsc_0_15_i_qa_d => peaseNTT_core_inst_xt_rsc_0_15_i_qa_d,
      xt_rsc_0_16_i_qa_d => peaseNTT_core_inst_xt_rsc_0_16_i_qa_d,
      xt_rsc_0_17_i_qa_d => peaseNTT_core_inst_xt_rsc_0_17_i_qa_d,
      xt_rsc_0_18_i_qa_d => peaseNTT_core_inst_xt_rsc_0_18_i_qa_d,
      xt_rsc_0_19_i_qa_d => peaseNTT_core_inst_xt_rsc_0_19_i_qa_d,
      xt_rsc_0_20_i_qa_d => peaseNTT_core_inst_xt_rsc_0_20_i_qa_d,
      xt_rsc_0_21_i_qa_d => peaseNTT_core_inst_xt_rsc_0_21_i_qa_d,
      xt_rsc_0_22_i_qa_d => peaseNTT_core_inst_xt_rsc_0_22_i_qa_d,
      xt_rsc_0_23_i_qa_d => peaseNTT_core_inst_xt_rsc_0_23_i_qa_d,
      xt_rsc_0_24_i_qa_d => peaseNTT_core_inst_xt_rsc_0_24_i_qa_d,
      xt_rsc_0_25_i_qa_d => peaseNTT_core_inst_xt_rsc_0_25_i_qa_d,
      xt_rsc_0_26_i_qa_d => peaseNTT_core_inst_xt_rsc_0_26_i_qa_d,
      xt_rsc_0_27_i_qa_d => peaseNTT_core_inst_xt_rsc_0_27_i_qa_d,
      xt_rsc_0_28_i_qa_d => peaseNTT_core_inst_xt_rsc_0_28_i_qa_d,
      xt_rsc_0_29_i_qa_d => peaseNTT_core_inst_xt_rsc_0_29_i_qa_d,
      xt_rsc_0_30_i_qa_d => peaseNTT_core_inst_xt_rsc_0_30_i_qa_d,
      xt_rsc_0_31_i_qa_d => peaseNTT_core_inst_xt_rsc_0_31_i_qa_d,
      xt_rsc_1_0_i_qa_d => peaseNTT_core_inst_xt_rsc_1_0_i_qa_d,
      xt_rsc_1_1_i_qa_d => peaseNTT_core_inst_xt_rsc_1_1_i_qa_d,
      xt_rsc_1_2_i_qa_d => peaseNTT_core_inst_xt_rsc_1_2_i_qa_d,
      xt_rsc_1_3_i_qa_d => peaseNTT_core_inst_xt_rsc_1_3_i_qa_d,
      xt_rsc_1_4_i_qa_d => peaseNTT_core_inst_xt_rsc_1_4_i_qa_d,
      xt_rsc_1_5_i_qa_d => peaseNTT_core_inst_xt_rsc_1_5_i_qa_d,
      xt_rsc_1_6_i_qa_d => peaseNTT_core_inst_xt_rsc_1_6_i_qa_d,
      xt_rsc_1_7_i_qa_d => peaseNTT_core_inst_xt_rsc_1_7_i_qa_d,
      xt_rsc_1_8_i_qa_d => peaseNTT_core_inst_xt_rsc_1_8_i_qa_d,
      xt_rsc_1_9_i_qa_d => peaseNTT_core_inst_xt_rsc_1_9_i_qa_d,
      xt_rsc_1_10_i_qa_d => peaseNTT_core_inst_xt_rsc_1_10_i_qa_d,
      xt_rsc_1_11_i_qa_d => peaseNTT_core_inst_xt_rsc_1_11_i_qa_d,
      xt_rsc_1_12_i_qa_d => peaseNTT_core_inst_xt_rsc_1_12_i_qa_d,
      xt_rsc_1_13_i_qa_d => peaseNTT_core_inst_xt_rsc_1_13_i_qa_d,
      xt_rsc_1_14_i_qa_d => peaseNTT_core_inst_xt_rsc_1_14_i_qa_d,
      xt_rsc_1_15_i_qa_d => peaseNTT_core_inst_xt_rsc_1_15_i_qa_d,
      xt_rsc_1_16_i_qa_d => peaseNTT_core_inst_xt_rsc_1_16_i_qa_d,
      xt_rsc_1_17_i_qa_d => peaseNTT_core_inst_xt_rsc_1_17_i_qa_d,
      xt_rsc_1_18_i_qa_d => peaseNTT_core_inst_xt_rsc_1_18_i_qa_d,
      xt_rsc_1_19_i_qa_d => peaseNTT_core_inst_xt_rsc_1_19_i_qa_d,
      xt_rsc_1_20_i_qa_d => peaseNTT_core_inst_xt_rsc_1_20_i_qa_d,
      xt_rsc_1_21_i_qa_d => peaseNTT_core_inst_xt_rsc_1_21_i_qa_d,
      xt_rsc_1_22_i_qa_d => peaseNTT_core_inst_xt_rsc_1_22_i_qa_d,
      xt_rsc_1_23_i_qa_d => peaseNTT_core_inst_xt_rsc_1_23_i_qa_d,
      xt_rsc_1_24_i_qa_d => peaseNTT_core_inst_xt_rsc_1_24_i_qa_d,
      xt_rsc_1_25_i_qa_d => peaseNTT_core_inst_xt_rsc_1_25_i_qa_d,
      xt_rsc_1_26_i_qa_d => peaseNTT_core_inst_xt_rsc_1_26_i_qa_d,
      xt_rsc_1_27_i_qa_d => peaseNTT_core_inst_xt_rsc_1_27_i_qa_d,
      xt_rsc_1_28_i_qa_d => peaseNTT_core_inst_xt_rsc_1_28_i_qa_d,
      xt_rsc_1_29_i_qa_d => peaseNTT_core_inst_xt_rsc_1_29_i_qa_d,
      xt_rsc_1_30_i_qa_d => peaseNTT_core_inst_xt_rsc_1_30_i_qa_d,
      xt_rsc_1_31_i_qa_d => peaseNTT_core_inst_xt_rsc_1_31_i_qa_d,
      xt_rsc_2_0_i_qa_d => peaseNTT_core_inst_xt_rsc_2_0_i_qa_d,
      xt_rsc_2_1_i_qa_d => peaseNTT_core_inst_xt_rsc_2_1_i_qa_d,
      xt_rsc_2_2_i_qa_d => peaseNTT_core_inst_xt_rsc_2_2_i_qa_d,
      xt_rsc_2_3_i_qa_d => peaseNTT_core_inst_xt_rsc_2_3_i_qa_d,
      xt_rsc_2_4_i_qa_d => peaseNTT_core_inst_xt_rsc_2_4_i_qa_d,
      xt_rsc_2_5_i_qa_d => peaseNTT_core_inst_xt_rsc_2_5_i_qa_d,
      xt_rsc_2_6_i_qa_d => peaseNTT_core_inst_xt_rsc_2_6_i_qa_d,
      xt_rsc_2_7_i_qa_d => peaseNTT_core_inst_xt_rsc_2_7_i_qa_d,
      xt_rsc_2_8_i_qa_d => peaseNTT_core_inst_xt_rsc_2_8_i_qa_d,
      xt_rsc_2_9_i_qa_d => peaseNTT_core_inst_xt_rsc_2_9_i_qa_d,
      xt_rsc_2_10_i_qa_d => peaseNTT_core_inst_xt_rsc_2_10_i_qa_d,
      xt_rsc_2_11_i_qa_d => peaseNTT_core_inst_xt_rsc_2_11_i_qa_d,
      xt_rsc_2_12_i_qa_d => peaseNTT_core_inst_xt_rsc_2_12_i_qa_d,
      xt_rsc_2_13_i_qa_d => peaseNTT_core_inst_xt_rsc_2_13_i_qa_d,
      xt_rsc_2_14_i_qa_d => peaseNTT_core_inst_xt_rsc_2_14_i_qa_d,
      xt_rsc_2_15_i_qa_d => peaseNTT_core_inst_xt_rsc_2_15_i_qa_d,
      xt_rsc_2_16_i_qa_d => peaseNTT_core_inst_xt_rsc_2_16_i_qa_d,
      xt_rsc_2_17_i_qa_d => peaseNTT_core_inst_xt_rsc_2_17_i_qa_d,
      xt_rsc_2_18_i_qa_d => peaseNTT_core_inst_xt_rsc_2_18_i_qa_d,
      xt_rsc_2_19_i_qa_d => peaseNTT_core_inst_xt_rsc_2_19_i_qa_d,
      xt_rsc_2_20_i_qa_d => peaseNTT_core_inst_xt_rsc_2_20_i_qa_d,
      xt_rsc_2_21_i_qa_d => peaseNTT_core_inst_xt_rsc_2_21_i_qa_d,
      xt_rsc_2_22_i_qa_d => peaseNTT_core_inst_xt_rsc_2_22_i_qa_d,
      xt_rsc_2_23_i_qa_d => peaseNTT_core_inst_xt_rsc_2_23_i_qa_d,
      xt_rsc_2_24_i_qa_d => peaseNTT_core_inst_xt_rsc_2_24_i_qa_d,
      xt_rsc_2_25_i_qa_d => peaseNTT_core_inst_xt_rsc_2_25_i_qa_d,
      xt_rsc_2_26_i_qa_d => peaseNTT_core_inst_xt_rsc_2_26_i_qa_d,
      xt_rsc_2_27_i_qa_d => peaseNTT_core_inst_xt_rsc_2_27_i_qa_d,
      xt_rsc_2_28_i_qa_d => peaseNTT_core_inst_xt_rsc_2_28_i_qa_d,
      xt_rsc_2_29_i_qa_d => peaseNTT_core_inst_xt_rsc_2_29_i_qa_d,
      xt_rsc_2_30_i_qa_d => peaseNTT_core_inst_xt_rsc_2_30_i_qa_d,
      xt_rsc_2_31_i_qa_d => peaseNTT_core_inst_xt_rsc_2_31_i_qa_d,
      xt_rsc_3_0_i_qa_d => peaseNTT_core_inst_xt_rsc_3_0_i_qa_d,
      xt_rsc_3_1_i_qa_d => peaseNTT_core_inst_xt_rsc_3_1_i_qa_d,
      xt_rsc_3_2_i_qa_d => peaseNTT_core_inst_xt_rsc_3_2_i_qa_d,
      xt_rsc_3_3_i_qa_d => peaseNTT_core_inst_xt_rsc_3_3_i_qa_d,
      xt_rsc_3_4_i_qa_d => peaseNTT_core_inst_xt_rsc_3_4_i_qa_d,
      xt_rsc_3_5_i_qa_d => peaseNTT_core_inst_xt_rsc_3_5_i_qa_d,
      xt_rsc_3_6_i_qa_d => peaseNTT_core_inst_xt_rsc_3_6_i_qa_d,
      xt_rsc_3_7_i_qa_d => peaseNTT_core_inst_xt_rsc_3_7_i_qa_d,
      xt_rsc_3_8_i_qa_d => peaseNTT_core_inst_xt_rsc_3_8_i_qa_d,
      xt_rsc_3_9_i_qa_d => peaseNTT_core_inst_xt_rsc_3_9_i_qa_d,
      xt_rsc_3_10_i_qa_d => peaseNTT_core_inst_xt_rsc_3_10_i_qa_d,
      xt_rsc_3_11_i_qa_d => peaseNTT_core_inst_xt_rsc_3_11_i_qa_d,
      xt_rsc_3_12_i_qa_d => peaseNTT_core_inst_xt_rsc_3_12_i_qa_d,
      xt_rsc_3_13_i_qa_d => peaseNTT_core_inst_xt_rsc_3_13_i_qa_d,
      xt_rsc_3_14_i_qa_d => peaseNTT_core_inst_xt_rsc_3_14_i_qa_d,
      xt_rsc_3_15_i_qa_d => peaseNTT_core_inst_xt_rsc_3_15_i_qa_d,
      xt_rsc_3_16_i_qa_d => peaseNTT_core_inst_xt_rsc_3_16_i_qa_d,
      xt_rsc_3_17_i_qa_d => peaseNTT_core_inst_xt_rsc_3_17_i_qa_d,
      xt_rsc_3_18_i_qa_d => peaseNTT_core_inst_xt_rsc_3_18_i_qa_d,
      xt_rsc_3_19_i_qa_d => peaseNTT_core_inst_xt_rsc_3_19_i_qa_d,
      xt_rsc_3_20_i_qa_d => peaseNTT_core_inst_xt_rsc_3_20_i_qa_d,
      xt_rsc_3_21_i_qa_d => peaseNTT_core_inst_xt_rsc_3_21_i_qa_d,
      xt_rsc_3_22_i_qa_d => peaseNTT_core_inst_xt_rsc_3_22_i_qa_d,
      xt_rsc_3_23_i_qa_d => peaseNTT_core_inst_xt_rsc_3_23_i_qa_d,
      xt_rsc_3_24_i_qa_d => peaseNTT_core_inst_xt_rsc_3_24_i_qa_d,
      xt_rsc_3_25_i_qa_d => peaseNTT_core_inst_xt_rsc_3_25_i_qa_d,
      xt_rsc_3_26_i_qa_d => peaseNTT_core_inst_xt_rsc_3_26_i_qa_d,
      xt_rsc_3_27_i_qa_d => peaseNTT_core_inst_xt_rsc_3_27_i_qa_d,
      xt_rsc_3_28_i_qa_d => peaseNTT_core_inst_xt_rsc_3_28_i_qa_d,
      xt_rsc_3_29_i_qa_d => peaseNTT_core_inst_xt_rsc_3_29_i_qa_d,
      xt_rsc_3_30_i_qa_d => peaseNTT_core_inst_xt_rsc_3_30_i_qa_d,
      xt_rsc_3_31_i_qa_d => peaseNTT_core_inst_xt_rsc_3_31_i_qa_d,
      xt_rsc_4_0_i_qa_d => peaseNTT_core_inst_xt_rsc_4_0_i_qa_d,
      xt_rsc_4_1_i_qa_d => peaseNTT_core_inst_xt_rsc_4_1_i_qa_d,
      xt_rsc_4_2_i_qa_d => peaseNTT_core_inst_xt_rsc_4_2_i_qa_d,
      xt_rsc_4_3_i_qa_d => peaseNTT_core_inst_xt_rsc_4_3_i_qa_d,
      xt_rsc_4_4_i_qa_d => peaseNTT_core_inst_xt_rsc_4_4_i_qa_d,
      xt_rsc_4_5_i_qa_d => peaseNTT_core_inst_xt_rsc_4_5_i_qa_d,
      xt_rsc_4_6_i_qa_d => peaseNTT_core_inst_xt_rsc_4_6_i_qa_d,
      xt_rsc_4_7_i_qa_d => peaseNTT_core_inst_xt_rsc_4_7_i_qa_d,
      xt_rsc_4_8_i_qa_d => peaseNTT_core_inst_xt_rsc_4_8_i_qa_d,
      xt_rsc_4_9_i_qa_d => peaseNTT_core_inst_xt_rsc_4_9_i_qa_d,
      xt_rsc_4_10_i_qa_d => peaseNTT_core_inst_xt_rsc_4_10_i_qa_d,
      xt_rsc_4_11_i_qa_d => peaseNTT_core_inst_xt_rsc_4_11_i_qa_d,
      xt_rsc_4_12_i_qa_d => peaseNTT_core_inst_xt_rsc_4_12_i_qa_d,
      xt_rsc_4_13_i_qa_d => peaseNTT_core_inst_xt_rsc_4_13_i_qa_d,
      xt_rsc_4_14_i_qa_d => peaseNTT_core_inst_xt_rsc_4_14_i_qa_d,
      xt_rsc_4_15_i_qa_d => peaseNTT_core_inst_xt_rsc_4_15_i_qa_d,
      xt_rsc_4_16_i_qa_d => peaseNTT_core_inst_xt_rsc_4_16_i_qa_d,
      xt_rsc_4_17_i_qa_d => peaseNTT_core_inst_xt_rsc_4_17_i_qa_d,
      xt_rsc_4_18_i_qa_d => peaseNTT_core_inst_xt_rsc_4_18_i_qa_d,
      xt_rsc_4_19_i_qa_d => peaseNTT_core_inst_xt_rsc_4_19_i_qa_d,
      xt_rsc_4_20_i_qa_d => peaseNTT_core_inst_xt_rsc_4_20_i_qa_d,
      xt_rsc_4_21_i_qa_d => peaseNTT_core_inst_xt_rsc_4_21_i_qa_d,
      xt_rsc_4_22_i_qa_d => peaseNTT_core_inst_xt_rsc_4_22_i_qa_d,
      xt_rsc_4_23_i_qa_d => peaseNTT_core_inst_xt_rsc_4_23_i_qa_d,
      xt_rsc_4_24_i_qa_d => peaseNTT_core_inst_xt_rsc_4_24_i_qa_d,
      xt_rsc_4_25_i_qa_d => peaseNTT_core_inst_xt_rsc_4_25_i_qa_d,
      xt_rsc_4_26_i_qa_d => peaseNTT_core_inst_xt_rsc_4_26_i_qa_d,
      xt_rsc_4_27_i_qa_d => peaseNTT_core_inst_xt_rsc_4_27_i_qa_d,
      xt_rsc_4_28_i_qa_d => peaseNTT_core_inst_xt_rsc_4_28_i_qa_d,
      xt_rsc_4_29_i_qa_d => peaseNTT_core_inst_xt_rsc_4_29_i_qa_d,
      xt_rsc_4_30_i_qa_d => peaseNTT_core_inst_xt_rsc_4_30_i_qa_d,
      xt_rsc_4_31_i_qa_d => peaseNTT_core_inst_xt_rsc_4_31_i_qa_d,
      xt_rsc_5_0_i_qa_d => peaseNTT_core_inst_xt_rsc_5_0_i_qa_d,
      xt_rsc_5_1_i_qa_d => peaseNTT_core_inst_xt_rsc_5_1_i_qa_d,
      xt_rsc_5_2_i_qa_d => peaseNTT_core_inst_xt_rsc_5_2_i_qa_d,
      xt_rsc_5_3_i_qa_d => peaseNTT_core_inst_xt_rsc_5_3_i_qa_d,
      xt_rsc_5_4_i_qa_d => peaseNTT_core_inst_xt_rsc_5_4_i_qa_d,
      xt_rsc_5_5_i_qa_d => peaseNTT_core_inst_xt_rsc_5_5_i_qa_d,
      xt_rsc_5_6_i_qa_d => peaseNTT_core_inst_xt_rsc_5_6_i_qa_d,
      xt_rsc_5_7_i_qa_d => peaseNTT_core_inst_xt_rsc_5_7_i_qa_d,
      xt_rsc_5_8_i_qa_d => peaseNTT_core_inst_xt_rsc_5_8_i_qa_d,
      xt_rsc_5_9_i_qa_d => peaseNTT_core_inst_xt_rsc_5_9_i_qa_d,
      xt_rsc_5_10_i_qa_d => peaseNTT_core_inst_xt_rsc_5_10_i_qa_d,
      xt_rsc_5_11_i_qa_d => peaseNTT_core_inst_xt_rsc_5_11_i_qa_d,
      xt_rsc_5_12_i_qa_d => peaseNTT_core_inst_xt_rsc_5_12_i_qa_d,
      xt_rsc_5_13_i_qa_d => peaseNTT_core_inst_xt_rsc_5_13_i_qa_d,
      xt_rsc_5_14_i_qa_d => peaseNTT_core_inst_xt_rsc_5_14_i_qa_d,
      xt_rsc_5_15_i_qa_d => peaseNTT_core_inst_xt_rsc_5_15_i_qa_d,
      xt_rsc_5_16_i_qa_d => peaseNTT_core_inst_xt_rsc_5_16_i_qa_d,
      xt_rsc_5_17_i_qa_d => peaseNTT_core_inst_xt_rsc_5_17_i_qa_d,
      xt_rsc_5_18_i_qa_d => peaseNTT_core_inst_xt_rsc_5_18_i_qa_d,
      xt_rsc_5_19_i_qa_d => peaseNTT_core_inst_xt_rsc_5_19_i_qa_d,
      xt_rsc_5_20_i_qa_d => peaseNTT_core_inst_xt_rsc_5_20_i_qa_d,
      xt_rsc_5_21_i_qa_d => peaseNTT_core_inst_xt_rsc_5_21_i_qa_d,
      xt_rsc_5_22_i_qa_d => peaseNTT_core_inst_xt_rsc_5_22_i_qa_d,
      xt_rsc_5_23_i_qa_d => peaseNTT_core_inst_xt_rsc_5_23_i_qa_d,
      xt_rsc_5_24_i_qa_d => peaseNTT_core_inst_xt_rsc_5_24_i_qa_d,
      xt_rsc_5_25_i_qa_d => peaseNTT_core_inst_xt_rsc_5_25_i_qa_d,
      xt_rsc_5_26_i_qa_d => peaseNTT_core_inst_xt_rsc_5_26_i_qa_d,
      xt_rsc_5_27_i_qa_d => peaseNTT_core_inst_xt_rsc_5_27_i_qa_d,
      xt_rsc_5_28_i_qa_d => peaseNTT_core_inst_xt_rsc_5_28_i_qa_d,
      xt_rsc_5_29_i_qa_d => peaseNTT_core_inst_xt_rsc_5_29_i_qa_d,
      xt_rsc_5_30_i_qa_d => peaseNTT_core_inst_xt_rsc_5_30_i_qa_d,
      xt_rsc_5_31_i_qa_d => peaseNTT_core_inst_xt_rsc_5_31_i_qa_d,
      xt_rsc_6_0_i_qa_d => peaseNTT_core_inst_xt_rsc_6_0_i_qa_d,
      xt_rsc_6_1_i_qa_d => peaseNTT_core_inst_xt_rsc_6_1_i_qa_d,
      xt_rsc_6_2_i_qa_d => peaseNTT_core_inst_xt_rsc_6_2_i_qa_d,
      xt_rsc_6_3_i_qa_d => peaseNTT_core_inst_xt_rsc_6_3_i_qa_d,
      xt_rsc_6_4_i_qa_d => peaseNTT_core_inst_xt_rsc_6_4_i_qa_d,
      xt_rsc_6_5_i_qa_d => peaseNTT_core_inst_xt_rsc_6_5_i_qa_d,
      xt_rsc_6_6_i_qa_d => peaseNTT_core_inst_xt_rsc_6_6_i_qa_d,
      xt_rsc_6_7_i_qa_d => peaseNTT_core_inst_xt_rsc_6_7_i_qa_d,
      xt_rsc_6_8_i_qa_d => peaseNTT_core_inst_xt_rsc_6_8_i_qa_d,
      xt_rsc_6_9_i_qa_d => peaseNTT_core_inst_xt_rsc_6_9_i_qa_d,
      xt_rsc_6_10_i_qa_d => peaseNTT_core_inst_xt_rsc_6_10_i_qa_d,
      xt_rsc_6_11_i_qa_d => peaseNTT_core_inst_xt_rsc_6_11_i_qa_d,
      xt_rsc_6_12_i_qa_d => peaseNTT_core_inst_xt_rsc_6_12_i_qa_d,
      xt_rsc_6_13_i_qa_d => peaseNTT_core_inst_xt_rsc_6_13_i_qa_d,
      xt_rsc_6_14_i_qa_d => peaseNTT_core_inst_xt_rsc_6_14_i_qa_d,
      xt_rsc_6_15_i_qa_d => peaseNTT_core_inst_xt_rsc_6_15_i_qa_d,
      xt_rsc_6_16_i_qa_d => peaseNTT_core_inst_xt_rsc_6_16_i_qa_d,
      xt_rsc_6_17_i_qa_d => peaseNTT_core_inst_xt_rsc_6_17_i_qa_d,
      xt_rsc_6_18_i_qa_d => peaseNTT_core_inst_xt_rsc_6_18_i_qa_d,
      xt_rsc_6_19_i_qa_d => peaseNTT_core_inst_xt_rsc_6_19_i_qa_d,
      xt_rsc_6_20_i_qa_d => peaseNTT_core_inst_xt_rsc_6_20_i_qa_d,
      xt_rsc_6_21_i_qa_d => peaseNTT_core_inst_xt_rsc_6_21_i_qa_d,
      xt_rsc_6_22_i_qa_d => peaseNTT_core_inst_xt_rsc_6_22_i_qa_d,
      xt_rsc_6_23_i_qa_d => peaseNTT_core_inst_xt_rsc_6_23_i_qa_d,
      xt_rsc_6_24_i_qa_d => peaseNTT_core_inst_xt_rsc_6_24_i_qa_d,
      xt_rsc_6_25_i_qa_d => peaseNTT_core_inst_xt_rsc_6_25_i_qa_d,
      xt_rsc_6_26_i_qa_d => peaseNTT_core_inst_xt_rsc_6_26_i_qa_d,
      xt_rsc_6_27_i_qa_d => peaseNTT_core_inst_xt_rsc_6_27_i_qa_d,
      xt_rsc_6_28_i_qa_d => peaseNTT_core_inst_xt_rsc_6_28_i_qa_d,
      xt_rsc_6_29_i_qa_d => peaseNTT_core_inst_xt_rsc_6_29_i_qa_d,
      xt_rsc_6_30_i_qa_d => peaseNTT_core_inst_xt_rsc_6_30_i_qa_d,
      xt_rsc_6_31_i_qa_d => peaseNTT_core_inst_xt_rsc_6_31_i_qa_d,
      xt_rsc_7_0_i_qa_d => peaseNTT_core_inst_xt_rsc_7_0_i_qa_d,
      xt_rsc_7_1_i_qa_d => peaseNTT_core_inst_xt_rsc_7_1_i_qa_d,
      xt_rsc_7_2_i_qa_d => peaseNTT_core_inst_xt_rsc_7_2_i_qa_d,
      xt_rsc_7_3_i_qa_d => peaseNTT_core_inst_xt_rsc_7_3_i_qa_d,
      xt_rsc_7_4_i_qa_d => peaseNTT_core_inst_xt_rsc_7_4_i_qa_d,
      xt_rsc_7_5_i_qa_d => peaseNTT_core_inst_xt_rsc_7_5_i_qa_d,
      xt_rsc_7_6_i_qa_d => peaseNTT_core_inst_xt_rsc_7_6_i_qa_d,
      xt_rsc_7_7_i_qa_d => peaseNTT_core_inst_xt_rsc_7_7_i_qa_d,
      xt_rsc_7_8_i_qa_d => peaseNTT_core_inst_xt_rsc_7_8_i_qa_d,
      xt_rsc_7_9_i_qa_d => peaseNTT_core_inst_xt_rsc_7_9_i_qa_d,
      xt_rsc_7_10_i_qa_d => peaseNTT_core_inst_xt_rsc_7_10_i_qa_d,
      xt_rsc_7_11_i_qa_d => peaseNTT_core_inst_xt_rsc_7_11_i_qa_d,
      xt_rsc_7_12_i_qa_d => peaseNTT_core_inst_xt_rsc_7_12_i_qa_d,
      xt_rsc_7_13_i_qa_d => peaseNTT_core_inst_xt_rsc_7_13_i_qa_d,
      xt_rsc_7_14_i_qa_d => peaseNTT_core_inst_xt_rsc_7_14_i_qa_d,
      xt_rsc_7_15_i_qa_d => peaseNTT_core_inst_xt_rsc_7_15_i_qa_d,
      xt_rsc_7_16_i_qa_d => peaseNTT_core_inst_xt_rsc_7_16_i_qa_d,
      xt_rsc_7_17_i_qa_d => peaseNTT_core_inst_xt_rsc_7_17_i_qa_d,
      xt_rsc_7_18_i_qa_d => peaseNTT_core_inst_xt_rsc_7_18_i_qa_d,
      xt_rsc_7_19_i_qa_d => peaseNTT_core_inst_xt_rsc_7_19_i_qa_d,
      xt_rsc_7_20_i_qa_d => peaseNTT_core_inst_xt_rsc_7_20_i_qa_d,
      xt_rsc_7_21_i_qa_d => peaseNTT_core_inst_xt_rsc_7_21_i_qa_d,
      xt_rsc_7_22_i_qa_d => peaseNTT_core_inst_xt_rsc_7_22_i_qa_d,
      xt_rsc_7_23_i_qa_d => peaseNTT_core_inst_xt_rsc_7_23_i_qa_d,
      xt_rsc_7_24_i_qa_d => peaseNTT_core_inst_xt_rsc_7_24_i_qa_d,
      xt_rsc_7_25_i_qa_d => peaseNTT_core_inst_xt_rsc_7_25_i_qa_d,
      xt_rsc_7_26_i_qa_d => peaseNTT_core_inst_xt_rsc_7_26_i_qa_d,
      xt_rsc_7_27_i_qa_d => peaseNTT_core_inst_xt_rsc_7_27_i_qa_d,
      xt_rsc_7_28_i_qa_d => peaseNTT_core_inst_xt_rsc_7_28_i_qa_d,
      xt_rsc_7_29_i_qa_d => peaseNTT_core_inst_xt_rsc_7_29_i_qa_d,
      xt_rsc_7_30_i_qa_d => peaseNTT_core_inst_xt_rsc_7_30_i_qa_d,
      xt_rsc_7_31_i_qa_d => peaseNTT_core_inst_xt_rsc_7_31_i_qa_d,
      twiddle_rsc_0_0_i_adra_d => peaseNTT_core_inst_twiddle_rsc_0_0_i_adra_d,
      twiddle_rsc_0_0_i_qa_d => peaseNTT_core_inst_twiddle_rsc_0_0_i_qa_d,
      twiddle_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_twiddle_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_1_i_adra_d => peaseNTT_core_inst_twiddle_rsc_0_1_i_adra_d,
      twiddle_rsc_0_1_i_qa_d => peaseNTT_core_inst_twiddle_rsc_0_1_i_qa_d,
      twiddle_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_twiddle_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_2_i_adra_d => peaseNTT_core_inst_twiddle_rsc_0_2_i_adra_d,
      twiddle_rsc_0_2_i_qa_d => peaseNTT_core_inst_twiddle_rsc_0_2_i_qa_d,
      twiddle_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_twiddle_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_3_i_adra_d => peaseNTT_core_inst_twiddle_rsc_0_3_i_adra_d,
      twiddle_rsc_0_3_i_qa_d => peaseNTT_core_inst_twiddle_rsc_0_3_i_qa_d,
      twiddle_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_twiddle_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_4_i_adra_d => peaseNTT_core_inst_twiddle_rsc_0_4_i_adra_d,
      twiddle_rsc_0_4_i_qa_d => peaseNTT_core_inst_twiddle_rsc_0_4_i_qa_d,
      twiddle_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_twiddle_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_5_i_adra_d => peaseNTT_core_inst_twiddle_rsc_0_5_i_adra_d,
      twiddle_rsc_0_5_i_qa_d => peaseNTT_core_inst_twiddle_rsc_0_5_i_qa_d,
      twiddle_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_twiddle_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_6_i_adra_d => peaseNTT_core_inst_twiddle_rsc_0_6_i_adra_d,
      twiddle_rsc_0_6_i_qa_d => peaseNTT_core_inst_twiddle_rsc_0_6_i_qa_d,
      twiddle_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_twiddle_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_7_i_adra_d => peaseNTT_core_inst_twiddle_rsc_0_7_i_adra_d,
      twiddle_rsc_0_7_i_qa_d => peaseNTT_core_inst_twiddle_rsc_0_7_i_qa_d,
      twiddle_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_twiddle_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_8_i_adra_d => peaseNTT_core_inst_twiddle_rsc_0_8_i_adra_d,
      twiddle_rsc_0_8_i_qa_d => peaseNTT_core_inst_twiddle_rsc_0_8_i_qa_d,
      twiddle_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_twiddle_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_9_i_adra_d => peaseNTT_core_inst_twiddle_rsc_0_9_i_adra_d,
      twiddle_rsc_0_9_i_qa_d => peaseNTT_core_inst_twiddle_rsc_0_9_i_qa_d,
      twiddle_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_twiddle_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_10_i_adra_d => peaseNTT_core_inst_twiddle_rsc_0_10_i_adra_d,
      twiddle_rsc_0_10_i_qa_d => peaseNTT_core_inst_twiddle_rsc_0_10_i_qa_d,
      twiddle_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_twiddle_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_11_i_adra_d => peaseNTT_core_inst_twiddle_rsc_0_11_i_adra_d,
      twiddle_rsc_0_11_i_qa_d => peaseNTT_core_inst_twiddle_rsc_0_11_i_qa_d,
      twiddle_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_twiddle_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_12_i_adra_d => peaseNTT_core_inst_twiddle_rsc_0_12_i_adra_d,
      twiddle_rsc_0_12_i_qa_d => peaseNTT_core_inst_twiddle_rsc_0_12_i_qa_d,
      twiddle_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_twiddle_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_13_i_adra_d => peaseNTT_core_inst_twiddle_rsc_0_13_i_adra_d,
      twiddle_rsc_0_13_i_qa_d => peaseNTT_core_inst_twiddle_rsc_0_13_i_qa_d,
      twiddle_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_twiddle_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_14_i_adra_d => peaseNTT_core_inst_twiddle_rsc_0_14_i_adra_d,
      twiddle_rsc_0_14_i_qa_d => peaseNTT_core_inst_twiddle_rsc_0_14_i_qa_d,
      twiddle_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_twiddle_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_15_i_adra_d => peaseNTT_core_inst_twiddle_rsc_0_15_i_adra_d,
      twiddle_rsc_0_15_i_qa_d => peaseNTT_core_inst_twiddle_rsc_0_15_i_qa_d,
      twiddle_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_twiddle_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_0_i_adra_d => peaseNTT_core_inst_twiddle_h_rsc_0_0_i_adra_d,
      twiddle_h_rsc_0_0_i_qa_d => peaseNTT_core_inst_twiddle_h_rsc_0_0_i_qa_d,
      twiddle_h_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_twiddle_h_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_1_i_adra_d => peaseNTT_core_inst_twiddle_h_rsc_0_1_i_adra_d,
      twiddle_h_rsc_0_1_i_qa_d => peaseNTT_core_inst_twiddle_h_rsc_0_1_i_qa_d,
      twiddle_h_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_twiddle_h_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_2_i_adra_d => peaseNTT_core_inst_twiddle_h_rsc_0_2_i_adra_d,
      twiddle_h_rsc_0_2_i_qa_d => peaseNTT_core_inst_twiddle_h_rsc_0_2_i_qa_d,
      twiddle_h_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_twiddle_h_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_3_i_adra_d => peaseNTT_core_inst_twiddle_h_rsc_0_3_i_adra_d,
      twiddle_h_rsc_0_3_i_qa_d => peaseNTT_core_inst_twiddle_h_rsc_0_3_i_qa_d,
      twiddle_h_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_twiddle_h_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_4_i_adra_d => peaseNTT_core_inst_twiddle_h_rsc_0_4_i_adra_d,
      twiddle_h_rsc_0_4_i_qa_d => peaseNTT_core_inst_twiddle_h_rsc_0_4_i_qa_d,
      twiddle_h_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_twiddle_h_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_5_i_adra_d => peaseNTT_core_inst_twiddle_h_rsc_0_5_i_adra_d,
      twiddle_h_rsc_0_5_i_qa_d => peaseNTT_core_inst_twiddle_h_rsc_0_5_i_qa_d,
      twiddle_h_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_twiddle_h_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_6_i_adra_d => peaseNTT_core_inst_twiddle_h_rsc_0_6_i_adra_d,
      twiddle_h_rsc_0_6_i_qa_d => peaseNTT_core_inst_twiddle_h_rsc_0_6_i_qa_d,
      twiddle_h_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_twiddle_h_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_7_i_adra_d => peaseNTT_core_inst_twiddle_h_rsc_0_7_i_adra_d,
      twiddle_h_rsc_0_7_i_qa_d => peaseNTT_core_inst_twiddle_h_rsc_0_7_i_qa_d,
      twiddle_h_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_twiddle_h_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_8_i_adra_d => peaseNTT_core_inst_twiddle_h_rsc_0_8_i_adra_d,
      twiddle_h_rsc_0_8_i_qa_d => peaseNTT_core_inst_twiddle_h_rsc_0_8_i_qa_d,
      twiddle_h_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_twiddle_h_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_9_i_adra_d => peaseNTT_core_inst_twiddle_h_rsc_0_9_i_adra_d,
      twiddle_h_rsc_0_9_i_qa_d => peaseNTT_core_inst_twiddle_h_rsc_0_9_i_qa_d,
      twiddle_h_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_twiddle_h_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_10_i_adra_d => peaseNTT_core_inst_twiddle_h_rsc_0_10_i_adra_d,
      twiddle_h_rsc_0_10_i_qa_d => peaseNTT_core_inst_twiddle_h_rsc_0_10_i_qa_d,
      twiddle_h_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_twiddle_h_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_11_i_adra_d => peaseNTT_core_inst_twiddle_h_rsc_0_11_i_adra_d,
      twiddle_h_rsc_0_11_i_qa_d => peaseNTT_core_inst_twiddle_h_rsc_0_11_i_qa_d,
      twiddle_h_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_twiddle_h_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_12_i_adra_d => peaseNTT_core_inst_twiddle_h_rsc_0_12_i_adra_d,
      twiddle_h_rsc_0_12_i_qa_d => peaseNTT_core_inst_twiddle_h_rsc_0_12_i_qa_d,
      twiddle_h_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_twiddle_h_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_13_i_adra_d => peaseNTT_core_inst_twiddle_h_rsc_0_13_i_adra_d,
      twiddle_h_rsc_0_13_i_qa_d => peaseNTT_core_inst_twiddle_h_rsc_0_13_i_qa_d,
      twiddle_h_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_twiddle_h_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_14_i_adra_d => peaseNTT_core_inst_twiddle_h_rsc_0_14_i_adra_d,
      twiddle_h_rsc_0_14_i_qa_d => peaseNTT_core_inst_twiddle_h_rsc_0_14_i_qa_d,
      twiddle_h_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_twiddle_h_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_15_i_adra_d => peaseNTT_core_inst_twiddle_h_rsc_0_15_i_adra_d,
      twiddle_h_rsc_0_15_i_qa_d => peaseNTT_core_inst_twiddle_h_rsc_0_15_i_qa_d,
      twiddle_h_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_twiddle_h_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yt_rsc_0_0_i_d_d_pff => peaseNTT_core_inst_yt_rsc_0_0_i_d_d_pff,
      yt_rsc_0_0_i_radr_d_pff => peaseNTT_core_inst_yt_rsc_0_0_i_radr_d_pff,
      yt_rsc_0_0_i_wadr_d_pff => peaseNTT_core_inst_yt_rsc_0_0_i_wadr_d_pff,
      yt_rsc_0_0_i_we_d_pff => yt_rsc_0_0_i_we_d_iff,
      yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_pff => yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff,
      yt_rsc_0_1_i_d_d_pff => peaseNTT_core_inst_yt_rsc_0_1_i_d_d_pff,
      yt_rsc_0_1_i_wadr_d_pff => peaseNTT_core_inst_yt_rsc_0_1_i_wadr_d_pff,
      yt_rsc_0_2_i_d_d_pff => peaseNTT_core_inst_yt_rsc_0_2_i_d_d_pff,
      yt_rsc_0_2_i_wadr_d_pff => peaseNTT_core_inst_yt_rsc_0_2_i_wadr_d_pff,
      yt_rsc_0_3_i_d_d_pff => peaseNTT_core_inst_yt_rsc_0_3_i_d_d_pff,
      yt_rsc_0_3_i_wadr_d_pff => peaseNTT_core_inst_yt_rsc_0_3_i_wadr_d_pff,
      yt_rsc_0_4_i_d_d_pff => peaseNTT_core_inst_yt_rsc_0_4_i_d_d_pff,
      yt_rsc_0_4_i_wadr_d_pff => peaseNTT_core_inst_yt_rsc_0_4_i_wadr_d_pff,
      yt_rsc_0_5_i_d_d_pff => peaseNTT_core_inst_yt_rsc_0_5_i_d_d_pff,
      yt_rsc_0_5_i_wadr_d_pff => peaseNTT_core_inst_yt_rsc_0_5_i_wadr_d_pff,
      yt_rsc_0_6_i_d_d_pff => peaseNTT_core_inst_yt_rsc_0_6_i_d_d_pff,
      yt_rsc_0_6_i_wadr_d_pff => peaseNTT_core_inst_yt_rsc_0_6_i_wadr_d_pff,
      yt_rsc_0_7_i_d_d_pff => peaseNTT_core_inst_yt_rsc_0_7_i_d_d_pff,
      yt_rsc_0_8_i_d_d_pff => peaseNTT_core_inst_yt_rsc_0_8_i_d_d_pff,
      yt_rsc_0_9_i_d_d_pff => peaseNTT_core_inst_yt_rsc_0_9_i_d_d_pff,
      yt_rsc_0_10_i_d_d_pff => peaseNTT_core_inst_yt_rsc_0_10_i_d_d_pff,
      yt_rsc_0_10_i_wadr_d_pff => peaseNTT_core_inst_yt_rsc_0_10_i_wadr_d_pff,
      yt_rsc_0_11_i_d_d_pff => peaseNTT_core_inst_yt_rsc_0_11_i_d_d_pff,
      yt_rsc_0_11_i_wadr_d_pff => peaseNTT_core_inst_yt_rsc_0_11_i_wadr_d_pff,
      yt_rsc_0_12_i_d_d_pff => peaseNTT_core_inst_yt_rsc_0_12_i_d_d_pff,
      yt_rsc_0_13_i_d_d_pff => peaseNTT_core_inst_yt_rsc_0_13_i_d_d_pff,
      yt_rsc_0_14_i_d_d_pff => peaseNTT_core_inst_yt_rsc_0_14_i_d_d_pff,
      yt_rsc_0_15_i_d_d_pff => peaseNTT_core_inst_yt_rsc_0_15_i_d_d_pff,
      yt_rsc_0_16_i_we_d_pff => yt_rsc_0_16_i_we_d_iff,
      yt_rsc_1_0_i_we_d_pff => yt_rsc_1_0_i_we_d_iff,
      yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_pff => yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff,
      yt_rsc_1_16_i_we_d_pff => yt_rsc_1_16_i_we_d_iff,
      yt_rsc_2_0_i_we_d_pff => yt_rsc_2_0_i_we_d_iff,
      yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_pff => yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff,
      yt_rsc_2_16_i_we_d_pff => yt_rsc_2_16_i_we_d_iff,
      yt_rsc_3_0_i_we_d_pff => yt_rsc_3_0_i_we_d_iff,
      yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_pff => yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff,
      yt_rsc_3_16_i_we_d_pff => yt_rsc_3_16_i_we_d_iff,
      yt_rsc_4_0_i_d_d_pff => peaseNTT_core_inst_yt_rsc_4_0_i_d_d_pff,
      yt_rsc_4_0_i_wadr_d_pff => peaseNTT_core_inst_yt_rsc_4_0_i_wadr_d_pff,
      yt_rsc_4_0_i_we_d_pff => yt_rsc_4_0_i_we_d_iff,
      yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_pff => yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff,
      yt_rsc_4_1_i_d_d_pff => peaseNTT_core_inst_yt_rsc_4_1_i_d_d_pff,
      yt_rsc_4_1_i_wadr_d_pff => peaseNTT_core_inst_yt_rsc_4_1_i_wadr_d_pff,
      yt_rsc_4_2_i_d_d_pff => peaseNTT_core_inst_yt_rsc_4_2_i_d_d_pff,
      yt_rsc_4_2_i_wadr_d_pff => peaseNTT_core_inst_yt_rsc_4_2_i_wadr_d_pff,
      yt_rsc_4_3_i_d_d_pff => peaseNTT_core_inst_yt_rsc_4_3_i_d_d_pff,
      yt_rsc_4_3_i_wadr_d_pff => peaseNTT_core_inst_yt_rsc_4_3_i_wadr_d_pff,
      yt_rsc_4_4_i_d_d_pff => peaseNTT_core_inst_yt_rsc_4_4_i_d_d_pff,
      yt_rsc_4_4_i_wadr_d_pff => peaseNTT_core_inst_yt_rsc_4_4_i_wadr_d_pff,
      yt_rsc_4_5_i_d_d_pff => peaseNTT_core_inst_yt_rsc_4_5_i_d_d_pff,
      yt_rsc_4_5_i_wadr_d_pff => peaseNTT_core_inst_yt_rsc_4_5_i_wadr_d_pff,
      yt_rsc_4_6_i_d_d_pff => peaseNTT_core_inst_yt_rsc_4_6_i_d_d_pff,
      yt_rsc_4_6_i_wadr_d_pff => peaseNTT_core_inst_yt_rsc_4_6_i_wadr_d_pff,
      yt_rsc_4_7_i_d_d_pff => peaseNTT_core_inst_yt_rsc_4_7_i_d_d_pff,
      yt_rsc_4_8_i_d_d_pff => peaseNTT_core_inst_yt_rsc_4_8_i_d_d_pff,
      yt_rsc_4_9_i_d_d_pff => peaseNTT_core_inst_yt_rsc_4_9_i_d_d_pff,
      yt_rsc_4_9_i_wadr_d_pff => peaseNTT_core_inst_yt_rsc_4_9_i_wadr_d_pff,
      yt_rsc_4_10_i_d_d_pff => peaseNTT_core_inst_yt_rsc_4_10_i_d_d_pff,
      yt_rsc_4_10_i_wadr_d_pff => peaseNTT_core_inst_yt_rsc_4_10_i_wadr_d_pff,
      yt_rsc_4_11_i_d_d_pff => peaseNTT_core_inst_yt_rsc_4_11_i_d_d_pff,
      yt_rsc_4_11_i_wadr_d_pff => peaseNTT_core_inst_yt_rsc_4_11_i_wadr_d_pff,
      yt_rsc_4_12_i_d_d_pff => peaseNTT_core_inst_yt_rsc_4_12_i_d_d_pff,
      yt_rsc_4_13_i_d_d_pff => peaseNTT_core_inst_yt_rsc_4_13_i_d_d_pff,
      yt_rsc_4_14_i_d_d_pff => peaseNTT_core_inst_yt_rsc_4_14_i_d_d_pff,
      yt_rsc_4_15_i_d_d_pff => peaseNTT_core_inst_yt_rsc_4_15_i_d_d_pff,
      yt_rsc_4_16_i_we_d_pff => yt_rsc_4_16_i_we_d_iff,
      yt_rsc_5_0_i_we_d_pff => yt_rsc_5_0_i_we_d_iff,
      yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_pff => yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff,
      yt_rsc_5_16_i_we_d_pff => yt_rsc_5_16_i_we_d_iff,
      yt_rsc_6_0_i_we_d_pff => yt_rsc_6_0_i_we_d_iff,
      yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_pff => yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff,
      yt_rsc_6_16_i_we_d_pff => yt_rsc_6_16_i_we_d_iff,
      yt_rsc_7_0_i_we_d_pff => yt_rsc_7_0_i_we_d_iff,
      yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_pff => yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff,
      yt_rsc_7_16_i_we_d_pff => yt_rsc_7_16_i_we_d_iff,
      xt_rsc_0_0_i_adra_d_pff => peaseNTT_core_inst_xt_rsc_0_0_i_adra_d_pff,
      xt_rsc_0_0_i_da_d_pff => peaseNTT_core_inst_xt_rsc_0_0_i_da_d_pff,
      xt_rsc_0_0_i_wea_d_pff => xt_rsc_0_0_i_wea_d_iff,
      xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff => xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      xt_rsc_0_1_i_adra_d_pff => peaseNTT_core_inst_xt_rsc_0_1_i_adra_d_pff,
      xt_rsc_0_1_i_da_d_pff => peaseNTT_core_inst_xt_rsc_0_1_i_da_d_pff,
      xt_rsc_0_2_i_adra_d_pff => peaseNTT_core_inst_xt_rsc_0_2_i_adra_d_pff,
      xt_rsc_0_2_i_da_d_pff => peaseNTT_core_inst_xt_rsc_0_2_i_da_d_pff,
      xt_rsc_0_3_i_adra_d_pff => peaseNTT_core_inst_xt_rsc_0_3_i_adra_d_pff,
      xt_rsc_0_3_i_da_d_pff => peaseNTT_core_inst_xt_rsc_0_3_i_da_d_pff,
      xt_rsc_0_4_i_adra_d_pff => peaseNTT_core_inst_xt_rsc_0_4_i_adra_d_pff,
      xt_rsc_0_4_i_da_d_pff => peaseNTT_core_inst_xt_rsc_0_4_i_da_d_pff,
      xt_rsc_0_5_i_adra_d_pff => peaseNTT_core_inst_xt_rsc_0_5_i_adra_d_pff,
      xt_rsc_0_5_i_da_d_pff => peaseNTT_core_inst_xt_rsc_0_5_i_da_d_pff,
      xt_rsc_0_6_i_adra_d_pff => peaseNTT_core_inst_xt_rsc_0_6_i_adra_d_pff,
      xt_rsc_0_6_i_da_d_pff => peaseNTT_core_inst_xt_rsc_0_6_i_da_d_pff,
      xt_rsc_0_7_i_adra_d_pff => peaseNTT_core_inst_xt_rsc_0_7_i_adra_d_pff,
      xt_rsc_0_7_i_da_d_pff => peaseNTT_core_inst_xt_rsc_0_7_i_da_d_pff,
      xt_rsc_0_8_i_adra_d_pff => peaseNTT_core_inst_xt_rsc_0_8_i_adra_d_pff,
      xt_rsc_0_8_i_da_d_pff => peaseNTT_core_inst_xt_rsc_0_8_i_da_d_pff,
      xt_rsc_0_9_i_adra_d_pff => peaseNTT_core_inst_xt_rsc_0_9_i_adra_d_pff,
      xt_rsc_0_9_i_da_d_pff => peaseNTT_core_inst_xt_rsc_0_9_i_da_d_pff,
      xt_rsc_0_10_i_adra_d_pff => peaseNTT_core_inst_xt_rsc_0_10_i_adra_d_pff,
      xt_rsc_0_10_i_da_d_pff => peaseNTT_core_inst_xt_rsc_0_10_i_da_d_pff,
      xt_rsc_0_11_i_adra_d_pff => peaseNTT_core_inst_xt_rsc_0_11_i_adra_d_pff,
      xt_rsc_0_11_i_da_d_pff => peaseNTT_core_inst_xt_rsc_0_11_i_da_d_pff,
      xt_rsc_0_12_i_adra_d_pff => peaseNTT_core_inst_xt_rsc_0_12_i_adra_d_pff,
      xt_rsc_0_12_i_da_d_pff => peaseNTT_core_inst_xt_rsc_0_12_i_da_d_pff,
      xt_rsc_0_13_i_adra_d_pff => peaseNTT_core_inst_xt_rsc_0_13_i_adra_d_pff,
      xt_rsc_0_13_i_da_d_pff => peaseNTT_core_inst_xt_rsc_0_13_i_da_d_pff,
      xt_rsc_0_14_i_adra_d_pff => peaseNTT_core_inst_xt_rsc_0_14_i_adra_d_pff,
      xt_rsc_0_14_i_da_d_pff => peaseNTT_core_inst_xt_rsc_0_14_i_da_d_pff,
      xt_rsc_0_15_i_adra_d_pff => peaseNTT_core_inst_xt_rsc_0_15_i_adra_d_pff,
      xt_rsc_0_15_i_da_d_pff => peaseNTT_core_inst_xt_rsc_0_15_i_da_d_pff,
      xt_rsc_0_16_i_wea_d_pff => xt_rsc_0_16_i_wea_d_iff,
      xt_rsc_1_0_i_wea_d_pff => xt_rsc_1_0_i_wea_d_iff,
      xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff => xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      xt_rsc_1_16_i_wea_d_pff => xt_rsc_1_16_i_wea_d_iff,
      xt_rsc_2_0_i_wea_d_pff => xt_rsc_2_0_i_wea_d_iff,
      xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff => xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      xt_rsc_2_16_i_wea_d_pff => xt_rsc_2_16_i_wea_d_iff,
      xt_rsc_3_0_i_wea_d_pff => xt_rsc_3_0_i_wea_d_iff,
      xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff => xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      xt_rsc_3_16_i_wea_d_pff => xt_rsc_3_16_i_wea_d_iff,
      xt_rsc_4_0_i_da_d_pff => peaseNTT_core_inst_xt_rsc_4_0_i_da_d_pff,
      xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff => xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      xt_rsc_4_1_i_adra_d_pff => peaseNTT_core_inst_xt_rsc_4_1_i_adra_d_pff,
      xt_rsc_4_1_i_da_d_pff => peaseNTT_core_inst_xt_rsc_4_1_i_da_d_pff,
      xt_rsc_4_2_i_adra_d_pff => peaseNTT_core_inst_xt_rsc_4_2_i_adra_d_pff,
      xt_rsc_4_2_i_da_d_pff => peaseNTT_core_inst_xt_rsc_4_2_i_da_d_pff,
      xt_rsc_4_3_i_da_d_pff => peaseNTT_core_inst_xt_rsc_4_3_i_da_d_pff,
      xt_rsc_4_4_i_da_d_pff => peaseNTT_core_inst_xt_rsc_4_4_i_da_d_pff,
      xt_rsc_4_5_i_da_d_pff => peaseNTT_core_inst_xt_rsc_4_5_i_da_d_pff,
      xt_rsc_4_6_i_da_d_pff => peaseNTT_core_inst_xt_rsc_4_6_i_da_d_pff,
      xt_rsc_4_7_i_da_d_pff => peaseNTT_core_inst_xt_rsc_4_7_i_da_d_pff,
      xt_rsc_4_8_i_da_d_pff => peaseNTT_core_inst_xt_rsc_4_8_i_da_d_pff,
      xt_rsc_4_9_i_adra_d_pff => peaseNTT_core_inst_xt_rsc_4_9_i_adra_d_pff,
      xt_rsc_4_9_i_da_d_pff => peaseNTT_core_inst_xt_rsc_4_9_i_da_d_pff,
      xt_rsc_4_10_i_adra_d_pff => peaseNTT_core_inst_xt_rsc_4_10_i_adra_d_pff,
      xt_rsc_4_10_i_da_d_pff => peaseNTT_core_inst_xt_rsc_4_10_i_da_d_pff,
      xt_rsc_4_11_i_da_d_pff => peaseNTT_core_inst_xt_rsc_4_11_i_da_d_pff,
      xt_rsc_4_12_i_da_d_pff => peaseNTT_core_inst_xt_rsc_4_12_i_da_d_pff,
      xt_rsc_4_13_i_da_d_pff => peaseNTT_core_inst_xt_rsc_4_13_i_da_d_pff,
      xt_rsc_4_14_i_da_d_pff => peaseNTT_core_inst_xt_rsc_4_14_i_da_d_pff,
      xt_rsc_4_15_i_da_d_pff => peaseNTT_core_inst_xt_rsc_4_15_i_da_d_pff,
      xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff => xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff => xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff => xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff
    );
  peaseNTT_core_inst_p_rsc_dat <= p_rsc_dat;
  peaseNTT_core_inst_yt_rsc_0_0_i_q_d <= yt_rsc_0_0_i_q_d;
  peaseNTT_core_inst_yt_rsc_0_1_i_q_d <= yt_rsc_0_1_i_q_d;
  peaseNTT_core_inst_yt_rsc_0_2_i_q_d <= yt_rsc_0_2_i_q_d;
  peaseNTT_core_inst_yt_rsc_0_3_i_q_d <= yt_rsc_0_3_i_q_d;
  peaseNTT_core_inst_yt_rsc_0_4_i_q_d <= yt_rsc_0_4_i_q_d;
  peaseNTT_core_inst_yt_rsc_0_5_i_q_d <= yt_rsc_0_5_i_q_d;
  peaseNTT_core_inst_yt_rsc_0_6_i_q_d <= yt_rsc_0_6_i_q_d;
  peaseNTT_core_inst_yt_rsc_0_7_i_q_d <= yt_rsc_0_7_i_q_d;
  peaseNTT_core_inst_yt_rsc_0_8_i_q_d <= yt_rsc_0_8_i_q_d;
  peaseNTT_core_inst_yt_rsc_0_9_i_q_d <= yt_rsc_0_9_i_q_d;
  peaseNTT_core_inst_yt_rsc_0_10_i_q_d <= yt_rsc_0_10_i_q_d;
  peaseNTT_core_inst_yt_rsc_0_11_i_q_d <= yt_rsc_0_11_i_q_d;
  peaseNTT_core_inst_yt_rsc_0_12_i_q_d <= yt_rsc_0_12_i_q_d;
  peaseNTT_core_inst_yt_rsc_0_13_i_q_d <= yt_rsc_0_13_i_q_d;
  peaseNTT_core_inst_yt_rsc_0_14_i_q_d <= yt_rsc_0_14_i_q_d;
  peaseNTT_core_inst_yt_rsc_0_15_i_q_d <= yt_rsc_0_15_i_q_d;
  peaseNTT_core_inst_yt_rsc_0_16_i_q_d <= yt_rsc_0_16_i_q_d;
  peaseNTT_core_inst_yt_rsc_0_17_i_q_d <= yt_rsc_0_17_i_q_d;
  peaseNTT_core_inst_yt_rsc_0_18_i_q_d <= yt_rsc_0_18_i_q_d;
  peaseNTT_core_inst_yt_rsc_0_19_i_q_d <= yt_rsc_0_19_i_q_d;
  peaseNTT_core_inst_yt_rsc_0_20_i_q_d <= yt_rsc_0_20_i_q_d;
  peaseNTT_core_inst_yt_rsc_0_21_i_q_d <= yt_rsc_0_21_i_q_d;
  peaseNTT_core_inst_yt_rsc_0_22_i_q_d <= yt_rsc_0_22_i_q_d;
  peaseNTT_core_inst_yt_rsc_0_23_i_q_d <= yt_rsc_0_23_i_q_d;
  peaseNTT_core_inst_yt_rsc_0_24_i_q_d <= yt_rsc_0_24_i_q_d;
  peaseNTT_core_inst_yt_rsc_0_25_i_q_d <= yt_rsc_0_25_i_q_d;
  peaseNTT_core_inst_yt_rsc_0_26_i_q_d <= yt_rsc_0_26_i_q_d;
  peaseNTT_core_inst_yt_rsc_0_27_i_q_d <= yt_rsc_0_27_i_q_d;
  peaseNTT_core_inst_yt_rsc_0_28_i_q_d <= yt_rsc_0_28_i_q_d;
  peaseNTT_core_inst_yt_rsc_0_29_i_q_d <= yt_rsc_0_29_i_q_d;
  peaseNTT_core_inst_yt_rsc_0_30_i_q_d <= yt_rsc_0_30_i_q_d;
  peaseNTT_core_inst_yt_rsc_0_31_i_q_d <= yt_rsc_0_31_i_q_d;
  peaseNTT_core_inst_yt_rsc_1_0_i_q_d <= yt_rsc_1_0_i_q_d;
  peaseNTT_core_inst_yt_rsc_1_1_i_q_d <= yt_rsc_1_1_i_q_d;
  peaseNTT_core_inst_yt_rsc_1_2_i_q_d <= yt_rsc_1_2_i_q_d;
  peaseNTT_core_inst_yt_rsc_1_3_i_q_d <= yt_rsc_1_3_i_q_d;
  peaseNTT_core_inst_yt_rsc_1_4_i_q_d <= yt_rsc_1_4_i_q_d;
  peaseNTT_core_inst_yt_rsc_1_5_i_q_d <= yt_rsc_1_5_i_q_d;
  peaseNTT_core_inst_yt_rsc_1_6_i_q_d <= yt_rsc_1_6_i_q_d;
  peaseNTT_core_inst_yt_rsc_1_7_i_q_d <= yt_rsc_1_7_i_q_d;
  peaseNTT_core_inst_yt_rsc_1_8_i_q_d <= yt_rsc_1_8_i_q_d;
  peaseNTT_core_inst_yt_rsc_1_9_i_q_d <= yt_rsc_1_9_i_q_d;
  peaseNTT_core_inst_yt_rsc_1_10_i_q_d <= yt_rsc_1_10_i_q_d;
  peaseNTT_core_inst_yt_rsc_1_11_i_q_d <= yt_rsc_1_11_i_q_d;
  peaseNTT_core_inst_yt_rsc_1_12_i_q_d <= yt_rsc_1_12_i_q_d;
  peaseNTT_core_inst_yt_rsc_1_13_i_q_d <= yt_rsc_1_13_i_q_d;
  peaseNTT_core_inst_yt_rsc_1_14_i_q_d <= yt_rsc_1_14_i_q_d;
  peaseNTT_core_inst_yt_rsc_1_15_i_q_d <= yt_rsc_1_15_i_q_d;
  peaseNTT_core_inst_yt_rsc_1_16_i_q_d <= yt_rsc_1_16_i_q_d;
  peaseNTT_core_inst_yt_rsc_1_17_i_q_d <= yt_rsc_1_17_i_q_d;
  peaseNTT_core_inst_yt_rsc_1_18_i_q_d <= yt_rsc_1_18_i_q_d;
  peaseNTT_core_inst_yt_rsc_1_19_i_q_d <= yt_rsc_1_19_i_q_d;
  peaseNTT_core_inst_yt_rsc_1_20_i_q_d <= yt_rsc_1_20_i_q_d;
  peaseNTT_core_inst_yt_rsc_1_21_i_q_d <= yt_rsc_1_21_i_q_d;
  peaseNTT_core_inst_yt_rsc_1_22_i_q_d <= yt_rsc_1_22_i_q_d;
  peaseNTT_core_inst_yt_rsc_1_23_i_q_d <= yt_rsc_1_23_i_q_d;
  peaseNTT_core_inst_yt_rsc_1_24_i_q_d <= yt_rsc_1_24_i_q_d;
  peaseNTT_core_inst_yt_rsc_1_25_i_q_d <= yt_rsc_1_25_i_q_d;
  peaseNTT_core_inst_yt_rsc_1_26_i_q_d <= yt_rsc_1_26_i_q_d;
  peaseNTT_core_inst_yt_rsc_1_27_i_q_d <= yt_rsc_1_27_i_q_d;
  peaseNTT_core_inst_yt_rsc_1_28_i_q_d <= yt_rsc_1_28_i_q_d;
  peaseNTT_core_inst_yt_rsc_1_29_i_q_d <= yt_rsc_1_29_i_q_d;
  peaseNTT_core_inst_yt_rsc_1_30_i_q_d <= yt_rsc_1_30_i_q_d;
  peaseNTT_core_inst_yt_rsc_1_31_i_q_d <= yt_rsc_1_31_i_q_d;
  peaseNTT_core_inst_yt_rsc_2_0_i_q_d <= yt_rsc_2_0_i_q_d;
  peaseNTT_core_inst_yt_rsc_2_1_i_q_d <= yt_rsc_2_1_i_q_d;
  peaseNTT_core_inst_yt_rsc_2_2_i_q_d <= yt_rsc_2_2_i_q_d;
  peaseNTT_core_inst_yt_rsc_2_3_i_q_d <= yt_rsc_2_3_i_q_d;
  peaseNTT_core_inst_yt_rsc_2_4_i_q_d <= yt_rsc_2_4_i_q_d;
  peaseNTT_core_inst_yt_rsc_2_5_i_q_d <= yt_rsc_2_5_i_q_d;
  peaseNTT_core_inst_yt_rsc_2_6_i_q_d <= yt_rsc_2_6_i_q_d;
  peaseNTT_core_inst_yt_rsc_2_7_i_q_d <= yt_rsc_2_7_i_q_d;
  peaseNTT_core_inst_yt_rsc_2_8_i_q_d <= yt_rsc_2_8_i_q_d;
  peaseNTT_core_inst_yt_rsc_2_9_i_q_d <= yt_rsc_2_9_i_q_d;
  peaseNTT_core_inst_yt_rsc_2_10_i_q_d <= yt_rsc_2_10_i_q_d;
  peaseNTT_core_inst_yt_rsc_2_11_i_q_d <= yt_rsc_2_11_i_q_d;
  peaseNTT_core_inst_yt_rsc_2_12_i_q_d <= yt_rsc_2_12_i_q_d;
  peaseNTT_core_inst_yt_rsc_2_13_i_q_d <= yt_rsc_2_13_i_q_d;
  peaseNTT_core_inst_yt_rsc_2_14_i_q_d <= yt_rsc_2_14_i_q_d;
  peaseNTT_core_inst_yt_rsc_2_15_i_q_d <= yt_rsc_2_15_i_q_d;
  peaseNTT_core_inst_yt_rsc_2_16_i_q_d <= yt_rsc_2_16_i_q_d;
  peaseNTT_core_inst_yt_rsc_2_17_i_q_d <= yt_rsc_2_17_i_q_d;
  peaseNTT_core_inst_yt_rsc_2_18_i_q_d <= yt_rsc_2_18_i_q_d;
  peaseNTT_core_inst_yt_rsc_2_19_i_q_d <= yt_rsc_2_19_i_q_d;
  peaseNTT_core_inst_yt_rsc_2_20_i_q_d <= yt_rsc_2_20_i_q_d;
  peaseNTT_core_inst_yt_rsc_2_21_i_q_d <= yt_rsc_2_21_i_q_d;
  peaseNTT_core_inst_yt_rsc_2_22_i_q_d <= yt_rsc_2_22_i_q_d;
  peaseNTT_core_inst_yt_rsc_2_23_i_q_d <= yt_rsc_2_23_i_q_d;
  peaseNTT_core_inst_yt_rsc_2_24_i_q_d <= yt_rsc_2_24_i_q_d;
  peaseNTT_core_inst_yt_rsc_2_25_i_q_d <= yt_rsc_2_25_i_q_d;
  peaseNTT_core_inst_yt_rsc_2_26_i_q_d <= yt_rsc_2_26_i_q_d;
  peaseNTT_core_inst_yt_rsc_2_27_i_q_d <= yt_rsc_2_27_i_q_d;
  peaseNTT_core_inst_yt_rsc_2_28_i_q_d <= yt_rsc_2_28_i_q_d;
  peaseNTT_core_inst_yt_rsc_2_29_i_q_d <= yt_rsc_2_29_i_q_d;
  peaseNTT_core_inst_yt_rsc_2_30_i_q_d <= yt_rsc_2_30_i_q_d;
  peaseNTT_core_inst_yt_rsc_2_31_i_q_d <= yt_rsc_2_31_i_q_d;
  peaseNTT_core_inst_yt_rsc_3_0_i_q_d <= yt_rsc_3_0_i_q_d;
  peaseNTT_core_inst_yt_rsc_3_1_i_q_d <= yt_rsc_3_1_i_q_d;
  peaseNTT_core_inst_yt_rsc_3_2_i_q_d <= yt_rsc_3_2_i_q_d;
  peaseNTT_core_inst_yt_rsc_3_3_i_q_d <= yt_rsc_3_3_i_q_d;
  peaseNTT_core_inst_yt_rsc_3_4_i_q_d <= yt_rsc_3_4_i_q_d;
  peaseNTT_core_inst_yt_rsc_3_5_i_q_d <= yt_rsc_3_5_i_q_d;
  peaseNTT_core_inst_yt_rsc_3_6_i_q_d <= yt_rsc_3_6_i_q_d;
  peaseNTT_core_inst_yt_rsc_3_7_i_q_d <= yt_rsc_3_7_i_q_d;
  peaseNTT_core_inst_yt_rsc_3_8_i_q_d <= yt_rsc_3_8_i_q_d;
  peaseNTT_core_inst_yt_rsc_3_9_i_q_d <= yt_rsc_3_9_i_q_d;
  peaseNTT_core_inst_yt_rsc_3_10_i_q_d <= yt_rsc_3_10_i_q_d;
  peaseNTT_core_inst_yt_rsc_3_11_i_q_d <= yt_rsc_3_11_i_q_d;
  peaseNTT_core_inst_yt_rsc_3_12_i_q_d <= yt_rsc_3_12_i_q_d;
  peaseNTT_core_inst_yt_rsc_3_13_i_q_d <= yt_rsc_3_13_i_q_d;
  peaseNTT_core_inst_yt_rsc_3_14_i_q_d <= yt_rsc_3_14_i_q_d;
  peaseNTT_core_inst_yt_rsc_3_15_i_q_d <= yt_rsc_3_15_i_q_d;
  peaseNTT_core_inst_yt_rsc_3_16_i_q_d <= yt_rsc_3_16_i_q_d;
  peaseNTT_core_inst_yt_rsc_3_17_i_q_d <= yt_rsc_3_17_i_q_d;
  peaseNTT_core_inst_yt_rsc_3_18_i_q_d <= yt_rsc_3_18_i_q_d;
  peaseNTT_core_inst_yt_rsc_3_19_i_q_d <= yt_rsc_3_19_i_q_d;
  peaseNTT_core_inst_yt_rsc_3_20_i_q_d <= yt_rsc_3_20_i_q_d;
  peaseNTT_core_inst_yt_rsc_3_21_i_q_d <= yt_rsc_3_21_i_q_d;
  peaseNTT_core_inst_yt_rsc_3_22_i_q_d <= yt_rsc_3_22_i_q_d;
  peaseNTT_core_inst_yt_rsc_3_23_i_q_d <= yt_rsc_3_23_i_q_d;
  peaseNTT_core_inst_yt_rsc_3_24_i_q_d <= yt_rsc_3_24_i_q_d;
  peaseNTT_core_inst_yt_rsc_3_25_i_q_d <= yt_rsc_3_25_i_q_d;
  peaseNTT_core_inst_yt_rsc_3_26_i_q_d <= yt_rsc_3_26_i_q_d;
  peaseNTT_core_inst_yt_rsc_3_27_i_q_d <= yt_rsc_3_27_i_q_d;
  peaseNTT_core_inst_yt_rsc_3_28_i_q_d <= yt_rsc_3_28_i_q_d;
  peaseNTT_core_inst_yt_rsc_3_29_i_q_d <= yt_rsc_3_29_i_q_d;
  peaseNTT_core_inst_yt_rsc_3_30_i_q_d <= yt_rsc_3_30_i_q_d;
  peaseNTT_core_inst_yt_rsc_3_31_i_q_d <= yt_rsc_3_31_i_q_d;
  peaseNTT_core_inst_yt_rsc_4_0_i_q_d <= yt_rsc_4_0_i_q_d;
  peaseNTT_core_inst_yt_rsc_4_1_i_q_d <= yt_rsc_4_1_i_q_d;
  peaseNTT_core_inst_yt_rsc_4_2_i_q_d <= yt_rsc_4_2_i_q_d;
  peaseNTT_core_inst_yt_rsc_4_3_i_q_d <= yt_rsc_4_3_i_q_d;
  peaseNTT_core_inst_yt_rsc_4_4_i_q_d <= yt_rsc_4_4_i_q_d;
  peaseNTT_core_inst_yt_rsc_4_5_i_q_d <= yt_rsc_4_5_i_q_d;
  peaseNTT_core_inst_yt_rsc_4_6_i_q_d <= yt_rsc_4_6_i_q_d;
  peaseNTT_core_inst_yt_rsc_4_7_i_q_d <= yt_rsc_4_7_i_q_d;
  peaseNTT_core_inst_yt_rsc_4_8_i_q_d <= yt_rsc_4_8_i_q_d;
  peaseNTT_core_inst_yt_rsc_4_9_i_q_d <= yt_rsc_4_9_i_q_d;
  peaseNTT_core_inst_yt_rsc_4_10_i_q_d <= yt_rsc_4_10_i_q_d;
  peaseNTT_core_inst_yt_rsc_4_11_i_q_d <= yt_rsc_4_11_i_q_d;
  peaseNTT_core_inst_yt_rsc_4_12_i_q_d <= yt_rsc_4_12_i_q_d;
  peaseNTT_core_inst_yt_rsc_4_13_i_q_d <= yt_rsc_4_13_i_q_d;
  peaseNTT_core_inst_yt_rsc_4_14_i_q_d <= yt_rsc_4_14_i_q_d;
  peaseNTT_core_inst_yt_rsc_4_15_i_q_d <= yt_rsc_4_15_i_q_d;
  peaseNTT_core_inst_yt_rsc_4_16_i_q_d <= yt_rsc_4_16_i_q_d;
  peaseNTT_core_inst_yt_rsc_4_17_i_q_d <= yt_rsc_4_17_i_q_d;
  peaseNTT_core_inst_yt_rsc_4_18_i_q_d <= yt_rsc_4_18_i_q_d;
  peaseNTT_core_inst_yt_rsc_4_19_i_q_d <= yt_rsc_4_19_i_q_d;
  peaseNTT_core_inst_yt_rsc_4_20_i_q_d <= yt_rsc_4_20_i_q_d;
  peaseNTT_core_inst_yt_rsc_4_21_i_q_d <= yt_rsc_4_21_i_q_d;
  peaseNTT_core_inst_yt_rsc_4_22_i_q_d <= yt_rsc_4_22_i_q_d;
  peaseNTT_core_inst_yt_rsc_4_23_i_q_d <= yt_rsc_4_23_i_q_d;
  peaseNTT_core_inst_yt_rsc_4_24_i_q_d <= yt_rsc_4_24_i_q_d;
  peaseNTT_core_inst_yt_rsc_4_25_i_q_d <= yt_rsc_4_25_i_q_d;
  peaseNTT_core_inst_yt_rsc_4_26_i_q_d <= yt_rsc_4_26_i_q_d;
  peaseNTT_core_inst_yt_rsc_4_27_i_q_d <= yt_rsc_4_27_i_q_d;
  peaseNTT_core_inst_yt_rsc_4_28_i_q_d <= yt_rsc_4_28_i_q_d;
  peaseNTT_core_inst_yt_rsc_4_29_i_q_d <= yt_rsc_4_29_i_q_d;
  peaseNTT_core_inst_yt_rsc_4_30_i_q_d <= yt_rsc_4_30_i_q_d;
  peaseNTT_core_inst_yt_rsc_4_31_i_q_d <= yt_rsc_4_31_i_q_d;
  peaseNTT_core_inst_yt_rsc_5_0_i_q_d <= yt_rsc_5_0_i_q_d;
  peaseNTT_core_inst_yt_rsc_5_1_i_q_d <= yt_rsc_5_1_i_q_d;
  peaseNTT_core_inst_yt_rsc_5_2_i_q_d <= yt_rsc_5_2_i_q_d;
  peaseNTT_core_inst_yt_rsc_5_3_i_q_d <= yt_rsc_5_3_i_q_d;
  peaseNTT_core_inst_yt_rsc_5_4_i_q_d <= yt_rsc_5_4_i_q_d;
  peaseNTT_core_inst_yt_rsc_5_5_i_q_d <= yt_rsc_5_5_i_q_d;
  peaseNTT_core_inst_yt_rsc_5_6_i_q_d <= yt_rsc_5_6_i_q_d;
  peaseNTT_core_inst_yt_rsc_5_7_i_q_d <= yt_rsc_5_7_i_q_d;
  peaseNTT_core_inst_yt_rsc_5_8_i_q_d <= yt_rsc_5_8_i_q_d;
  peaseNTT_core_inst_yt_rsc_5_9_i_q_d <= yt_rsc_5_9_i_q_d;
  peaseNTT_core_inst_yt_rsc_5_10_i_q_d <= yt_rsc_5_10_i_q_d;
  peaseNTT_core_inst_yt_rsc_5_11_i_q_d <= yt_rsc_5_11_i_q_d;
  peaseNTT_core_inst_yt_rsc_5_12_i_q_d <= yt_rsc_5_12_i_q_d;
  peaseNTT_core_inst_yt_rsc_5_13_i_q_d <= yt_rsc_5_13_i_q_d;
  peaseNTT_core_inst_yt_rsc_5_14_i_q_d <= yt_rsc_5_14_i_q_d;
  peaseNTT_core_inst_yt_rsc_5_15_i_q_d <= yt_rsc_5_15_i_q_d;
  peaseNTT_core_inst_yt_rsc_5_16_i_q_d <= yt_rsc_5_16_i_q_d;
  peaseNTT_core_inst_yt_rsc_5_17_i_q_d <= yt_rsc_5_17_i_q_d;
  peaseNTT_core_inst_yt_rsc_5_18_i_q_d <= yt_rsc_5_18_i_q_d;
  peaseNTT_core_inst_yt_rsc_5_19_i_q_d <= yt_rsc_5_19_i_q_d;
  peaseNTT_core_inst_yt_rsc_5_20_i_q_d <= yt_rsc_5_20_i_q_d;
  peaseNTT_core_inst_yt_rsc_5_21_i_q_d <= yt_rsc_5_21_i_q_d;
  peaseNTT_core_inst_yt_rsc_5_22_i_q_d <= yt_rsc_5_22_i_q_d;
  peaseNTT_core_inst_yt_rsc_5_23_i_q_d <= yt_rsc_5_23_i_q_d;
  peaseNTT_core_inst_yt_rsc_5_24_i_q_d <= yt_rsc_5_24_i_q_d;
  peaseNTT_core_inst_yt_rsc_5_25_i_q_d <= yt_rsc_5_25_i_q_d;
  peaseNTT_core_inst_yt_rsc_5_26_i_q_d <= yt_rsc_5_26_i_q_d;
  peaseNTT_core_inst_yt_rsc_5_27_i_q_d <= yt_rsc_5_27_i_q_d;
  peaseNTT_core_inst_yt_rsc_5_28_i_q_d <= yt_rsc_5_28_i_q_d;
  peaseNTT_core_inst_yt_rsc_5_29_i_q_d <= yt_rsc_5_29_i_q_d;
  peaseNTT_core_inst_yt_rsc_5_30_i_q_d <= yt_rsc_5_30_i_q_d;
  peaseNTT_core_inst_yt_rsc_5_31_i_q_d <= yt_rsc_5_31_i_q_d;
  peaseNTT_core_inst_yt_rsc_6_0_i_q_d <= yt_rsc_6_0_i_q_d;
  peaseNTT_core_inst_yt_rsc_6_1_i_q_d <= yt_rsc_6_1_i_q_d;
  peaseNTT_core_inst_yt_rsc_6_2_i_q_d <= yt_rsc_6_2_i_q_d;
  peaseNTT_core_inst_yt_rsc_6_3_i_q_d <= yt_rsc_6_3_i_q_d;
  peaseNTT_core_inst_yt_rsc_6_4_i_q_d <= yt_rsc_6_4_i_q_d;
  peaseNTT_core_inst_yt_rsc_6_5_i_q_d <= yt_rsc_6_5_i_q_d;
  peaseNTT_core_inst_yt_rsc_6_6_i_q_d <= yt_rsc_6_6_i_q_d;
  peaseNTT_core_inst_yt_rsc_6_7_i_q_d <= yt_rsc_6_7_i_q_d;
  peaseNTT_core_inst_yt_rsc_6_8_i_q_d <= yt_rsc_6_8_i_q_d;
  peaseNTT_core_inst_yt_rsc_6_9_i_q_d <= yt_rsc_6_9_i_q_d;
  peaseNTT_core_inst_yt_rsc_6_10_i_q_d <= yt_rsc_6_10_i_q_d;
  peaseNTT_core_inst_yt_rsc_6_11_i_q_d <= yt_rsc_6_11_i_q_d;
  peaseNTT_core_inst_yt_rsc_6_12_i_q_d <= yt_rsc_6_12_i_q_d;
  peaseNTT_core_inst_yt_rsc_6_13_i_q_d <= yt_rsc_6_13_i_q_d;
  peaseNTT_core_inst_yt_rsc_6_14_i_q_d <= yt_rsc_6_14_i_q_d;
  peaseNTT_core_inst_yt_rsc_6_15_i_q_d <= yt_rsc_6_15_i_q_d;
  peaseNTT_core_inst_yt_rsc_6_16_i_q_d <= yt_rsc_6_16_i_q_d;
  peaseNTT_core_inst_yt_rsc_6_17_i_q_d <= yt_rsc_6_17_i_q_d;
  peaseNTT_core_inst_yt_rsc_6_18_i_q_d <= yt_rsc_6_18_i_q_d;
  peaseNTT_core_inst_yt_rsc_6_19_i_q_d <= yt_rsc_6_19_i_q_d;
  peaseNTT_core_inst_yt_rsc_6_20_i_q_d <= yt_rsc_6_20_i_q_d;
  peaseNTT_core_inst_yt_rsc_6_21_i_q_d <= yt_rsc_6_21_i_q_d;
  peaseNTT_core_inst_yt_rsc_6_22_i_q_d <= yt_rsc_6_22_i_q_d;
  peaseNTT_core_inst_yt_rsc_6_23_i_q_d <= yt_rsc_6_23_i_q_d;
  peaseNTT_core_inst_yt_rsc_6_24_i_q_d <= yt_rsc_6_24_i_q_d;
  peaseNTT_core_inst_yt_rsc_6_25_i_q_d <= yt_rsc_6_25_i_q_d;
  peaseNTT_core_inst_yt_rsc_6_26_i_q_d <= yt_rsc_6_26_i_q_d;
  peaseNTT_core_inst_yt_rsc_6_27_i_q_d <= yt_rsc_6_27_i_q_d;
  peaseNTT_core_inst_yt_rsc_6_28_i_q_d <= yt_rsc_6_28_i_q_d;
  peaseNTT_core_inst_yt_rsc_6_29_i_q_d <= yt_rsc_6_29_i_q_d;
  peaseNTT_core_inst_yt_rsc_6_30_i_q_d <= yt_rsc_6_30_i_q_d;
  peaseNTT_core_inst_yt_rsc_6_31_i_q_d <= yt_rsc_6_31_i_q_d;
  peaseNTT_core_inst_yt_rsc_7_0_i_q_d <= yt_rsc_7_0_i_q_d;
  peaseNTT_core_inst_yt_rsc_7_1_i_q_d <= yt_rsc_7_1_i_q_d;
  peaseNTT_core_inst_yt_rsc_7_2_i_q_d <= yt_rsc_7_2_i_q_d;
  peaseNTT_core_inst_yt_rsc_7_3_i_q_d <= yt_rsc_7_3_i_q_d;
  peaseNTT_core_inst_yt_rsc_7_4_i_q_d <= yt_rsc_7_4_i_q_d;
  peaseNTT_core_inst_yt_rsc_7_5_i_q_d <= yt_rsc_7_5_i_q_d;
  peaseNTT_core_inst_yt_rsc_7_6_i_q_d <= yt_rsc_7_6_i_q_d;
  peaseNTT_core_inst_yt_rsc_7_7_i_q_d <= yt_rsc_7_7_i_q_d;
  peaseNTT_core_inst_yt_rsc_7_8_i_q_d <= yt_rsc_7_8_i_q_d;
  peaseNTT_core_inst_yt_rsc_7_9_i_q_d <= yt_rsc_7_9_i_q_d;
  peaseNTT_core_inst_yt_rsc_7_10_i_q_d <= yt_rsc_7_10_i_q_d;
  peaseNTT_core_inst_yt_rsc_7_11_i_q_d <= yt_rsc_7_11_i_q_d;
  peaseNTT_core_inst_yt_rsc_7_12_i_q_d <= yt_rsc_7_12_i_q_d;
  peaseNTT_core_inst_yt_rsc_7_13_i_q_d <= yt_rsc_7_13_i_q_d;
  peaseNTT_core_inst_yt_rsc_7_14_i_q_d <= yt_rsc_7_14_i_q_d;
  peaseNTT_core_inst_yt_rsc_7_15_i_q_d <= yt_rsc_7_15_i_q_d;
  peaseNTT_core_inst_yt_rsc_7_16_i_q_d <= yt_rsc_7_16_i_q_d;
  peaseNTT_core_inst_yt_rsc_7_17_i_q_d <= yt_rsc_7_17_i_q_d;
  peaseNTT_core_inst_yt_rsc_7_18_i_q_d <= yt_rsc_7_18_i_q_d;
  peaseNTT_core_inst_yt_rsc_7_19_i_q_d <= yt_rsc_7_19_i_q_d;
  peaseNTT_core_inst_yt_rsc_7_20_i_q_d <= yt_rsc_7_20_i_q_d;
  peaseNTT_core_inst_yt_rsc_7_21_i_q_d <= yt_rsc_7_21_i_q_d;
  peaseNTT_core_inst_yt_rsc_7_22_i_q_d <= yt_rsc_7_22_i_q_d;
  peaseNTT_core_inst_yt_rsc_7_23_i_q_d <= yt_rsc_7_23_i_q_d;
  peaseNTT_core_inst_yt_rsc_7_24_i_q_d <= yt_rsc_7_24_i_q_d;
  peaseNTT_core_inst_yt_rsc_7_25_i_q_d <= yt_rsc_7_25_i_q_d;
  peaseNTT_core_inst_yt_rsc_7_26_i_q_d <= yt_rsc_7_26_i_q_d;
  peaseNTT_core_inst_yt_rsc_7_27_i_q_d <= yt_rsc_7_27_i_q_d;
  peaseNTT_core_inst_yt_rsc_7_28_i_q_d <= yt_rsc_7_28_i_q_d;
  peaseNTT_core_inst_yt_rsc_7_29_i_q_d <= yt_rsc_7_29_i_q_d;
  peaseNTT_core_inst_yt_rsc_7_30_i_q_d <= yt_rsc_7_30_i_q_d;
  peaseNTT_core_inst_yt_rsc_7_31_i_q_d <= yt_rsc_7_31_i_q_d;
  peaseNTT_core_inst_xt_rsc_0_0_i_qa_d <= xt_rsc_0_0_i_qa_d;
  peaseNTT_core_inst_xt_rsc_0_1_i_qa_d <= xt_rsc_0_1_i_qa_d;
  peaseNTT_core_inst_xt_rsc_0_2_i_qa_d <= xt_rsc_0_2_i_qa_d;
  peaseNTT_core_inst_xt_rsc_0_3_i_qa_d <= xt_rsc_0_3_i_qa_d;
  peaseNTT_core_inst_xt_rsc_0_4_i_qa_d <= xt_rsc_0_4_i_qa_d;
  peaseNTT_core_inst_xt_rsc_0_5_i_qa_d <= xt_rsc_0_5_i_qa_d;
  peaseNTT_core_inst_xt_rsc_0_6_i_qa_d <= xt_rsc_0_6_i_qa_d;
  peaseNTT_core_inst_xt_rsc_0_7_i_qa_d <= xt_rsc_0_7_i_qa_d;
  peaseNTT_core_inst_xt_rsc_0_8_i_qa_d <= xt_rsc_0_8_i_qa_d;
  peaseNTT_core_inst_xt_rsc_0_9_i_qa_d <= xt_rsc_0_9_i_qa_d;
  peaseNTT_core_inst_xt_rsc_0_10_i_qa_d <= xt_rsc_0_10_i_qa_d;
  peaseNTT_core_inst_xt_rsc_0_11_i_qa_d <= xt_rsc_0_11_i_qa_d;
  peaseNTT_core_inst_xt_rsc_0_12_i_qa_d <= xt_rsc_0_12_i_qa_d;
  peaseNTT_core_inst_xt_rsc_0_13_i_qa_d <= xt_rsc_0_13_i_qa_d;
  peaseNTT_core_inst_xt_rsc_0_14_i_qa_d <= xt_rsc_0_14_i_qa_d;
  peaseNTT_core_inst_xt_rsc_0_15_i_qa_d <= xt_rsc_0_15_i_qa_d;
  peaseNTT_core_inst_xt_rsc_0_16_i_qa_d <= xt_rsc_0_16_i_qa_d;
  peaseNTT_core_inst_xt_rsc_0_17_i_qa_d <= xt_rsc_0_17_i_qa_d;
  peaseNTT_core_inst_xt_rsc_0_18_i_qa_d <= xt_rsc_0_18_i_qa_d;
  peaseNTT_core_inst_xt_rsc_0_19_i_qa_d <= xt_rsc_0_19_i_qa_d;
  peaseNTT_core_inst_xt_rsc_0_20_i_qa_d <= xt_rsc_0_20_i_qa_d;
  peaseNTT_core_inst_xt_rsc_0_21_i_qa_d <= xt_rsc_0_21_i_qa_d;
  peaseNTT_core_inst_xt_rsc_0_22_i_qa_d <= xt_rsc_0_22_i_qa_d;
  peaseNTT_core_inst_xt_rsc_0_23_i_qa_d <= xt_rsc_0_23_i_qa_d;
  peaseNTT_core_inst_xt_rsc_0_24_i_qa_d <= xt_rsc_0_24_i_qa_d;
  peaseNTT_core_inst_xt_rsc_0_25_i_qa_d <= xt_rsc_0_25_i_qa_d;
  peaseNTT_core_inst_xt_rsc_0_26_i_qa_d <= xt_rsc_0_26_i_qa_d;
  peaseNTT_core_inst_xt_rsc_0_27_i_qa_d <= xt_rsc_0_27_i_qa_d;
  peaseNTT_core_inst_xt_rsc_0_28_i_qa_d <= xt_rsc_0_28_i_qa_d;
  peaseNTT_core_inst_xt_rsc_0_29_i_qa_d <= xt_rsc_0_29_i_qa_d;
  peaseNTT_core_inst_xt_rsc_0_30_i_qa_d <= xt_rsc_0_30_i_qa_d;
  peaseNTT_core_inst_xt_rsc_0_31_i_qa_d <= xt_rsc_0_31_i_qa_d;
  peaseNTT_core_inst_xt_rsc_1_0_i_qa_d <= xt_rsc_1_0_i_qa_d;
  peaseNTT_core_inst_xt_rsc_1_1_i_qa_d <= xt_rsc_1_1_i_qa_d;
  peaseNTT_core_inst_xt_rsc_1_2_i_qa_d <= xt_rsc_1_2_i_qa_d;
  peaseNTT_core_inst_xt_rsc_1_3_i_qa_d <= xt_rsc_1_3_i_qa_d;
  peaseNTT_core_inst_xt_rsc_1_4_i_qa_d <= xt_rsc_1_4_i_qa_d;
  peaseNTT_core_inst_xt_rsc_1_5_i_qa_d <= xt_rsc_1_5_i_qa_d;
  peaseNTT_core_inst_xt_rsc_1_6_i_qa_d <= xt_rsc_1_6_i_qa_d;
  peaseNTT_core_inst_xt_rsc_1_7_i_qa_d <= xt_rsc_1_7_i_qa_d;
  peaseNTT_core_inst_xt_rsc_1_8_i_qa_d <= xt_rsc_1_8_i_qa_d;
  peaseNTT_core_inst_xt_rsc_1_9_i_qa_d <= xt_rsc_1_9_i_qa_d;
  peaseNTT_core_inst_xt_rsc_1_10_i_qa_d <= xt_rsc_1_10_i_qa_d;
  peaseNTT_core_inst_xt_rsc_1_11_i_qa_d <= xt_rsc_1_11_i_qa_d;
  peaseNTT_core_inst_xt_rsc_1_12_i_qa_d <= xt_rsc_1_12_i_qa_d;
  peaseNTT_core_inst_xt_rsc_1_13_i_qa_d <= xt_rsc_1_13_i_qa_d;
  peaseNTT_core_inst_xt_rsc_1_14_i_qa_d <= xt_rsc_1_14_i_qa_d;
  peaseNTT_core_inst_xt_rsc_1_15_i_qa_d <= xt_rsc_1_15_i_qa_d;
  peaseNTT_core_inst_xt_rsc_1_16_i_qa_d <= xt_rsc_1_16_i_qa_d;
  peaseNTT_core_inst_xt_rsc_1_17_i_qa_d <= xt_rsc_1_17_i_qa_d;
  peaseNTT_core_inst_xt_rsc_1_18_i_qa_d <= xt_rsc_1_18_i_qa_d;
  peaseNTT_core_inst_xt_rsc_1_19_i_qa_d <= xt_rsc_1_19_i_qa_d;
  peaseNTT_core_inst_xt_rsc_1_20_i_qa_d <= xt_rsc_1_20_i_qa_d;
  peaseNTT_core_inst_xt_rsc_1_21_i_qa_d <= xt_rsc_1_21_i_qa_d;
  peaseNTT_core_inst_xt_rsc_1_22_i_qa_d <= xt_rsc_1_22_i_qa_d;
  peaseNTT_core_inst_xt_rsc_1_23_i_qa_d <= xt_rsc_1_23_i_qa_d;
  peaseNTT_core_inst_xt_rsc_1_24_i_qa_d <= xt_rsc_1_24_i_qa_d;
  peaseNTT_core_inst_xt_rsc_1_25_i_qa_d <= xt_rsc_1_25_i_qa_d;
  peaseNTT_core_inst_xt_rsc_1_26_i_qa_d <= xt_rsc_1_26_i_qa_d;
  peaseNTT_core_inst_xt_rsc_1_27_i_qa_d <= xt_rsc_1_27_i_qa_d;
  peaseNTT_core_inst_xt_rsc_1_28_i_qa_d <= xt_rsc_1_28_i_qa_d;
  peaseNTT_core_inst_xt_rsc_1_29_i_qa_d <= xt_rsc_1_29_i_qa_d;
  peaseNTT_core_inst_xt_rsc_1_30_i_qa_d <= xt_rsc_1_30_i_qa_d;
  peaseNTT_core_inst_xt_rsc_1_31_i_qa_d <= xt_rsc_1_31_i_qa_d;
  peaseNTT_core_inst_xt_rsc_2_0_i_qa_d <= xt_rsc_2_0_i_qa_d;
  peaseNTT_core_inst_xt_rsc_2_1_i_qa_d <= xt_rsc_2_1_i_qa_d;
  peaseNTT_core_inst_xt_rsc_2_2_i_qa_d <= xt_rsc_2_2_i_qa_d;
  peaseNTT_core_inst_xt_rsc_2_3_i_qa_d <= xt_rsc_2_3_i_qa_d;
  peaseNTT_core_inst_xt_rsc_2_4_i_qa_d <= xt_rsc_2_4_i_qa_d;
  peaseNTT_core_inst_xt_rsc_2_5_i_qa_d <= xt_rsc_2_5_i_qa_d;
  peaseNTT_core_inst_xt_rsc_2_6_i_qa_d <= xt_rsc_2_6_i_qa_d;
  peaseNTT_core_inst_xt_rsc_2_7_i_qa_d <= xt_rsc_2_7_i_qa_d;
  peaseNTT_core_inst_xt_rsc_2_8_i_qa_d <= xt_rsc_2_8_i_qa_d;
  peaseNTT_core_inst_xt_rsc_2_9_i_qa_d <= xt_rsc_2_9_i_qa_d;
  peaseNTT_core_inst_xt_rsc_2_10_i_qa_d <= xt_rsc_2_10_i_qa_d;
  peaseNTT_core_inst_xt_rsc_2_11_i_qa_d <= xt_rsc_2_11_i_qa_d;
  peaseNTT_core_inst_xt_rsc_2_12_i_qa_d <= xt_rsc_2_12_i_qa_d;
  peaseNTT_core_inst_xt_rsc_2_13_i_qa_d <= xt_rsc_2_13_i_qa_d;
  peaseNTT_core_inst_xt_rsc_2_14_i_qa_d <= xt_rsc_2_14_i_qa_d;
  peaseNTT_core_inst_xt_rsc_2_15_i_qa_d <= xt_rsc_2_15_i_qa_d;
  peaseNTT_core_inst_xt_rsc_2_16_i_qa_d <= xt_rsc_2_16_i_qa_d;
  peaseNTT_core_inst_xt_rsc_2_17_i_qa_d <= xt_rsc_2_17_i_qa_d;
  peaseNTT_core_inst_xt_rsc_2_18_i_qa_d <= xt_rsc_2_18_i_qa_d;
  peaseNTT_core_inst_xt_rsc_2_19_i_qa_d <= xt_rsc_2_19_i_qa_d;
  peaseNTT_core_inst_xt_rsc_2_20_i_qa_d <= xt_rsc_2_20_i_qa_d;
  peaseNTT_core_inst_xt_rsc_2_21_i_qa_d <= xt_rsc_2_21_i_qa_d;
  peaseNTT_core_inst_xt_rsc_2_22_i_qa_d <= xt_rsc_2_22_i_qa_d;
  peaseNTT_core_inst_xt_rsc_2_23_i_qa_d <= xt_rsc_2_23_i_qa_d;
  peaseNTT_core_inst_xt_rsc_2_24_i_qa_d <= xt_rsc_2_24_i_qa_d;
  peaseNTT_core_inst_xt_rsc_2_25_i_qa_d <= xt_rsc_2_25_i_qa_d;
  peaseNTT_core_inst_xt_rsc_2_26_i_qa_d <= xt_rsc_2_26_i_qa_d;
  peaseNTT_core_inst_xt_rsc_2_27_i_qa_d <= xt_rsc_2_27_i_qa_d;
  peaseNTT_core_inst_xt_rsc_2_28_i_qa_d <= xt_rsc_2_28_i_qa_d;
  peaseNTT_core_inst_xt_rsc_2_29_i_qa_d <= xt_rsc_2_29_i_qa_d;
  peaseNTT_core_inst_xt_rsc_2_30_i_qa_d <= xt_rsc_2_30_i_qa_d;
  peaseNTT_core_inst_xt_rsc_2_31_i_qa_d <= xt_rsc_2_31_i_qa_d;
  peaseNTT_core_inst_xt_rsc_3_0_i_qa_d <= xt_rsc_3_0_i_qa_d;
  peaseNTT_core_inst_xt_rsc_3_1_i_qa_d <= xt_rsc_3_1_i_qa_d;
  peaseNTT_core_inst_xt_rsc_3_2_i_qa_d <= xt_rsc_3_2_i_qa_d;
  peaseNTT_core_inst_xt_rsc_3_3_i_qa_d <= xt_rsc_3_3_i_qa_d;
  peaseNTT_core_inst_xt_rsc_3_4_i_qa_d <= xt_rsc_3_4_i_qa_d;
  peaseNTT_core_inst_xt_rsc_3_5_i_qa_d <= xt_rsc_3_5_i_qa_d;
  peaseNTT_core_inst_xt_rsc_3_6_i_qa_d <= xt_rsc_3_6_i_qa_d;
  peaseNTT_core_inst_xt_rsc_3_7_i_qa_d <= xt_rsc_3_7_i_qa_d;
  peaseNTT_core_inst_xt_rsc_3_8_i_qa_d <= xt_rsc_3_8_i_qa_d;
  peaseNTT_core_inst_xt_rsc_3_9_i_qa_d <= xt_rsc_3_9_i_qa_d;
  peaseNTT_core_inst_xt_rsc_3_10_i_qa_d <= xt_rsc_3_10_i_qa_d;
  peaseNTT_core_inst_xt_rsc_3_11_i_qa_d <= xt_rsc_3_11_i_qa_d;
  peaseNTT_core_inst_xt_rsc_3_12_i_qa_d <= xt_rsc_3_12_i_qa_d;
  peaseNTT_core_inst_xt_rsc_3_13_i_qa_d <= xt_rsc_3_13_i_qa_d;
  peaseNTT_core_inst_xt_rsc_3_14_i_qa_d <= xt_rsc_3_14_i_qa_d;
  peaseNTT_core_inst_xt_rsc_3_15_i_qa_d <= xt_rsc_3_15_i_qa_d;
  peaseNTT_core_inst_xt_rsc_3_16_i_qa_d <= xt_rsc_3_16_i_qa_d;
  peaseNTT_core_inst_xt_rsc_3_17_i_qa_d <= xt_rsc_3_17_i_qa_d;
  peaseNTT_core_inst_xt_rsc_3_18_i_qa_d <= xt_rsc_3_18_i_qa_d;
  peaseNTT_core_inst_xt_rsc_3_19_i_qa_d <= xt_rsc_3_19_i_qa_d;
  peaseNTT_core_inst_xt_rsc_3_20_i_qa_d <= xt_rsc_3_20_i_qa_d;
  peaseNTT_core_inst_xt_rsc_3_21_i_qa_d <= xt_rsc_3_21_i_qa_d;
  peaseNTT_core_inst_xt_rsc_3_22_i_qa_d <= xt_rsc_3_22_i_qa_d;
  peaseNTT_core_inst_xt_rsc_3_23_i_qa_d <= xt_rsc_3_23_i_qa_d;
  peaseNTT_core_inst_xt_rsc_3_24_i_qa_d <= xt_rsc_3_24_i_qa_d;
  peaseNTT_core_inst_xt_rsc_3_25_i_qa_d <= xt_rsc_3_25_i_qa_d;
  peaseNTT_core_inst_xt_rsc_3_26_i_qa_d <= xt_rsc_3_26_i_qa_d;
  peaseNTT_core_inst_xt_rsc_3_27_i_qa_d <= xt_rsc_3_27_i_qa_d;
  peaseNTT_core_inst_xt_rsc_3_28_i_qa_d <= xt_rsc_3_28_i_qa_d;
  peaseNTT_core_inst_xt_rsc_3_29_i_qa_d <= xt_rsc_3_29_i_qa_d;
  peaseNTT_core_inst_xt_rsc_3_30_i_qa_d <= xt_rsc_3_30_i_qa_d;
  peaseNTT_core_inst_xt_rsc_3_31_i_qa_d <= xt_rsc_3_31_i_qa_d;
  peaseNTT_core_inst_xt_rsc_4_0_i_qa_d <= xt_rsc_4_0_i_qa_d;
  peaseNTT_core_inst_xt_rsc_4_1_i_qa_d <= xt_rsc_4_1_i_qa_d;
  peaseNTT_core_inst_xt_rsc_4_2_i_qa_d <= xt_rsc_4_2_i_qa_d;
  peaseNTT_core_inst_xt_rsc_4_3_i_qa_d <= xt_rsc_4_3_i_qa_d;
  peaseNTT_core_inst_xt_rsc_4_4_i_qa_d <= xt_rsc_4_4_i_qa_d;
  peaseNTT_core_inst_xt_rsc_4_5_i_qa_d <= xt_rsc_4_5_i_qa_d;
  peaseNTT_core_inst_xt_rsc_4_6_i_qa_d <= xt_rsc_4_6_i_qa_d;
  peaseNTT_core_inst_xt_rsc_4_7_i_qa_d <= xt_rsc_4_7_i_qa_d;
  peaseNTT_core_inst_xt_rsc_4_8_i_qa_d <= xt_rsc_4_8_i_qa_d;
  peaseNTT_core_inst_xt_rsc_4_9_i_qa_d <= xt_rsc_4_9_i_qa_d;
  peaseNTT_core_inst_xt_rsc_4_10_i_qa_d <= xt_rsc_4_10_i_qa_d;
  peaseNTT_core_inst_xt_rsc_4_11_i_qa_d <= xt_rsc_4_11_i_qa_d;
  peaseNTT_core_inst_xt_rsc_4_12_i_qa_d <= xt_rsc_4_12_i_qa_d;
  peaseNTT_core_inst_xt_rsc_4_13_i_qa_d <= xt_rsc_4_13_i_qa_d;
  peaseNTT_core_inst_xt_rsc_4_14_i_qa_d <= xt_rsc_4_14_i_qa_d;
  peaseNTT_core_inst_xt_rsc_4_15_i_qa_d <= xt_rsc_4_15_i_qa_d;
  peaseNTT_core_inst_xt_rsc_4_16_i_qa_d <= xt_rsc_4_16_i_qa_d;
  peaseNTT_core_inst_xt_rsc_4_17_i_qa_d <= xt_rsc_4_17_i_qa_d;
  peaseNTT_core_inst_xt_rsc_4_18_i_qa_d <= xt_rsc_4_18_i_qa_d;
  peaseNTT_core_inst_xt_rsc_4_19_i_qa_d <= xt_rsc_4_19_i_qa_d;
  peaseNTT_core_inst_xt_rsc_4_20_i_qa_d <= xt_rsc_4_20_i_qa_d;
  peaseNTT_core_inst_xt_rsc_4_21_i_qa_d <= xt_rsc_4_21_i_qa_d;
  peaseNTT_core_inst_xt_rsc_4_22_i_qa_d <= xt_rsc_4_22_i_qa_d;
  peaseNTT_core_inst_xt_rsc_4_23_i_qa_d <= xt_rsc_4_23_i_qa_d;
  peaseNTT_core_inst_xt_rsc_4_24_i_qa_d <= xt_rsc_4_24_i_qa_d;
  peaseNTT_core_inst_xt_rsc_4_25_i_qa_d <= xt_rsc_4_25_i_qa_d;
  peaseNTT_core_inst_xt_rsc_4_26_i_qa_d <= xt_rsc_4_26_i_qa_d;
  peaseNTT_core_inst_xt_rsc_4_27_i_qa_d <= xt_rsc_4_27_i_qa_d;
  peaseNTT_core_inst_xt_rsc_4_28_i_qa_d <= xt_rsc_4_28_i_qa_d;
  peaseNTT_core_inst_xt_rsc_4_29_i_qa_d <= xt_rsc_4_29_i_qa_d;
  peaseNTT_core_inst_xt_rsc_4_30_i_qa_d <= xt_rsc_4_30_i_qa_d;
  peaseNTT_core_inst_xt_rsc_4_31_i_qa_d <= xt_rsc_4_31_i_qa_d;
  peaseNTT_core_inst_xt_rsc_5_0_i_qa_d <= xt_rsc_5_0_i_qa_d;
  peaseNTT_core_inst_xt_rsc_5_1_i_qa_d <= xt_rsc_5_1_i_qa_d;
  peaseNTT_core_inst_xt_rsc_5_2_i_qa_d <= xt_rsc_5_2_i_qa_d;
  peaseNTT_core_inst_xt_rsc_5_3_i_qa_d <= xt_rsc_5_3_i_qa_d;
  peaseNTT_core_inst_xt_rsc_5_4_i_qa_d <= xt_rsc_5_4_i_qa_d;
  peaseNTT_core_inst_xt_rsc_5_5_i_qa_d <= xt_rsc_5_5_i_qa_d;
  peaseNTT_core_inst_xt_rsc_5_6_i_qa_d <= xt_rsc_5_6_i_qa_d;
  peaseNTT_core_inst_xt_rsc_5_7_i_qa_d <= xt_rsc_5_7_i_qa_d;
  peaseNTT_core_inst_xt_rsc_5_8_i_qa_d <= xt_rsc_5_8_i_qa_d;
  peaseNTT_core_inst_xt_rsc_5_9_i_qa_d <= xt_rsc_5_9_i_qa_d;
  peaseNTT_core_inst_xt_rsc_5_10_i_qa_d <= xt_rsc_5_10_i_qa_d;
  peaseNTT_core_inst_xt_rsc_5_11_i_qa_d <= xt_rsc_5_11_i_qa_d;
  peaseNTT_core_inst_xt_rsc_5_12_i_qa_d <= xt_rsc_5_12_i_qa_d;
  peaseNTT_core_inst_xt_rsc_5_13_i_qa_d <= xt_rsc_5_13_i_qa_d;
  peaseNTT_core_inst_xt_rsc_5_14_i_qa_d <= xt_rsc_5_14_i_qa_d;
  peaseNTT_core_inst_xt_rsc_5_15_i_qa_d <= xt_rsc_5_15_i_qa_d;
  peaseNTT_core_inst_xt_rsc_5_16_i_qa_d <= xt_rsc_5_16_i_qa_d;
  peaseNTT_core_inst_xt_rsc_5_17_i_qa_d <= xt_rsc_5_17_i_qa_d;
  peaseNTT_core_inst_xt_rsc_5_18_i_qa_d <= xt_rsc_5_18_i_qa_d;
  peaseNTT_core_inst_xt_rsc_5_19_i_qa_d <= xt_rsc_5_19_i_qa_d;
  peaseNTT_core_inst_xt_rsc_5_20_i_qa_d <= xt_rsc_5_20_i_qa_d;
  peaseNTT_core_inst_xt_rsc_5_21_i_qa_d <= xt_rsc_5_21_i_qa_d;
  peaseNTT_core_inst_xt_rsc_5_22_i_qa_d <= xt_rsc_5_22_i_qa_d;
  peaseNTT_core_inst_xt_rsc_5_23_i_qa_d <= xt_rsc_5_23_i_qa_d;
  peaseNTT_core_inst_xt_rsc_5_24_i_qa_d <= xt_rsc_5_24_i_qa_d;
  peaseNTT_core_inst_xt_rsc_5_25_i_qa_d <= xt_rsc_5_25_i_qa_d;
  peaseNTT_core_inst_xt_rsc_5_26_i_qa_d <= xt_rsc_5_26_i_qa_d;
  peaseNTT_core_inst_xt_rsc_5_27_i_qa_d <= xt_rsc_5_27_i_qa_d;
  peaseNTT_core_inst_xt_rsc_5_28_i_qa_d <= xt_rsc_5_28_i_qa_d;
  peaseNTT_core_inst_xt_rsc_5_29_i_qa_d <= xt_rsc_5_29_i_qa_d;
  peaseNTT_core_inst_xt_rsc_5_30_i_qa_d <= xt_rsc_5_30_i_qa_d;
  peaseNTT_core_inst_xt_rsc_5_31_i_qa_d <= xt_rsc_5_31_i_qa_d;
  peaseNTT_core_inst_xt_rsc_6_0_i_qa_d <= xt_rsc_6_0_i_qa_d;
  peaseNTT_core_inst_xt_rsc_6_1_i_qa_d <= xt_rsc_6_1_i_qa_d;
  peaseNTT_core_inst_xt_rsc_6_2_i_qa_d <= xt_rsc_6_2_i_qa_d;
  peaseNTT_core_inst_xt_rsc_6_3_i_qa_d <= xt_rsc_6_3_i_qa_d;
  peaseNTT_core_inst_xt_rsc_6_4_i_qa_d <= xt_rsc_6_4_i_qa_d;
  peaseNTT_core_inst_xt_rsc_6_5_i_qa_d <= xt_rsc_6_5_i_qa_d;
  peaseNTT_core_inst_xt_rsc_6_6_i_qa_d <= xt_rsc_6_6_i_qa_d;
  peaseNTT_core_inst_xt_rsc_6_7_i_qa_d <= xt_rsc_6_7_i_qa_d;
  peaseNTT_core_inst_xt_rsc_6_8_i_qa_d <= xt_rsc_6_8_i_qa_d;
  peaseNTT_core_inst_xt_rsc_6_9_i_qa_d <= xt_rsc_6_9_i_qa_d;
  peaseNTT_core_inst_xt_rsc_6_10_i_qa_d <= xt_rsc_6_10_i_qa_d;
  peaseNTT_core_inst_xt_rsc_6_11_i_qa_d <= xt_rsc_6_11_i_qa_d;
  peaseNTT_core_inst_xt_rsc_6_12_i_qa_d <= xt_rsc_6_12_i_qa_d;
  peaseNTT_core_inst_xt_rsc_6_13_i_qa_d <= xt_rsc_6_13_i_qa_d;
  peaseNTT_core_inst_xt_rsc_6_14_i_qa_d <= xt_rsc_6_14_i_qa_d;
  peaseNTT_core_inst_xt_rsc_6_15_i_qa_d <= xt_rsc_6_15_i_qa_d;
  peaseNTT_core_inst_xt_rsc_6_16_i_qa_d <= xt_rsc_6_16_i_qa_d;
  peaseNTT_core_inst_xt_rsc_6_17_i_qa_d <= xt_rsc_6_17_i_qa_d;
  peaseNTT_core_inst_xt_rsc_6_18_i_qa_d <= xt_rsc_6_18_i_qa_d;
  peaseNTT_core_inst_xt_rsc_6_19_i_qa_d <= xt_rsc_6_19_i_qa_d;
  peaseNTT_core_inst_xt_rsc_6_20_i_qa_d <= xt_rsc_6_20_i_qa_d;
  peaseNTT_core_inst_xt_rsc_6_21_i_qa_d <= xt_rsc_6_21_i_qa_d;
  peaseNTT_core_inst_xt_rsc_6_22_i_qa_d <= xt_rsc_6_22_i_qa_d;
  peaseNTT_core_inst_xt_rsc_6_23_i_qa_d <= xt_rsc_6_23_i_qa_d;
  peaseNTT_core_inst_xt_rsc_6_24_i_qa_d <= xt_rsc_6_24_i_qa_d;
  peaseNTT_core_inst_xt_rsc_6_25_i_qa_d <= xt_rsc_6_25_i_qa_d;
  peaseNTT_core_inst_xt_rsc_6_26_i_qa_d <= xt_rsc_6_26_i_qa_d;
  peaseNTT_core_inst_xt_rsc_6_27_i_qa_d <= xt_rsc_6_27_i_qa_d;
  peaseNTT_core_inst_xt_rsc_6_28_i_qa_d <= xt_rsc_6_28_i_qa_d;
  peaseNTT_core_inst_xt_rsc_6_29_i_qa_d <= xt_rsc_6_29_i_qa_d;
  peaseNTT_core_inst_xt_rsc_6_30_i_qa_d <= xt_rsc_6_30_i_qa_d;
  peaseNTT_core_inst_xt_rsc_6_31_i_qa_d <= xt_rsc_6_31_i_qa_d;
  peaseNTT_core_inst_xt_rsc_7_0_i_qa_d <= xt_rsc_7_0_i_qa_d;
  peaseNTT_core_inst_xt_rsc_7_1_i_qa_d <= xt_rsc_7_1_i_qa_d;
  peaseNTT_core_inst_xt_rsc_7_2_i_qa_d <= xt_rsc_7_2_i_qa_d;
  peaseNTT_core_inst_xt_rsc_7_3_i_qa_d <= xt_rsc_7_3_i_qa_d;
  peaseNTT_core_inst_xt_rsc_7_4_i_qa_d <= xt_rsc_7_4_i_qa_d;
  peaseNTT_core_inst_xt_rsc_7_5_i_qa_d <= xt_rsc_7_5_i_qa_d;
  peaseNTT_core_inst_xt_rsc_7_6_i_qa_d <= xt_rsc_7_6_i_qa_d;
  peaseNTT_core_inst_xt_rsc_7_7_i_qa_d <= xt_rsc_7_7_i_qa_d;
  peaseNTT_core_inst_xt_rsc_7_8_i_qa_d <= xt_rsc_7_8_i_qa_d;
  peaseNTT_core_inst_xt_rsc_7_9_i_qa_d <= xt_rsc_7_9_i_qa_d;
  peaseNTT_core_inst_xt_rsc_7_10_i_qa_d <= xt_rsc_7_10_i_qa_d;
  peaseNTT_core_inst_xt_rsc_7_11_i_qa_d <= xt_rsc_7_11_i_qa_d;
  peaseNTT_core_inst_xt_rsc_7_12_i_qa_d <= xt_rsc_7_12_i_qa_d;
  peaseNTT_core_inst_xt_rsc_7_13_i_qa_d <= xt_rsc_7_13_i_qa_d;
  peaseNTT_core_inst_xt_rsc_7_14_i_qa_d <= xt_rsc_7_14_i_qa_d;
  peaseNTT_core_inst_xt_rsc_7_15_i_qa_d <= xt_rsc_7_15_i_qa_d;
  peaseNTT_core_inst_xt_rsc_7_16_i_qa_d <= xt_rsc_7_16_i_qa_d;
  peaseNTT_core_inst_xt_rsc_7_17_i_qa_d <= xt_rsc_7_17_i_qa_d;
  peaseNTT_core_inst_xt_rsc_7_18_i_qa_d <= xt_rsc_7_18_i_qa_d;
  peaseNTT_core_inst_xt_rsc_7_19_i_qa_d <= xt_rsc_7_19_i_qa_d;
  peaseNTT_core_inst_xt_rsc_7_20_i_qa_d <= xt_rsc_7_20_i_qa_d;
  peaseNTT_core_inst_xt_rsc_7_21_i_qa_d <= xt_rsc_7_21_i_qa_d;
  peaseNTT_core_inst_xt_rsc_7_22_i_qa_d <= xt_rsc_7_22_i_qa_d;
  peaseNTT_core_inst_xt_rsc_7_23_i_qa_d <= xt_rsc_7_23_i_qa_d;
  peaseNTT_core_inst_xt_rsc_7_24_i_qa_d <= xt_rsc_7_24_i_qa_d;
  peaseNTT_core_inst_xt_rsc_7_25_i_qa_d <= xt_rsc_7_25_i_qa_d;
  peaseNTT_core_inst_xt_rsc_7_26_i_qa_d <= xt_rsc_7_26_i_qa_d;
  peaseNTT_core_inst_xt_rsc_7_27_i_qa_d <= xt_rsc_7_27_i_qa_d;
  peaseNTT_core_inst_xt_rsc_7_28_i_qa_d <= xt_rsc_7_28_i_qa_d;
  peaseNTT_core_inst_xt_rsc_7_29_i_qa_d <= xt_rsc_7_29_i_qa_d;
  peaseNTT_core_inst_xt_rsc_7_30_i_qa_d <= xt_rsc_7_30_i_qa_d;
  peaseNTT_core_inst_xt_rsc_7_31_i_qa_d <= xt_rsc_7_31_i_qa_d;
  twiddle_rsc_0_0_i_adra_d <= peaseNTT_core_inst_twiddle_rsc_0_0_i_adra_d;
  peaseNTT_core_inst_twiddle_rsc_0_0_i_qa_d <= twiddle_rsc_0_0_i_qa_d;
  twiddle_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_twiddle_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_rsc_0_1_i_adra_d <= peaseNTT_core_inst_twiddle_rsc_0_1_i_adra_d;
  peaseNTT_core_inst_twiddle_rsc_0_1_i_qa_d <= twiddle_rsc_0_1_i_qa_d;
  twiddle_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_twiddle_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_rsc_0_2_i_adra_d <= peaseNTT_core_inst_twiddle_rsc_0_2_i_adra_d;
  peaseNTT_core_inst_twiddle_rsc_0_2_i_qa_d <= twiddle_rsc_0_2_i_qa_d;
  twiddle_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_twiddle_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_rsc_0_3_i_adra_d <= peaseNTT_core_inst_twiddle_rsc_0_3_i_adra_d;
  peaseNTT_core_inst_twiddle_rsc_0_3_i_qa_d <= twiddle_rsc_0_3_i_qa_d;
  twiddle_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_twiddle_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_rsc_0_4_i_adra_d <= peaseNTT_core_inst_twiddle_rsc_0_4_i_adra_d;
  peaseNTT_core_inst_twiddle_rsc_0_4_i_qa_d <= twiddle_rsc_0_4_i_qa_d;
  twiddle_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_twiddle_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_rsc_0_5_i_adra_d <= peaseNTT_core_inst_twiddle_rsc_0_5_i_adra_d;
  peaseNTT_core_inst_twiddle_rsc_0_5_i_qa_d <= twiddle_rsc_0_5_i_qa_d;
  twiddle_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_twiddle_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_rsc_0_6_i_adra_d <= peaseNTT_core_inst_twiddle_rsc_0_6_i_adra_d;
  peaseNTT_core_inst_twiddle_rsc_0_6_i_qa_d <= twiddle_rsc_0_6_i_qa_d;
  twiddle_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_twiddle_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_rsc_0_7_i_adra_d <= peaseNTT_core_inst_twiddle_rsc_0_7_i_adra_d;
  peaseNTT_core_inst_twiddle_rsc_0_7_i_qa_d <= twiddle_rsc_0_7_i_qa_d;
  twiddle_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_twiddle_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_rsc_0_8_i_adra_d <= peaseNTT_core_inst_twiddle_rsc_0_8_i_adra_d;
  peaseNTT_core_inst_twiddle_rsc_0_8_i_qa_d <= twiddle_rsc_0_8_i_qa_d;
  twiddle_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_twiddle_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_rsc_0_9_i_adra_d <= peaseNTT_core_inst_twiddle_rsc_0_9_i_adra_d;
  peaseNTT_core_inst_twiddle_rsc_0_9_i_qa_d <= twiddle_rsc_0_9_i_qa_d;
  twiddle_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_twiddle_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_rsc_0_10_i_adra_d <= peaseNTT_core_inst_twiddle_rsc_0_10_i_adra_d;
  peaseNTT_core_inst_twiddle_rsc_0_10_i_qa_d <= twiddle_rsc_0_10_i_qa_d;
  twiddle_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_twiddle_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_rsc_0_11_i_adra_d <= peaseNTT_core_inst_twiddle_rsc_0_11_i_adra_d;
  peaseNTT_core_inst_twiddle_rsc_0_11_i_qa_d <= twiddle_rsc_0_11_i_qa_d;
  twiddle_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_twiddle_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_rsc_0_12_i_adra_d <= peaseNTT_core_inst_twiddle_rsc_0_12_i_adra_d;
  peaseNTT_core_inst_twiddle_rsc_0_12_i_qa_d <= twiddle_rsc_0_12_i_qa_d;
  twiddle_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_twiddle_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_rsc_0_13_i_adra_d <= peaseNTT_core_inst_twiddle_rsc_0_13_i_adra_d;
  peaseNTT_core_inst_twiddle_rsc_0_13_i_qa_d <= twiddle_rsc_0_13_i_qa_d;
  twiddle_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_twiddle_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_rsc_0_14_i_adra_d <= peaseNTT_core_inst_twiddle_rsc_0_14_i_adra_d;
  peaseNTT_core_inst_twiddle_rsc_0_14_i_qa_d <= twiddle_rsc_0_14_i_qa_d;
  twiddle_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_twiddle_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_rsc_0_15_i_adra_d <= peaseNTT_core_inst_twiddle_rsc_0_15_i_adra_d;
  peaseNTT_core_inst_twiddle_rsc_0_15_i_qa_d <= twiddle_rsc_0_15_i_qa_d;
  twiddle_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_twiddle_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_h_rsc_0_0_i_adra_d <= peaseNTT_core_inst_twiddle_h_rsc_0_0_i_adra_d;
  peaseNTT_core_inst_twiddle_h_rsc_0_0_i_qa_d <= twiddle_h_rsc_0_0_i_qa_d;
  twiddle_h_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_twiddle_h_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_h_rsc_0_1_i_adra_d <= peaseNTT_core_inst_twiddle_h_rsc_0_1_i_adra_d;
  peaseNTT_core_inst_twiddle_h_rsc_0_1_i_qa_d <= twiddle_h_rsc_0_1_i_qa_d;
  twiddle_h_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_twiddle_h_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_h_rsc_0_2_i_adra_d <= peaseNTT_core_inst_twiddle_h_rsc_0_2_i_adra_d;
  peaseNTT_core_inst_twiddle_h_rsc_0_2_i_qa_d <= twiddle_h_rsc_0_2_i_qa_d;
  twiddle_h_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_twiddle_h_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_h_rsc_0_3_i_adra_d <= peaseNTT_core_inst_twiddle_h_rsc_0_3_i_adra_d;
  peaseNTT_core_inst_twiddle_h_rsc_0_3_i_qa_d <= twiddle_h_rsc_0_3_i_qa_d;
  twiddle_h_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_twiddle_h_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_h_rsc_0_4_i_adra_d <= peaseNTT_core_inst_twiddle_h_rsc_0_4_i_adra_d;
  peaseNTT_core_inst_twiddle_h_rsc_0_4_i_qa_d <= twiddle_h_rsc_0_4_i_qa_d;
  twiddle_h_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_twiddle_h_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_h_rsc_0_5_i_adra_d <= peaseNTT_core_inst_twiddle_h_rsc_0_5_i_adra_d;
  peaseNTT_core_inst_twiddle_h_rsc_0_5_i_qa_d <= twiddle_h_rsc_0_5_i_qa_d;
  twiddle_h_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_twiddle_h_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_h_rsc_0_6_i_adra_d <= peaseNTT_core_inst_twiddle_h_rsc_0_6_i_adra_d;
  peaseNTT_core_inst_twiddle_h_rsc_0_6_i_qa_d <= twiddle_h_rsc_0_6_i_qa_d;
  twiddle_h_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_twiddle_h_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_h_rsc_0_7_i_adra_d <= peaseNTT_core_inst_twiddle_h_rsc_0_7_i_adra_d;
  peaseNTT_core_inst_twiddle_h_rsc_0_7_i_qa_d <= twiddle_h_rsc_0_7_i_qa_d;
  twiddle_h_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_twiddle_h_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_h_rsc_0_8_i_adra_d <= peaseNTT_core_inst_twiddle_h_rsc_0_8_i_adra_d;
  peaseNTT_core_inst_twiddle_h_rsc_0_8_i_qa_d <= twiddle_h_rsc_0_8_i_qa_d;
  twiddle_h_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_twiddle_h_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_h_rsc_0_9_i_adra_d <= peaseNTT_core_inst_twiddle_h_rsc_0_9_i_adra_d;
  peaseNTT_core_inst_twiddle_h_rsc_0_9_i_qa_d <= twiddle_h_rsc_0_9_i_qa_d;
  twiddle_h_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_twiddle_h_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_h_rsc_0_10_i_adra_d <= peaseNTT_core_inst_twiddle_h_rsc_0_10_i_adra_d;
  peaseNTT_core_inst_twiddle_h_rsc_0_10_i_qa_d <= twiddle_h_rsc_0_10_i_qa_d;
  twiddle_h_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_twiddle_h_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_h_rsc_0_11_i_adra_d <= peaseNTT_core_inst_twiddle_h_rsc_0_11_i_adra_d;
  peaseNTT_core_inst_twiddle_h_rsc_0_11_i_qa_d <= twiddle_h_rsc_0_11_i_qa_d;
  twiddle_h_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_twiddle_h_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_h_rsc_0_12_i_adra_d <= peaseNTT_core_inst_twiddle_h_rsc_0_12_i_adra_d;
  peaseNTT_core_inst_twiddle_h_rsc_0_12_i_qa_d <= twiddle_h_rsc_0_12_i_qa_d;
  twiddle_h_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_twiddle_h_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_h_rsc_0_13_i_adra_d <= peaseNTT_core_inst_twiddle_h_rsc_0_13_i_adra_d;
  peaseNTT_core_inst_twiddle_h_rsc_0_13_i_qa_d <= twiddle_h_rsc_0_13_i_qa_d;
  twiddle_h_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_twiddle_h_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_h_rsc_0_14_i_adra_d <= peaseNTT_core_inst_twiddle_h_rsc_0_14_i_adra_d;
  peaseNTT_core_inst_twiddle_h_rsc_0_14_i_qa_d <= twiddle_h_rsc_0_14_i_qa_d;
  twiddle_h_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_twiddle_h_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_h_rsc_0_15_i_adra_d <= peaseNTT_core_inst_twiddle_h_rsc_0_15_i_adra_d;
  peaseNTT_core_inst_twiddle_h_rsc_0_15_i_qa_d <= twiddle_h_rsc_0_15_i_qa_d;
  twiddle_h_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_twiddle_h_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yt_rsc_0_0_i_d_d_iff <= peaseNTT_core_inst_yt_rsc_0_0_i_d_d_pff;
  yt_rsc_0_0_i_radr_d_iff <= peaseNTT_core_inst_yt_rsc_0_0_i_radr_d_pff;
  yt_rsc_0_0_i_wadr_d_iff <= peaseNTT_core_inst_yt_rsc_0_0_i_wadr_d_pff;
  yt_rsc_0_1_i_d_d_iff <= peaseNTT_core_inst_yt_rsc_0_1_i_d_d_pff;
  yt_rsc_0_1_i_wadr_d_iff <= peaseNTT_core_inst_yt_rsc_0_1_i_wadr_d_pff;
  yt_rsc_0_2_i_d_d_iff <= peaseNTT_core_inst_yt_rsc_0_2_i_d_d_pff;
  yt_rsc_0_2_i_wadr_d_iff <= peaseNTT_core_inst_yt_rsc_0_2_i_wadr_d_pff;
  yt_rsc_0_3_i_d_d_iff <= peaseNTT_core_inst_yt_rsc_0_3_i_d_d_pff;
  yt_rsc_0_3_i_wadr_d_iff <= peaseNTT_core_inst_yt_rsc_0_3_i_wadr_d_pff;
  yt_rsc_0_4_i_d_d_iff <= peaseNTT_core_inst_yt_rsc_0_4_i_d_d_pff;
  yt_rsc_0_4_i_wadr_d_iff <= peaseNTT_core_inst_yt_rsc_0_4_i_wadr_d_pff;
  yt_rsc_0_5_i_d_d_iff <= peaseNTT_core_inst_yt_rsc_0_5_i_d_d_pff;
  yt_rsc_0_5_i_wadr_d_iff <= peaseNTT_core_inst_yt_rsc_0_5_i_wadr_d_pff;
  yt_rsc_0_6_i_d_d_iff <= peaseNTT_core_inst_yt_rsc_0_6_i_d_d_pff;
  yt_rsc_0_6_i_wadr_d_iff <= peaseNTT_core_inst_yt_rsc_0_6_i_wadr_d_pff;
  yt_rsc_0_7_i_d_d_iff <= peaseNTT_core_inst_yt_rsc_0_7_i_d_d_pff;
  yt_rsc_0_8_i_d_d_iff <= peaseNTT_core_inst_yt_rsc_0_8_i_d_d_pff;
  yt_rsc_0_9_i_d_d_iff <= peaseNTT_core_inst_yt_rsc_0_9_i_d_d_pff;
  yt_rsc_0_10_i_d_d_iff <= peaseNTT_core_inst_yt_rsc_0_10_i_d_d_pff;
  yt_rsc_0_10_i_wadr_d_iff <= peaseNTT_core_inst_yt_rsc_0_10_i_wadr_d_pff;
  yt_rsc_0_11_i_d_d_iff <= peaseNTT_core_inst_yt_rsc_0_11_i_d_d_pff;
  yt_rsc_0_11_i_wadr_d_iff <= peaseNTT_core_inst_yt_rsc_0_11_i_wadr_d_pff;
  yt_rsc_0_12_i_d_d_iff <= peaseNTT_core_inst_yt_rsc_0_12_i_d_d_pff;
  yt_rsc_0_13_i_d_d_iff <= peaseNTT_core_inst_yt_rsc_0_13_i_d_d_pff;
  yt_rsc_0_14_i_d_d_iff <= peaseNTT_core_inst_yt_rsc_0_14_i_d_d_pff;
  yt_rsc_0_15_i_d_d_iff <= peaseNTT_core_inst_yt_rsc_0_15_i_d_d_pff;
  yt_rsc_4_0_i_d_d_iff <= peaseNTT_core_inst_yt_rsc_4_0_i_d_d_pff;
  yt_rsc_4_0_i_wadr_d_iff <= peaseNTT_core_inst_yt_rsc_4_0_i_wadr_d_pff;
  yt_rsc_4_1_i_d_d_iff <= peaseNTT_core_inst_yt_rsc_4_1_i_d_d_pff;
  yt_rsc_4_1_i_wadr_d_iff <= peaseNTT_core_inst_yt_rsc_4_1_i_wadr_d_pff;
  yt_rsc_4_2_i_d_d_iff <= peaseNTT_core_inst_yt_rsc_4_2_i_d_d_pff;
  yt_rsc_4_2_i_wadr_d_iff <= peaseNTT_core_inst_yt_rsc_4_2_i_wadr_d_pff;
  yt_rsc_4_3_i_d_d_iff <= peaseNTT_core_inst_yt_rsc_4_3_i_d_d_pff;
  yt_rsc_4_3_i_wadr_d_iff <= peaseNTT_core_inst_yt_rsc_4_3_i_wadr_d_pff;
  yt_rsc_4_4_i_d_d_iff <= peaseNTT_core_inst_yt_rsc_4_4_i_d_d_pff;
  yt_rsc_4_4_i_wadr_d_iff <= peaseNTT_core_inst_yt_rsc_4_4_i_wadr_d_pff;
  yt_rsc_4_5_i_d_d_iff <= peaseNTT_core_inst_yt_rsc_4_5_i_d_d_pff;
  yt_rsc_4_5_i_wadr_d_iff <= peaseNTT_core_inst_yt_rsc_4_5_i_wadr_d_pff;
  yt_rsc_4_6_i_d_d_iff <= peaseNTT_core_inst_yt_rsc_4_6_i_d_d_pff;
  yt_rsc_4_6_i_wadr_d_iff <= peaseNTT_core_inst_yt_rsc_4_6_i_wadr_d_pff;
  yt_rsc_4_7_i_d_d_iff <= peaseNTT_core_inst_yt_rsc_4_7_i_d_d_pff;
  yt_rsc_4_8_i_d_d_iff <= peaseNTT_core_inst_yt_rsc_4_8_i_d_d_pff;
  yt_rsc_4_9_i_d_d_iff <= peaseNTT_core_inst_yt_rsc_4_9_i_d_d_pff;
  yt_rsc_4_9_i_wadr_d_iff <= peaseNTT_core_inst_yt_rsc_4_9_i_wadr_d_pff;
  yt_rsc_4_10_i_d_d_iff <= peaseNTT_core_inst_yt_rsc_4_10_i_d_d_pff;
  yt_rsc_4_10_i_wadr_d_iff <= peaseNTT_core_inst_yt_rsc_4_10_i_wadr_d_pff;
  yt_rsc_4_11_i_d_d_iff <= peaseNTT_core_inst_yt_rsc_4_11_i_d_d_pff;
  yt_rsc_4_11_i_wadr_d_iff <= peaseNTT_core_inst_yt_rsc_4_11_i_wadr_d_pff;
  yt_rsc_4_12_i_d_d_iff <= peaseNTT_core_inst_yt_rsc_4_12_i_d_d_pff;
  yt_rsc_4_13_i_d_d_iff <= peaseNTT_core_inst_yt_rsc_4_13_i_d_d_pff;
  yt_rsc_4_14_i_d_d_iff <= peaseNTT_core_inst_yt_rsc_4_14_i_d_d_pff;
  yt_rsc_4_15_i_d_d_iff <= peaseNTT_core_inst_yt_rsc_4_15_i_d_d_pff;
  xt_rsc_0_0_i_adra_d_iff <= peaseNTT_core_inst_xt_rsc_0_0_i_adra_d_pff;
  xt_rsc_0_0_i_da_d_iff <= peaseNTT_core_inst_xt_rsc_0_0_i_da_d_pff;
  xt_rsc_0_1_i_adra_d_iff <= peaseNTT_core_inst_xt_rsc_0_1_i_adra_d_pff;
  xt_rsc_0_1_i_da_d_iff <= peaseNTT_core_inst_xt_rsc_0_1_i_da_d_pff;
  xt_rsc_0_2_i_adra_d_iff <= peaseNTT_core_inst_xt_rsc_0_2_i_adra_d_pff;
  xt_rsc_0_2_i_da_d_iff <= peaseNTT_core_inst_xt_rsc_0_2_i_da_d_pff;
  xt_rsc_0_3_i_adra_d_iff <= peaseNTT_core_inst_xt_rsc_0_3_i_adra_d_pff;
  xt_rsc_0_3_i_da_d_iff <= peaseNTT_core_inst_xt_rsc_0_3_i_da_d_pff;
  xt_rsc_0_4_i_adra_d_iff <= peaseNTT_core_inst_xt_rsc_0_4_i_adra_d_pff;
  xt_rsc_0_4_i_da_d_iff <= peaseNTT_core_inst_xt_rsc_0_4_i_da_d_pff;
  xt_rsc_0_5_i_adra_d_iff <= peaseNTT_core_inst_xt_rsc_0_5_i_adra_d_pff;
  xt_rsc_0_5_i_da_d_iff <= peaseNTT_core_inst_xt_rsc_0_5_i_da_d_pff;
  xt_rsc_0_6_i_adra_d_iff <= peaseNTT_core_inst_xt_rsc_0_6_i_adra_d_pff;
  xt_rsc_0_6_i_da_d_iff <= peaseNTT_core_inst_xt_rsc_0_6_i_da_d_pff;
  xt_rsc_0_7_i_adra_d_iff <= peaseNTT_core_inst_xt_rsc_0_7_i_adra_d_pff;
  xt_rsc_0_7_i_da_d_iff <= peaseNTT_core_inst_xt_rsc_0_7_i_da_d_pff;
  xt_rsc_0_8_i_adra_d_iff <= peaseNTT_core_inst_xt_rsc_0_8_i_adra_d_pff;
  xt_rsc_0_8_i_da_d_iff <= peaseNTT_core_inst_xt_rsc_0_8_i_da_d_pff;
  xt_rsc_0_9_i_adra_d_iff <= peaseNTT_core_inst_xt_rsc_0_9_i_adra_d_pff;
  xt_rsc_0_9_i_da_d_iff <= peaseNTT_core_inst_xt_rsc_0_9_i_da_d_pff;
  xt_rsc_0_10_i_adra_d_iff <= peaseNTT_core_inst_xt_rsc_0_10_i_adra_d_pff;
  xt_rsc_0_10_i_da_d_iff <= peaseNTT_core_inst_xt_rsc_0_10_i_da_d_pff;
  xt_rsc_0_11_i_adra_d_iff <= peaseNTT_core_inst_xt_rsc_0_11_i_adra_d_pff;
  xt_rsc_0_11_i_da_d_iff <= peaseNTT_core_inst_xt_rsc_0_11_i_da_d_pff;
  xt_rsc_0_12_i_adra_d_iff <= peaseNTT_core_inst_xt_rsc_0_12_i_adra_d_pff;
  xt_rsc_0_12_i_da_d_iff <= peaseNTT_core_inst_xt_rsc_0_12_i_da_d_pff;
  xt_rsc_0_13_i_adra_d_iff <= peaseNTT_core_inst_xt_rsc_0_13_i_adra_d_pff;
  xt_rsc_0_13_i_da_d_iff <= peaseNTT_core_inst_xt_rsc_0_13_i_da_d_pff;
  xt_rsc_0_14_i_adra_d_iff <= peaseNTT_core_inst_xt_rsc_0_14_i_adra_d_pff;
  xt_rsc_0_14_i_da_d_iff <= peaseNTT_core_inst_xt_rsc_0_14_i_da_d_pff;
  xt_rsc_0_15_i_adra_d_iff <= peaseNTT_core_inst_xt_rsc_0_15_i_adra_d_pff;
  xt_rsc_0_15_i_da_d_iff <= peaseNTT_core_inst_xt_rsc_0_15_i_da_d_pff;
  xt_rsc_4_0_i_da_d_iff <= peaseNTT_core_inst_xt_rsc_4_0_i_da_d_pff;
  xt_rsc_4_1_i_adra_d_iff <= peaseNTT_core_inst_xt_rsc_4_1_i_adra_d_pff;
  xt_rsc_4_1_i_da_d_iff <= peaseNTT_core_inst_xt_rsc_4_1_i_da_d_pff;
  xt_rsc_4_2_i_adra_d_iff <= peaseNTT_core_inst_xt_rsc_4_2_i_adra_d_pff;
  xt_rsc_4_2_i_da_d_iff <= peaseNTT_core_inst_xt_rsc_4_2_i_da_d_pff;
  xt_rsc_4_3_i_da_d_iff <= peaseNTT_core_inst_xt_rsc_4_3_i_da_d_pff;
  xt_rsc_4_4_i_da_d_iff <= peaseNTT_core_inst_xt_rsc_4_4_i_da_d_pff;
  xt_rsc_4_5_i_da_d_iff <= peaseNTT_core_inst_xt_rsc_4_5_i_da_d_pff;
  xt_rsc_4_6_i_da_d_iff <= peaseNTT_core_inst_xt_rsc_4_6_i_da_d_pff;
  xt_rsc_4_7_i_da_d_iff <= peaseNTT_core_inst_xt_rsc_4_7_i_da_d_pff;
  xt_rsc_4_8_i_da_d_iff <= peaseNTT_core_inst_xt_rsc_4_8_i_da_d_pff;
  xt_rsc_4_9_i_adra_d_iff <= peaseNTT_core_inst_xt_rsc_4_9_i_adra_d_pff;
  xt_rsc_4_9_i_da_d_iff <= peaseNTT_core_inst_xt_rsc_4_9_i_da_d_pff;
  xt_rsc_4_10_i_adra_d_iff <= peaseNTT_core_inst_xt_rsc_4_10_i_adra_d_pff;
  xt_rsc_4_10_i_da_d_iff <= peaseNTT_core_inst_xt_rsc_4_10_i_da_d_pff;
  xt_rsc_4_11_i_da_d_iff <= peaseNTT_core_inst_xt_rsc_4_11_i_da_d_pff;
  xt_rsc_4_12_i_da_d_iff <= peaseNTT_core_inst_xt_rsc_4_12_i_da_d_pff;
  xt_rsc_4_13_i_da_d_iff <= peaseNTT_core_inst_xt_rsc_4_13_i_da_d_pff;
  xt_rsc_4_14_i_da_d_iff <= peaseNTT_core_inst_xt_rsc_4_14_i_da_d_pff;
  xt_rsc_4_15_i_da_d_iff <= peaseNTT_core_inst_xt_rsc_4_15_i_da_d_pff;

END v14;



