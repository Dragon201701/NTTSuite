
--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/ccs_in_v1.vhd 
--------------------------------------------------------------------------------
-- Catapult Synthesis - Sample I/O Port Library
--
-- Copyright (c) 2003-2017 Mentor Graphics Corp.
--       All Rights Reserved
--
-- This document may be used and distributed without restriction provided that
-- this copyright statement is not removed from the file and that any derivative
-- work contains this copyright notice.
--
-- The design information contained in this file is intended to be an example
-- of the functionality which the end user may study in preparation for creating
-- their own custom interfaces. This design does not necessarily present a 
-- complete implementation of the named protocol or standard.
--
--------------------------------------------------------------------------------

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;

PACKAGE ccs_in_pkg_v1 IS

COMPONENT ccs_in_v1
  GENERIC (
    rscid    : INTEGER;
    width    : INTEGER
  );
  PORT (
    idat   : OUT std_logic_vector(width-1 DOWNTO 0);
    dat    : IN  std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

END ccs_in_pkg_v1;

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all; -- Prevent STARC 2.1.1.2 violation

ENTITY ccs_in_v1 IS
  GENERIC (
    rscid : INTEGER;
    width : INTEGER
  );
  PORT (
    idat  : OUT std_logic_vector(width-1 DOWNTO 0);
    dat   : IN  std_logic_vector(width-1 DOWNTO 0)
  );
END ccs_in_v1;

ARCHITECTURE beh OF ccs_in_v1 IS
BEGIN

  idat <= dat;

END beh;


--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_io_sync_v2.vhd 
--------------------------------------------------------------------------------
-- Catapult Synthesis - Sample I/O Port Library
--
-- Copyright (c) 2003-2017 Mentor Graphics Corp.
--       All Rights Reserved
--
-- This document may be used and distributed without restriction provided that
-- this copyright statement is not removed from the file and that any derivative
-- work contains this copyright notice.
--
-- The design information contained in this file is intended to be an example
-- of the functionality which the end user may study in preparation for creating
-- their own custom interfaces. This design does not necessarily present a 
-- complete implementation of the named protocol or standard.
--
--------------------------------------------------------------------------------

LIBRARY ieee;

USE ieee.std_logic_1164.all;
PACKAGE mgc_io_sync_pkg_v2 IS

COMPONENT mgc_io_sync_v2
  GENERIC (
    valid    : INTEGER RANGE 0 TO 1
  );
  PORT (
    ld       : IN    std_logic;
    lz       : OUT   std_logic
  );
END COMPONENT;

END mgc_io_sync_pkg_v2;

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all; -- Prevent STARC 2.1.1.2 violation

ENTITY mgc_io_sync_v2 IS
  GENERIC (
    valid    : INTEGER RANGE 0 TO 1
  );
  PORT (
    ld       : IN    std_logic;
    lz       : OUT   std_logic
  );
END mgc_io_sync_v2;

ARCHITECTURE beh OF mgc_io_sync_v2 IS
BEGIN

  lz <= ld;

END beh;


--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/src/funcs.vhd 

-- a package of attributes that give verification tools a hint about
-- the function being implemented
PACKAGE attributes IS
  ATTRIBUTE CALYPTO_FUNC : string;
  ATTRIBUTE CALYPTO_DATA_ORDER : string;
end attributes;

-----------------------------------------------------------------------
-- Package that declares synthesizable functions needed for RTL output
-----------------------------------------------------------------------

LIBRARY ieee;

use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;

PACKAGE funcs IS

-----------------------------------------------------------------
-- utility functions
-----------------------------------------------------------------

   FUNCTION TO_STDLOGIC(arg1: BOOLEAN) RETURN STD_LOGIC;
--   FUNCTION TO_STDLOGIC(arg1: STD_ULOGIC_VECTOR(0 DOWNTO 0)) RETURN STD_LOGIC;
   FUNCTION TO_STDLOGIC(arg1: STD_LOGIC_VECTOR(0 DOWNTO 0)) RETURN STD_LOGIC;
   FUNCTION TO_STDLOGIC(arg1: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION TO_STDLOGIC(arg1: SIGNED(0 DOWNTO 0)) RETURN STD_LOGIC;
   FUNCTION TO_STDLOGICVECTOR(arg1: STD_LOGIC) RETURN STD_LOGIC_VECTOR;

   FUNCTION maximum(arg1, arg2 : INTEGER) RETURN INTEGER;
   FUNCTION minimum(arg1, arg2 : INTEGER) RETURN INTEGER;
   FUNCTION ifeqsel(arg1, arg2, seleq, selne : INTEGER) RETURN INTEGER;
   FUNCTION resolve_std_logic_vector(input1: STD_LOGIC_VECTOR; input2 : STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR;
   
-----------------------------------------------------------------
-- logic functions
-----------------------------------------------------------------

   FUNCTION and_s(inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC;
   FUNCTION or_s (inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC;
   FUNCTION xor_s(inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC;

   FUNCTION and_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR;
   FUNCTION or_v (inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR;
   FUNCTION xor_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR;

-----------------------------------------------------------------
-- mux functions
-----------------------------------------------------------------

   FUNCTION mux_s(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC       ) RETURN STD_LOGIC;
   FUNCTION mux_s(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR) RETURN STD_LOGIC;
   FUNCTION mux_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC       ) RETURN STD_LOGIC_VECTOR;
   FUNCTION mux_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR;

-----------------------------------------------------------------
-- latch functions
-----------------------------------------------------------------
   FUNCTION lat_s(dinput: STD_LOGIC       ; clk: STD_LOGIC; doutput: STD_LOGIC       ) RETURN STD_LOGIC;
   FUNCTION lat_v(dinput: STD_LOGIC_VECTOR; clk: STD_LOGIC; doutput: STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR;

-----------------------------------------------------------------
-- tristate functions
-----------------------------------------------------------------
--   FUNCTION tri_s(dinput: STD_LOGIC       ; control: STD_LOGIC) RETURN STD_LOGIC;
--   FUNCTION tri_v(dinput: STD_LOGIC_VECTOR; control: STD_LOGIC) RETURN STD_LOGIC_VECTOR;

-----------------------------------------------------------------
-- compare functions returning STD_LOGIC
-- in contrast to the functions returning boolean
-----------------------------------------------------------------

   FUNCTION "=" (l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION "=" (l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION "/="(l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION "/="(l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION "<="(l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION "<="(l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION "<" (l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION "<" (l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION ">="(l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION ">="(l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION ">" (l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION ">" (l, r: SIGNED  ) RETURN STD_LOGIC;

   -- RETURN 2 bits (left => lt, right => eq)
   FUNCTION cmp (l, r: STD_LOGIC_VECTOR) RETURN STD_LOGIC;

-----------------------------------------------------------------
-- Vectorized Overloaded Arithmetic Operators
-----------------------------------------------------------------

   FUNCTION faccu(arg: UNSIGNED; width: NATURAL) RETURN UNSIGNED;
 
   FUNCTION fabs(arg1: SIGNED  ) RETURN UNSIGNED;

   FUNCTION "/"  (l, r: UNSIGNED) RETURN UNSIGNED;
   FUNCTION "MOD"(l, r: UNSIGNED) RETURN UNSIGNED;
   FUNCTION "REM"(l, r: UNSIGNED) RETURN UNSIGNED;
   FUNCTION "**" (l, r: UNSIGNED) RETURN UNSIGNED;

   FUNCTION "/"  (l, r: SIGNED  ) RETURN SIGNED  ;
   FUNCTION "MOD"(l, r: SIGNED  ) RETURN SIGNED  ;
   FUNCTION "REM"(l, r: SIGNED  ) RETURN SIGNED  ;
   FUNCTION "**" (l, r: SIGNED  ) RETURN SIGNED  ;

-----------------------------------------------------------------
--               S H I F T   F U C T I O N S
-- negative shift shifts the opposite direction
-- *_stdar functions use shift functions from std_logic_arith
-----------------------------------------------------------------

   FUNCTION fshl(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshl(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED;

   FUNCTION fshl(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshr(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshl(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshr(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED  ;

   FUNCTION fshl(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshl(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;

   FUNCTION frot(arg1: STD_LOGIC_VECTOR; arg2: STD_LOGIC_VECTOR; signd2: BOOLEAN; sdir: INTEGER range -1 TO 1) RETURN STD_LOGIC_VECTOR;
   FUNCTION frol(arg1: STD_LOGIC_VECTOR; arg2: UNSIGNED) RETURN STD_LOGIC_VECTOR;
   FUNCTION fror(arg1: STD_LOGIC_VECTOR; arg2: UNSIGNED) RETURN STD_LOGIC_VECTOR;
   FUNCTION frol(arg1: STD_LOGIC_VECTOR; arg2: SIGNED  ) RETURN STD_LOGIC_VECTOR;
   FUNCTION fror(arg1: STD_LOGIC_VECTOR; arg2: SIGNED  ) RETURN STD_LOGIC_VECTOR;

   -----------------------------------------------------------------
   -- *_stdar functions use shift functions from std_logic_arith
   -----------------------------------------------------------------
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED;

   FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshr_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshr_stdar(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED  ;

   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;

-----------------------------------------------------------------
-- indexing functions: LSB always has index 0
-----------------------------------------------------------------

   FUNCTION readindex(vec: STD_LOGIC_VECTOR; index: INTEGER                 ) RETURN STD_LOGIC;
   FUNCTION readslice(vec: STD_LOGIC_VECTOR; index: INTEGER; width: POSITIVE) RETURN STD_LOGIC_VECTOR;

   FUNCTION writeindex(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC       ; index: INTEGER) RETURN STD_LOGIC_VECTOR;
   FUNCTION n_bits(p: NATURAL) RETURN POSITIVE;
   --FUNCTION writeslice(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC_VECTOR; index: INTEGER) RETURN STD_LOGIC_VECTOR;
   FUNCTION writeslice(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC_VECTOR; enable: STD_LOGIC_VECTOR; byte_width: INTEGER;  index: INTEGER) RETURN STD_LOGIC_VECTOR ;

   FUNCTION ceil_log2(size : NATURAL) return NATURAL;
   FUNCTION bits(size : NATURAL) return NATURAL;    

   PROCEDURE csa(a, b, c: IN INTEGER; s, cout: OUT STD_LOGIC_VECTOR);
   PROCEDURE csha(a, b: IN INTEGER; s, cout: OUT STD_LOGIC_VECTOR);
   
END funcs;


--------------------------- B O D Y ----------------------------


PACKAGE BODY funcs IS

-----------------------------------------------------------------
-- utility functions
-----------------------------------------------------------------

   FUNCTION TO_STDLOGIC(arg1: BOOLEAN) RETURN STD_LOGIC IS
     BEGIN IF arg1 THEN RETURN '1'; ELSE RETURN '0'; END IF; END;
--   FUNCTION TO_STDLOGIC(arg1: STD_ULOGIC_VECTOR(0 DOWNTO 0)) RETURN STD_LOGIC IS
--     BEGIN RETURN arg1(0); END;
   FUNCTION TO_STDLOGIC(arg1: STD_LOGIC_VECTOR(0 DOWNTO 0)) RETURN STD_LOGIC IS
     BEGIN RETURN arg1(0); END;
   FUNCTION TO_STDLOGIC(arg1: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN arg1(0); END;
   FUNCTION TO_STDLOGIC(arg1: SIGNED(0 DOWNTO 0)) RETURN STD_LOGIC IS
     BEGIN RETURN arg1(0); END;

   FUNCTION TO_STDLOGICVECTOR(arg1: STD_LOGIC) RETURN STD_LOGIC_VECTOR IS
     VARIABLE result: STD_LOGIC_VECTOR(0 DOWNTO 0);
   BEGIN
     result := (0 => arg1);
     RETURN result;
   END;

   FUNCTION maximum (arg1,arg2: INTEGER) RETURN INTEGER IS
   BEGIN
     IF(arg1 > arg2) THEN
       RETURN(arg1) ;
     ELSE
       RETURN(arg2) ;
     END IF;
   END;

   FUNCTION minimum (arg1,arg2: INTEGER) RETURN INTEGER IS
   BEGIN
     IF(arg1 < arg2) THEN
       RETURN(arg1) ;
     ELSE
       RETURN(arg2) ;
     END IF;
   END;

   FUNCTION ifeqsel(arg1, arg2, seleq, selne : INTEGER) RETURN INTEGER IS
   BEGIN
     IF(arg1 = arg2) THEN
       RETURN(seleq) ;
     ELSE
       RETURN(selne) ;
     END IF;
   END;

   FUNCTION resolve_std_logic_vector(input1: STD_LOGIC_VECTOR; input2: STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR IS
     CONSTANT len: INTEGER := input1'LENGTH;
     ALIAS input1a: STD_LOGIC_VECTOR(len-1 DOWNTO 0) IS input1;
     ALIAS input2a: STD_LOGIC_VECTOR(len-1 DOWNTO 0) IS input2;
     VARIABLE result: STD_LOGIC_VECTOR(len-1 DOWNTO 0);
   BEGIN
     result := (others => '0');
     --synopsys translate_off
     FOR i IN len-1 DOWNTO 0 LOOP
       result(i) := resolved(input1a(i) & input2a(i));
     END LOOP;
     --synopsys translate_on
     RETURN result;
   END;

   FUNCTION resolve_unsigned(input1: UNSIGNED; input2: UNSIGNED) RETURN UNSIGNED IS
   BEGIN RETURN UNSIGNED(resolve_std_logic_vector(STD_LOGIC_VECTOR(input1), STD_LOGIC_VECTOR(input2))); END;

   FUNCTION resolve_signed(input1: SIGNED; input2: SIGNED) RETURN SIGNED IS
   BEGIN RETURN SIGNED(resolve_std_logic_vector(STD_LOGIC_VECTOR(input1), STD_LOGIC_VECTOR(input2))); END;

-----------------------------------------------------------------
-- Logic Functions
-----------------------------------------------------------------

   FUNCTION "not"(arg1: UNSIGNED) RETURN UNSIGNED IS
     BEGIN RETURN UNSIGNED(not STD_LOGIC_VECTOR(arg1)); END;
   FUNCTION and_s(inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
     BEGIN RETURN TO_STDLOGIC(and_v(inputs, 1)); END;
   FUNCTION or_s (inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
     BEGIN RETURN TO_STDLOGIC(or_v(inputs, 1)); END;
   FUNCTION xor_s(inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
     BEGIN RETURN TO_STDLOGIC(xor_v(inputs, 1)); END;

   FUNCTION and_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR IS
     CONSTANT ilen: POSITIVE := inputs'LENGTH;
     CONSTANT ilenM1: POSITIVE := ilen-1; --2.1.6.3
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT ilenMolenM1: INTEGER := ilen-olen-1; --2.1.6.3
     VARIABLE inputsx: STD_LOGIC_VECTOR(ilen-1 DOWNTO 0);
     CONSTANT icnt2: POSITIVE:= inputs'LENGTH/olen;
     VARIABLE result: STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT ilen REM olen = 0 SEVERITY FAILURE;
     --synopsys translate_on
     inputsx := inputs;
     result := inputsx(olenM1 DOWNTO 0);
     FOR i IN icnt2-1 DOWNTO 1 LOOP
       inputsx(ilenMolenM1 DOWNTO 0) := inputsx(ilenM1 DOWNTO olen);
       result := result AND inputsx(olenM1 DOWNTO 0);
     END LOOP;
     RETURN result;
   END;

   FUNCTION or_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR IS
     CONSTANT ilen: POSITIVE := inputs'LENGTH;
     CONSTANT ilenM1: POSITIVE := ilen-1; --2.1.6.3
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT ilenMolenM1: INTEGER := ilen-olen-1; --2.1.6.3
     VARIABLE inputsx: STD_LOGIC_VECTOR(ilen-1 DOWNTO 0);
     CONSTANT icnt2: POSITIVE:= inputs'LENGTH/olen;
     VARIABLE result: STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT ilen REM olen = 0 SEVERITY FAILURE;
     --synopsys translate_on
     inputsx := inputs;
     result := inputsx(olenM1 DOWNTO 0);
     -- this if is added as a quick fix for a bug in catapult evaluating the loop even if inputs'LENGTH==1
     -- see dts0100971279
     IF icnt2 > 1 THEN
       FOR i IN icnt2-1 DOWNTO 1 LOOP
         inputsx(ilenMolenM1 DOWNTO 0) := inputsx(ilenM1 DOWNTO olen);
         result := result OR inputsx(olenM1 DOWNTO 0);
       END LOOP;
     END IF;
     RETURN result;
   END;

   FUNCTION xor_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR IS
     CONSTANT ilen: POSITIVE := inputs'LENGTH;
     CONSTANT ilenM1: POSITIVE := ilen-1; --2.1.6.3
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT ilenMolenM1: INTEGER := ilen-olen-1; --2.1.6.3
     VARIABLE inputsx: STD_LOGIC_VECTOR(ilen-1 DOWNTO 0);
     CONSTANT icnt2: POSITIVE:= inputs'LENGTH/olen;
     VARIABLE result: STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT ilen REM olen = 0 SEVERITY FAILURE;
     --synopsys translate_on
     inputsx := inputs;
     result := inputsx(olenM1 DOWNTO 0);
     FOR i IN icnt2-1 DOWNTO 1 LOOP
       inputsx(ilenMolenM1 DOWNTO 0) := inputsx(ilenM1 DOWNTO olen);
       result := result XOR inputsx(olenM1 DOWNTO 0);
     END LOOP;
     RETURN result;
   END;

-----------------------------------------------------------------
-- Muxes
-----------------------------------------------------------------
   
   FUNCTION mux_sel2_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(1 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 4;
     ALIAS    inputs0: STD_LOGIC_VECTOR( inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector( size-1 DOWNTO 0);
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "00" =>
       result := inputs0(1*size-1 DOWNTO 0*size);
     WHEN "01" =>
       result := inputs0(2*size-1 DOWNTO 1*size);
     WHEN "10" =>
       result := inputs0(3*size-1 DOWNTO 2*size);
     WHEN "11" =>
       result := inputs0(4*size-1 DOWNTO 3*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;
   
   FUNCTION mux_sel3_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(2 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 8;
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector(size-1 DOWNTO 0);
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "000" =>
       result := inputs0(1*size-1 DOWNTO 0*size);
     WHEN "001" =>
       result := inputs0(2*size-1 DOWNTO 1*size);
     WHEN "010" =>
       result := inputs0(3*size-1 DOWNTO 2*size);
     WHEN "011" =>
       result := inputs0(4*size-1 DOWNTO 3*size);
     WHEN "100" =>
       result := inputs0(5*size-1 DOWNTO 4*size);
     WHEN "101" =>
       result := inputs0(6*size-1 DOWNTO 5*size);
     WHEN "110" =>
       result := inputs0(7*size-1 DOWNTO 6*size);
     WHEN "111" =>
       result := inputs0(8*size-1 DOWNTO 7*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;
   
   FUNCTION mux_sel4_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(3 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 16;
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector(size-1 DOWNTO 0);
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "0000" =>
       result := inputs0( 1*size-1 DOWNTO 0*size);
     WHEN "0001" =>
       result := inputs0( 2*size-1 DOWNTO 1*size);
     WHEN "0010" =>
       result := inputs0( 3*size-1 DOWNTO 2*size);
     WHEN "0011" =>
       result := inputs0( 4*size-1 DOWNTO 3*size);
     WHEN "0100" =>
       result := inputs0( 5*size-1 DOWNTO 4*size);
     WHEN "0101" =>
       result := inputs0( 6*size-1 DOWNTO 5*size);
     WHEN "0110" =>
       result := inputs0( 7*size-1 DOWNTO 6*size);
     WHEN "0111" =>
       result := inputs0( 8*size-1 DOWNTO 7*size);
     WHEN "1000" =>
       result := inputs0( 9*size-1 DOWNTO 8*size);
     WHEN "1001" =>
       result := inputs0( 10*size-1 DOWNTO 9*size);
     WHEN "1010" =>
       result := inputs0( 11*size-1 DOWNTO 10*size);
     WHEN "1011" =>
       result := inputs0( 12*size-1 DOWNTO 11*size);
     WHEN "1100" =>
       result := inputs0( 13*size-1 DOWNTO 12*size);
     WHEN "1101" =>
       result := inputs0( 14*size-1 DOWNTO 13*size);
     WHEN "1110" =>
       result := inputs0( 15*size-1 DOWNTO 14*size);
     WHEN "1111" =>
       result := inputs0( 16*size-1 DOWNTO 15*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;
   
   FUNCTION mux_sel5_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(4 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 32;
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector(size-1 DOWNTO 0 );
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "00000" =>
       result := inputs0( 1*size-1 DOWNTO 0*size);
     WHEN "00001" =>
       result := inputs0( 2*size-1 DOWNTO 1*size);
     WHEN "00010" =>
       result := inputs0( 3*size-1 DOWNTO 2*size);
     WHEN "00011" =>
       result := inputs0( 4*size-1 DOWNTO 3*size);
     WHEN "00100" =>
       result := inputs0( 5*size-1 DOWNTO 4*size);
     WHEN "00101" =>
       result := inputs0( 6*size-1 DOWNTO 5*size);
     WHEN "00110" =>
       result := inputs0( 7*size-1 DOWNTO 6*size);
     WHEN "00111" =>
       result := inputs0( 8*size-1 DOWNTO 7*size);
     WHEN "01000" =>
       result := inputs0( 9*size-1 DOWNTO 8*size);
     WHEN "01001" =>
       result := inputs0( 10*size-1 DOWNTO 9*size);
     WHEN "01010" =>
       result := inputs0( 11*size-1 DOWNTO 10*size);
     WHEN "01011" =>
       result := inputs0( 12*size-1 DOWNTO 11*size);
     WHEN "01100" =>
       result := inputs0( 13*size-1 DOWNTO 12*size);
     WHEN "01101" =>
       result := inputs0( 14*size-1 DOWNTO 13*size);
     WHEN "01110" =>
       result := inputs0( 15*size-1 DOWNTO 14*size);
     WHEN "01111" =>
       result := inputs0( 16*size-1 DOWNTO 15*size);
     WHEN "10000" =>
       result := inputs0( 17*size-1 DOWNTO 16*size);
     WHEN "10001" =>
       result := inputs0( 18*size-1 DOWNTO 17*size);
     WHEN "10010" =>
       result := inputs0( 19*size-1 DOWNTO 18*size);
     WHEN "10011" =>
       result := inputs0( 20*size-1 DOWNTO 19*size);
     WHEN "10100" =>
       result := inputs0( 21*size-1 DOWNTO 20*size);
     WHEN "10101" =>
       result := inputs0( 22*size-1 DOWNTO 21*size);
     WHEN "10110" =>
       result := inputs0( 23*size-1 DOWNTO 22*size);
     WHEN "10111" =>
       result := inputs0( 24*size-1 DOWNTO 23*size);
     WHEN "11000" =>
       result := inputs0( 25*size-1 DOWNTO 24*size);
     WHEN "11001" =>
       result := inputs0( 26*size-1 DOWNTO 25*size);
     WHEN "11010" =>
       result := inputs0( 27*size-1 DOWNTO 26*size);
     WHEN "11011" =>
       result := inputs0( 28*size-1 DOWNTO 27*size);
     WHEN "11100" =>
       result := inputs0( 29*size-1 DOWNTO 28*size);
     WHEN "11101" =>
       result := inputs0( 30*size-1 DOWNTO 29*size);
     WHEN "11110" =>
       result := inputs0( 31*size-1 DOWNTO 30*size);
     WHEN "11111" =>
       result := inputs0( 32*size-1 DOWNTO 31*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;
   
   FUNCTION mux_sel6_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(5 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 64;
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector(size-1 DOWNTO 0);
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "000000" =>
       result := inputs0( 1*size-1 DOWNTO 0*size);
     WHEN "000001" =>
       result := inputs0( 2*size-1 DOWNTO 1*size);
     WHEN "000010" =>
       result := inputs0( 3*size-1 DOWNTO 2*size);
     WHEN "000011" =>
       result := inputs0( 4*size-1 DOWNTO 3*size);
     WHEN "000100" =>
       result := inputs0( 5*size-1 DOWNTO 4*size);
     WHEN "000101" =>
       result := inputs0( 6*size-1 DOWNTO 5*size);
     WHEN "000110" =>
       result := inputs0( 7*size-1 DOWNTO 6*size);
     WHEN "000111" =>
       result := inputs0( 8*size-1 DOWNTO 7*size);
     WHEN "001000" =>
       result := inputs0( 9*size-1 DOWNTO 8*size);
     WHEN "001001" =>
       result := inputs0( 10*size-1 DOWNTO 9*size);
     WHEN "001010" =>
       result := inputs0( 11*size-1 DOWNTO 10*size);
     WHEN "001011" =>
       result := inputs0( 12*size-1 DOWNTO 11*size);
     WHEN "001100" =>
       result := inputs0( 13*size-1 DOWNTO 12*size);
     WHEN "001101" =>
       result := inputs0( 14*size-1 DOWNTO 13*size);
     WHEN "001110" =>
       result := inputs0( 15*size-1 DOWNTO 14*size);
     WHEN "001111" =>
       result := inputs0( 16*size-1 DOWNTO 15*size);
     WHEN "010000" =>
       result := inputs0( 17*size-1 DOWNTO 16*size);
     WHEN "010001" =>
       result := inputs0( 18*size-1 DOWNTO 17*size);
     WHEN "010010" =>
       result := inputs0( 19*size-1 DOWNTO 18*size);
     WHEN "010011" =>
       result := inputs0( 20*size-1 DOWNTO 19*size);
     WHEN "010100" =>
       result := inputs0( 21*size-1 DOWNTO 20*size);
     WHEN "010101" =>
       result := inputs0( 22*size-1 DOWNTO 21*size);
     WHEN "010110" =>
       result := inputs0( 23*size-1 DOWNTO 22*size);
     WHEN "010111" =>
       result := inputs0( 24*size-1 DOWNTO 23*size);
     WHEN "011000" =>
       result := inputs0( 25*size-1 DOWNTO 24*size);
     WHEN "011001" =>
       result := inputs0( 26*size-1 DOWNTO 25*size);
     WHEN "011010" =>
       result := inputs0( 27*size-1 DOWNTO 26*size);
     WHEN "011011" =>
       result := inputs0( 28*size-1 DOWNTO 27*size);
     WHEN "011100" =>
       result := inputs0( 29*size-1 DOWNTO 28*size);
     WHEN "011101" =>
       result := inputs0( 30*size-1 DOWNTO 29*size);
     WHEN "011110" =>
       result := inputs0( 31*size-1 DOWNTO 30*size);
     WHEN "011111" =>
       result := inputs0( 32*size-1 DOWNTO 31*size);
     WHEN "100000" =>
       result := inputs0( 33*size-1 DOWNTO 32*size);
     WHEN "100001" =>
       result := inputs0( 34*size-1 DOWNTO 33*size);
     WHEN "100010" =>
       result := inputs0( 35*size-1 DOWNTO 34*size);
     WHEN "100011" =>
       result := inputs0( 36*size-1 DOWNTO 35*size);
     WHEN "100100" =>
       result := inputs0( 37*size-1 DOWNTO 36*size);
     WHEN "100101" =>
       result := inputs0( 38*size-1 DOWNTO 37*size);
     WHEN "100110" =>
       result := inputs0( 39*size-1 DOWNTO 38*size);
     WHEN "100111" =>
       result := inputs0( 40*size-1 DOWNTO 39*size);
     WHEN "101000" =>
       result := inputs0( 41*size-1 DOWNTO 40*size);
     WHEN "101001" =>
       result := inputs0( 42*size-1 DOWNTO 41*size);
     WHEN "101010" =>
       result := inputs0( 43*size-1 DOWNTO 42*size);
     WHEN "101011" =>
       result := inputs0( 44*size-1 DOWNTO 43*size);
     WHEN "101100" =>
       result := inputs0( 45*size-1 DOWNTO 44*size);
     WHEN "101101" =>
       result := inputs0( 46*size-1 DOWNTO 45*size);
     WHEN "101110" =>
       result := inputs0( 47*size-1 DOWNTO 46*size);
     WHEN "101111" =>
       result := inputs0( 48*size-1 DOWNTO 47*size);
     WHEN "110000" =>
       result := inputs0( 49*size-1 DOWNTO 48*size);
     WHEN "110001" =>
       result := inputs0( 50*size-1 DOWNTO 49*size);
     WHEN "110010" =>
       result := inputs0( 51*size-1 DOWNTO 50*size);
     WHEN "110011" =>
       result := inputs0( 52*size-1 DOWNTO 51*size);
     WHEN "110100" =>
       result := inputs0( 53*size-1 DOWNTO 52*size);
     WHEN "110101" =>
       result := inputs0( 54*size-1 DOWNTO 53*size);
     WHEN "110110" =>
       result := inputs0( 55*size-1 DOWNTO 54*size);
     WHEN "110111" =>
       result := inputs0( 56*size-1 DOWNTO 55*size);
     WHEN "111000" =>
       result := inputs0( 57*size-1 DOWNTO 56*size);
     WHEN "111001" =>
       result := inputs0( 58*size-1 DOWNTO 57*size);
     WHEN "111010" =>
       result := inputs0( 59*size-1 DOWNTO 58*size);
     WHEN "111011" =>
       result := inputs0( 60*size-1 DOWNTO 59*size);
     WHEN "111100" =>
       result := inputs0( 61*size-1 DOWNTO 60*size);
     WHEN "111101" =>
       result := inputs0( 62*size-1 DOWNTO 61*size);
     WHEN "111110" =>
       result := inputs0( 63*size-1 DOWNTO 62*size);
     WHEN "111111" =>
       result := inputs0( 64*size-1 DOWNTO 63*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;

   FUNCTION mux_s(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC) RETURN STD_LOGIC IS
   BEGIN RETURN TO_STDLOGIC(mux_v(inputs, sel)); END;

   FUNCTION mux_s(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
   BEGIN RETURN TO_STDLOGIC(mux_v(inputs, sel)); END;

   FUNCTION mux_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC) RETURN STD_LOGIC_VECTOR IS  --pragma hls_map_to_operator mux
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     CONSTANT size   : POSITIVE := inputs'LENGTH / 2;
     CONSTANT olen   : POSITIVE := inputs'LENGTH / 2;
     VARIABLE result : STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT inputs'LENGTH = olen * 2 SEVERITY FAILURE;
     --synopsys translate_on
       CASE sel IS
       WHEN '1'
     --synopsys translate_off
            | 'H'
     --synopsys translate_on
            =>
         result := inputs0( size-1 DOWNTO 0);
       WHEN '0' 
     --synopsys translate_off
            | 'L'
     --synopsys translate_on
            =>
         result := inputs0(2*size-1  DOWNTO size);
       WHEN others =>
         --synopsys translate_off
         result := resolve_std_logic_vector(inputs0(size-1 DOWNTO 0), inputs0( 2*size-1 DOWNTO size));
         --synopsys translate_on
       END CASE;
       RETURN result;
   END;
--   BEGIN RETURN mux_v(inputs, TO_STDLOGICVECTOR(sel)); END;

   FUNCTION mux_v(inputs: STD_LOGIC_VECTOR; sel : STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR IS --pragma hls_map_to_operator mux
     ALIAS    inputs0: STD_LOGIC_VECTOR( inputs'LENGTH-1 DOWNTO 0) IS inputs;
     ALIAS    sel0   : STD_LOGIC_VECTOR( sel'LENGTH-1 DOWNTO 0 ) IS sel;

     VARIABLE sellen : INTEGER RANGE 2-sel'LENGTH TO sel'LENGTH;
     CONSTANT size   : POSITIVE := inputs'LENGTH / 2;
     CONSTANT olen   : POSITIVE := inputs'LENGTH / 2**sel'LENGTH;
     VARIABLE result : STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
     TYPE inputs_array_type is array(natural range <>) of std_logic_vector( olen - 1 DOWNTO 0);
     VARIABLE inputs_array : inputs_array_type( 2**sel'LENGTH - 1 DOWNTO 0);
   BEGIN
     sellen := sel'LENGTH;
     --synopsys translate_off
     ASSERT inputs'LENGTH = olen * 2**sellen SEVERITY FAILURE;
     sellen := 2-sellen;
     --synopsys translate_on
     CASE sellen IS
     WHEN 1 =>
       CASE sel0(0) IS

       WHEN '1' 
     --synopsys translate_off
            | 'H'
     --synopsys translate_on
            =>
         result := inputs0(  size-1 DOWNTO 0);
       WHEN '0' 
     --synopsys translate_off
            | 'L'
     --synopsys translate_on
            =>
         result := inputs0(2*size-1 DOWNTO size);
       WHEN others =>
         --synopsys translate_off
         result := resolve_std_logic_vector(inputs0( size-1 DOWNTO 0), inputs0( 2*size-1 DOWNTO size));
         --synopsys translate_on
       END CASE;
     WHEN 2 =>
       result := mux_sel2_v(inputs, not sel);
     WHEN 3 =>
       result := mux_sel3_v(inputs, not sel);
     WHEN 4 =>
       result := mux_sel4_v(inputs, not sel);
     WHEN 5 =>
       result := mux_sel5_v(inputs, not sel);
     WHEN 6 =>
       result := mux_sel6_v(inputs, not sel);
     WHEN others =>
       -- synopsys translate_off
       IF(Is_X(sel0)) THEN
         result := (others => 'X');
       ELSE
       -- synopsys translate_on
         FOR i in 0 to 2**sel'LENGTH - 1 LOOP
           inputs_array(i) := inputs0( ((i + 1) * olen) - 1  DOWNTO i*olen);
         END LOOP;
         result := inputs_array(CONV_INTEGER( (UNSIGNED(NOT sel0)) ));
       -- synopsys translate_off
       END IF;
       -- synopsys translate_on
     END CASE;
     RETURN result;
   END;

 
-----------------------------------------------------------------
-- Latches
-----------------------------------------------------------------

   FUNCTION lat_s(dinput: STD_LOGIC; clk: STD_LOGIC; doutput: STD_LOGIC) RETURN STD_LOGIC IS
   BEGIN RETURN mux_s(STD_LOGIC_VECTOR'(doutput & dinput), clk); END;

   FUNCTION lat_v(dinput: STD_LOGIC_VECTOR ; clk: STD_LOGIC; doutput: STD_LOGIC_VECTOR ) RETURN STD_LOGIC_VECTOR IS
   BEGIN
     --synopsys translate_off
     ASSERT dinput'LENGTH = doutput'LENGTH SEVERITY FAILURE;
     --synopsys translate_on
     RETURN mux_v(doutput & dinput, clk);
   END;

-----------------------------------------------------------------
-- Tri-States
-----------------------------------------------------------------
--   FUNCTION tri_s(dinput: STD_LOGIC; control: STD_LOGIC) RETURN STD_LOGIC IS
--   BEGIN RETURN TO_STDLOGIC(tri_v(TO_STDLOGICVECTOR(dinput), control)); END;
--
--   FUNCTION tri_v(dinput: STD_LOGIC_VECTOR ; control: STD_LOGIC) RETURN STD_LOGIC_VECTOR IS
--     VARIABLE result: STD_LOGIC_VECTOR(dinput'range);
--   BEGIN
--     CASE control IS
--     WHEN '0' | 'L' =>
--       result := (others => 'Z');
--     WHEN '1' | 'H' =>
--       FOR i IN dinput'range LOOP
--         result(i) := to_UX01(dinput(i));
--       END LOOP;
--     WHEN others =>
--       -- synopsys translate_off
--       result := (others => 'X');
--       -- synopsys translate_on
--     END CASE;
--     RETURN result;
--   END;

-----------------------------------------------------------------
-- compare functions returning STD_LOGIC
-- in contrast to the functions returning boolean
-----------------------------------------------------------------

   FUNCTION "=" (l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN not or_s(STD_LOGIC_VECTOR(l) xor STD_LOGIC_VECTOR(r)); END;
   FUNCTION "=" (l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN not or_s(STD_LOGIC_VECTOR(l) xor STD_LOGIC_VECTOR(r)); END;
   FUNCTION "/="(l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN or_s(STD_LOGIC_VECTOR(l) xor STD_LOGIC_VECTOR(r)); END;
   FUNCTION "/="(l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN or_s(STD_LOGIC_VECTOR(l) xor STD_LOGIC_VECTOR(r)); END;

   FUNCTION "<" (l, r: UNSIGNED) RETURN STD_LOGIC IS
     VARIABLE diff: UNSIGNED(l'LENGTH DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT l'LENGTH = r'LENGTH SEVERITY FAILURE;
     --synopsys translate_on
     diff := ('0'&l) - ('0'&r);
     RETURN diff(l'LENGTH);
   END;
   FUNCTION "<"(l, r: SIGNED  ) RETURN STD_LOGIC IS
   BEGIN
     RETURN (UNSIGNED(l) < UNSIGNED(r)) xor (l(l'LEFT) xor r(r'LEFT));
   END;

   FUNCTION "<="(l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN not STD_LOGIC'(r < l); END;
   FUNCTION "<=" (l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN not STD_LOGIC'(r < l); END;
   FUNCTION ">" (l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN r < l; END;
   FUNCTION ">"(l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN r < l; END;
   FUNCTION ">="(l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN not STD_LOGIC'(l < r); END;
   FUNCTION ">=" (l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN not STD_LOGIC'(l < r); END;

   FUNCTION cmp (l, r: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
   BEGIN
     --synopsys translate_off
     ASSERT l'LENGTH = r'LENGTH SEVERITY FAILURE;
     --synopsys translate_on
     RETURN not or_s(l xor r);
   END;

-----------------------------------------------------------------
-- Vectorized Overloaded Arithmetic Operators
-----------------------------------------------------------------

   --some functions to placate spyglass
   FUNCTION mult_natural(a,b : NATURAL) RETURN NATURAL IS
   BEGIN
     return a*b;
   END mult_natural;

   FUNCTION div_natural(a,b : NATURAL) RETURN NATURAL IS
   BEGIN
     return a/b;
   END div_natural;

   FUNCTION mod_natural(a,b : NATURAL) RETURN NATURAL IS
   BEGIN
     return a mod b;
   END mod_natural;

   FUNCTION add_unsigned(a,b : UNSIGNED) RETURN UNSIGNED IS
   BEGIN
     return a+b;
   END add_unsigned;

   FUNCTION sub_unsigned(a,b : UNSIGNED) RETURN UNSIGNED IS
   BEGIN
     return a-b;
   END sub_unsigned;

   FUNCTION sub_int(a,b : INTEGER) RETURN INTEGER IS
   BEGIN
     return a-b;
   END sub_int;

   FUNCTION concat_0(b : UNSIGNED) RETURN UNSIGNED IS
   BEGIN
     return '0' & b;
   END concat_0;

   FUNCTION concat_uns(a,b : UNSIGNED) RETURN UNSIGNED IS
   BEGIN
     return a&b;
   END concat_uns;

   FUNCTION concat_vect(a,b : STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR IS
   BEGIN
     return a&b;
   END concat_vect;





   FUNCTION faccu(arg: UNSIGNED; width: NATURAL) RETURN UNSIGNED IS
     CONSTANT ninps : NATURAL := arg'LENGTH / width;
     ALIAS    arg0  : UNSIGNED(arg'LENGTH-1 DOWNTO 0) IS arg;
     VARIABLE result: UNSIGNED(width-1 DOWNTO 0);
     VARIABLE from  : INTEGER;
     VARIABLE dto   : INTEGER;
   BEGIN
     --synopsys translate_off
     ASSERT arg'LENGTH = width * ninps SEVERITY FAILURE;
     --synopsys translate_on
     result := (OTHERS => '0');
     FOR i IN ninps-1 DOWNTO 0 LOOP
       --result := result + arg0((i+1)*width-1 DOWNTO i*width);
       from := mult_natural((i+1), width)-1; --2.1.6.3
       dto  := mult_natural(i,width); --2.1.6.3
       result := add_unsigned(result , arg0(from DOWNTO dto) );
     END LOOP;
     RETURN result;
   END faccu;

   FUNCTION  fabs (arg1: SIGNED) RETURN UNSIGNED IS
   BEGIN
     CASE arg1(arg1'LEFT) IS
     WHEN '1'
     --synopsys translate_off
          | 'H'
     --synopsys translate_on
       =>
       RETURN UNSIGNED'("0") - UNSIGNED(arg1);
     WHEN '0'
     --synopsys translate_off
          | 'L'
     --synopsys translate_on
       =>
       RETURN UNSIGNED(arg1);
     WHEN others =>
       RETURN resolve_unsigned(UNSIGNED(arg1), UNSIGNED'("0") - UNSIGNED(arg1));
     END CASE;
   END;

   PROCEDURE divmod(l, r: UNSIGNED; rdiv, rmod: OUT UNSIGNED) IS
     CONSTANT llen: INTEGER := l'LENGTH;
     CONSTANT rlen: INTEGER := r'LENGTH;
     CONSTANT llen_plus_rlen: INTEGER := llen + rlen;
     VARIABLE lbuf: UNSIGNED(llen+rlen-1 DOWNTO 0);
     VARIABLE diff: UNSIGNED(rlen DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT rdiv'LENGTH = llen AND rmod'LENGTH = rlen SEVERITY FAILURE;
     --synopsys translate_on
     lbuf := (others => '0');
     lbuf(llen-1 DOWNTO 0) := l;
     FOR i IN rdiv'range LOOP
       diff := sub_unsigned(lbuf(llen_plus_rlen-1 DOWNTO llen-1) ,(concat_0(r)));
       rdiv(i) := not diff(rlen);
       IF diff(rlen) = '0' THEN
         lbuf(llen_plus_rlen-1 DOWNTO llen-1) := diff;
       END IF;
       lbuf(llen_plus_rlen-1 DOWNTO 1) := lbuf(llen_plus_rlen-2 DOWNTO 0);
     END LOOP;
     rmod := lbuf(llen_plus_rlen-1 DOWNTO llen);
   END divmod;

   FUNCTION "/"  (l, r: UNSIGNED) RETURN UNSIGNED IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
   BEGIN
     divmod(l, r, rdiv, rmod);
     RETURN rdiv;
   END "/";

   FUNCTION "MOD"(l, r: UNSIGNED) RETURN UNSIGNED IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
   BEGIN
     divmod(l, r, rdiv, rmod);
     RETURN rmod;
   END;

   FUNCTION "REM"(l, r: UNSIGNED) RETURN UNSIGNED IS
     BEGIN RETURN l MOD r; END;

   FUNCTION "/"  (l, r: SIGNED  ) RETURN SIGNED  IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
   BEGIN
     divmod(fabs(l), fabs(r), rdiv, rmod);
     IF to_X01(l(l'LEFT)) /= to_X01(r(r'LEFT)) THEN
       rdiv := UNSIGNED'("0") - rdiv;
     END IF;
     RETURN SIGNED(rdiv); -- overflow problem "1000" / "11"
   END "/";

   FUNCTION "MOD"(l, r: SIGNED  ) RETURN SIGNED  IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
     CONSTANT rnul: UNSIGNED(r'LENGTH-1 DOWNTO 0) := (others => '0');
   BEGIN
     divmod(fabs(l), fabs(r), rdiv, rmod);
     IF to_X01(l(l'LEFT)) = '1' THEN
       rmod := UNSIGNED'("0") - rmod;
     END IF;
     IF rmod /= rnul AND to_X01(l(l'LEFT)) /= to_X01(r(r'LEFT)) THEN
       rmod := UNSIGNED(r) + rmod;
     END IF;
     RETURN SIGNED(rmod);
   END "MOD";

   FUNCTION "REM"(l, r: SIGNED  ) RETURN SIGNED  IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
   BEGIN
     divmod(fabs(l), fabs(r), rdiv, rmod);
     IF to_X01(l(l'LEFT)) = '1' THEN
       rmod := UNSIGNED'("0") - rmod;
     END IF;
     RETURN SIGNED(rmod);
   END "REM";

   FUNCTION mult_unsigned(l,r : UNSIGNED) return UNSIGNED is
   BEGIN
     return l*r; 
   END mult_unsigned;

   FUNCTION "**" (l, r : UNSIGNED) RETURN UNSIGNED IS
     CONSTANT llen  : NATURAL := l'LENGTH;
     VARIABLE result: UNSIGNED(llen-1 DOWNTO 0);
     VARIABLE fak   : UNSIGNED(llen-1 DOWNTO 0);
   BEGIN
     fak := l;
     result := (others => '0'); result(0) := '1';
     FOR i IN r'reverse_range LOOP
       --was:result := UNSIGNED(mux_v(STD_LOGIC_VECTOR(result & (result*fak)), r(i)));
       result := UNSIGNED(mux_v(STD_LOGIC_VECTOR( concat_uns(result , mult_unsigned(result,fak) )), r(i)));

       fak := mult_unsigned(fak , fak);
     END LOOP;
     RETURN result;
   END "**";

   FUNCTION "**" (l, r : SIGNED) RETURN SIGNED IS
     CONSTANT rlen  : NATURAL := r'LENGTH;
     ALIAS    r0    : SIGNED(0 TO r'LENGTH-1) IS r;
     VARIABLE result: SIGNED(l'range);
   BEGIN
     CASE r(r'LEFT) IS
     WHEN '0'
   --synopsys translate_off
          | 'L'
   --synopsys translate_on
     =>
       result := SIGNED(UNSIGNED(l) ** UNSIGNED(r0(1 TO r'LENGTH-1)));
     WHEN '1'
   --synopsys translate_off
          | 'H'
   --synopsys translate_on
     =>
       result := (others => '0');
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END "**";

-----------------------------------------------------------------
--               S H I F T   F U C T I O N S
-- negative shift shifts the opposite direction
-----------------------------------------------------------------

   FUNCTION add_nat(arg1 : NATURAL; arg2 : NATURAL ) RETURN NATURAL IS
   BEGIN
     return (arg1 + arg2);
   END;
   
--   FUNCTION UNSIGNED_2_BIT_VECTOR(arg1 : NATURAL; arg2 : NATURAL ) RETURN BIT_VECTOR IS
--   BEGIN
--     return (arg1 + arg2);
--   END;
   
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
     CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
   BEGIN
     result := (others => sbit);
     result(ilenub DOWNTO 0) := arg1;
     result := shl(result, arg2);
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshl_stdar(arg1: SIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
     CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: SIGNED(len-1 DOWNTO 0);
   BEGIN
     result := (others => sbit);
     result(ilenub DOWNTO 0) := arg1;
     result := shl(SIGNED(result), arg2);
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
     CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
   BEGIN
     result := (others => sbit);
     result(ilenub DOWNTO 0) := arg1;
     result := shr(result, arg2);
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshr_stdar(arg1: SIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
     CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: SIGNED(len-1 DOWNTO 0);
   BEGIN
     result := (others => sbit);
     result(ilenub DOWNTO 0) := arg1;
     result := shr(result, arg2);
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT arg1l: NATURAL := arg1'LENGTH - 1;
     ALIAS    arg1x: UNSIGNED(arg1l DOWNTO 0) IS arg1;
     CONSTANT arg2l: NATURAL := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE arg1x_pad: UNSIGNED(arg1l+1 DOWNTO 0);
     VARIABLE result: UNSIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others=>'0');
     arg1x_pad(arg1l+1) := sbit;
     arg1x_pad(arg1l downto 0) := arg1x;
     IF arg2l = 0 THEN
       RETURN fshr_stdar(arg1x_pad, UNSIGNED(arg2x), sbit, olen);
     -- ELSIF arg1l = 0 THEN
     --   RETURN fshl(sbit & arg1x, arg2x, sbit, olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
     --synopsys translate_off
            | 'L'
     --synopsys translate_on
       =>
         RETURN fshl_stdar(arg1x_pad, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN '1'
     --synopsys translate_off
            | 'H'
     --synopsys translate_on
       =>
         RETURN fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_unsigned(
           fshl_stdar(arg1x, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit,  olen),
           fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen)
         );
         --synopsys translate_on
         RETURN result;
       END CASE;
     END IF;
   END;

   FUNCTION fshl_stdar(arg1: SIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
     CONSTANT arg1l: NATURAL := arg1'LENGTH - 1;
     ALIAS    arg1x: SIGNED(arg1l DOWNTO 0) IS arg1;
     CONSTANT arg2l: NATURAL := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE arg1x_pad: SIGNED(arg1l+1 DOWNTO 0);
     VARIABLE result: SIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others=>'0');
     arg1x_pad(arg1l+1) := sbit;
     arg1x_pad(arg1l downto 0) := arg1x;
     IF arg2l = 0 THEN
       RETURN fshr_stdar(arg1x_pad, UNSIGNED(arg2x), sbit, olen);
     -- ELSIF arg1l = 0 THEN
     --   RETURN fshl(sbit & arg1x, arg2x, sbit, olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
       =>
         RETURN fshl_stdar(arg1x_pad, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
       =>
         RETURN fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_signed(
           fshl_stdar(arg1x, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit,  olen),
           fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen)
         );
         --synopsys translate_on
         RETURN result;
       END CASE;
     END IF;
   END;

   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT arg2l: INTEGER := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE result: UNSIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others => '0');
     IF arg2l = 0 THEN
       RETURN fshl_stdar(arg1, UNSIGNED(arg2x), olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
        =>
         RETURN fshr_stdar(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
        =>
         RETURN fshl_stdar(arg1 & '0', '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_unsigned(
           fshr_stdar(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen),
           fshl_stdar(arg1 & '0', '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen)
         );
         --synopsys translate_on
	 return result;
       END CASE;
     END IF;
   END;

   FUNCTION fshr_stdar(arg1: SIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
     CONSTANT arg2l: INTEGER := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE result: SIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others => '0');
     IF arg2l = 0 THEN
       RETURN fshl_stdar(arg1, UNSIGNED(arg2x), olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
       =>
         RETURN fshr_stdar(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
       =>
         RETURN fshl_stdar(arg1 & '0', '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_signed(
           fshr_stdar(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen),
           fshl_stdar(arg1 & '0', '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen)
         );
         --synopsys translate_on
	 return result;
       END CASE;
     END IF;
   END;

   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshl_stdar(arg1, arg2, '0', olen); END;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshr_stdar(arg1, arg2, '0', olen); END;
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshl_stdar(arg1, arg2, '0', olen); END;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshr_stdar(arg1, arg2, '0', olen); END;

   FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN fshl_stdar(arg1, arg2, arg1(arg1'LEFT), olen); END;
   FUNCTION fshr_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN fshr_stdar(arg1, arg2, arg1(arg1'LEFT), olen); END;
   FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN fshl_stdar(arg1, arg2, arg1(arg1'LEFT), olen); END;
   FUNCTION fshr_stdar(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN fshr_stdar(arg1, arg2, arg1(arg1'LEFT), olen); END;


   FUNCTION fshl(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
     VARIABLE temp: UNSIGNED(len-1 DOWNTO 0);
     --SUBTYPE  sw_range IS NATURAL range 1 TO len;
     VARIABLE sw: NATURAL range 1 TO len;
     VARIABLE temp_idx : INTEGER; --2.1.6.3
   BEGIN
     sw := 1;
     result := (others => sbit);
     result(ilen-1 DOWNTO 0) := arg1;
     FOR i IN arg2'reverse_range LOOP
       temp := (others => '0');
       FOR i2 IN len-1-sw DOWNTO 0 LOOP
         --was:temp(i2+sw) := result(i2);
         temp_idx := add_nat(i2,sw);
         temp(temp_idx) := result(i2);
       END LOOP;
       result := UNSIGNED(mux_v(STD_LOGIC_VECTOR(concat_uns(result,temp)), arg2(i)));
       sw := minimum(mult_natural(sw,2), len);
     END LOOP;
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshr(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
     VARIABLE temp: UNSIGNED(len-1 DOWNTO 0);
     SUBTYPE  sw_range IS NATURAL range 1 TO len;
     VARIABLE sw: sw_range;
     VARIABLE result_idx : INTEGER; --2.1.6.3
   BEGIN
     sw := 1;
     result := (others => sbit);
     result(ilen-1 DOWNTO 0) := arg1;
     FOR i IN arg2'reverse_range LOOP
       temp := (others => sbit);
       FOR i2 IN len-1-sw DOWNTO 0 LOOP
         -- was: temp(i2) := result(i2+sw);
         result_idx := add_nat(i2,sw);
         temp(i2) := result(result_idx);
       END LOOP;
       result := UNSIGNED(mux_v(STD_LOGIC_VECTOR(concat_uns(result,temp)), arg2(i)));
       sw := minimum(mult_natural(sw,2), len);
     END LOOP;
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshl(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT arg1l: NATURAL := arg1'LENGTH - 1;
     ALIAS    arg1x: UNSIGNED(arg1l DOWNTO 0) IS arg1;
     CONSTANT arg2l: NATURAL := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE arg1x_pad: UNSIGNED(arg1l+1 DOWNTO 0);
     VARIABLE result: UNSIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others=>'0');
     arg1x_pad(arg1l+1) := sbit;
     arg1x_pad(arg1l downto 0) := arg1x;
     IF arg2l = 0 THEN
       RETURN fshr(arg1x_pad, UNSIGNED(arg2x), sbit, olen);
     -- ELSIF arg1l = 0 THEN
     --   RETURN fshl(sbit & arg1x, arg2x, sbit, olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
       =>
         RETURN fshl(arg1x_pad, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);

       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
       =>
         RETURN fshr(arg1x_pad(arg1l+1 DOWNTO 1), not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);

       WHEN others =>
         --synopsys translate_off
         result := resolve_unsigned(
           fshl(arg1x_pad, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit,  olen),
           fshr(arg1x_pad(arg1l+1 DOWNTO 1), not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen)
         );
         --synopsys translate_on
         RETURN result;
       END CASE;
     END IF;
   END;

   FUNCTION fshr(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT arg2l: INTEGER := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE result: UNSIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others => '0');
     IF arg2l = 0 THEN
       RETURN fshl(arg1, UNSIGNED(arg2x), olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
       =>
         RETURN fshr(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);

       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
       =>
         RETURN fshl(arg1 & '0', not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_unsigned(
           fshr(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen),
           fshl(arg1 & '0', not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen)
         );
         --synopsys translate_on
	 return result;
       END CASE;
     END IF;
   END;

   FUNCTION fshl(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshl(arg1, arg2, '0', olen); END;
   FUNCTION fshr(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshr(arg1, arg2, '0', olen); END;
   FUNCTION fshl(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshl(arg1, arg2, '0', olen); END;
   FUNCTION fshr(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshr(arg1, arg2, '0', olen); END;

   FUNCTION fshl(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN SIGNED(fshl(UNSIGNED(arg1), arg2, arg1(arg1'LEFT), olen)); END;
   FUNCTION fshr(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN SIGNED(fshr(UNSIGNED(arg1), arg2, arg1(arg1'LEFT), olen)); END;
   FUNCTION fshl(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN SIGNED(fshl(UNSIGNED(arg1), arg2, arg1(arg1'LEFT), olen)); END;
   FUNCTION fshr(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN SIGNED(fshr(UNSIGNED(arg1), arg2, arg1(arg1'LEFT), olen)); END;


   FUNCTION frot(arg1: STD_LOGIC_VECTOR; arg2: STD_LOGIC_VECTOR; signd2: BOOLEAN; sdir: INTEGER range -1 TO 1) RETURN STD_LOGIC_VECTOR IS
     CONSTANT len: INTEGER := arg1'LENGTH;
     VARIABLE result: STD_LOGIC_VECTOR(len-1 DOWNTO 0);
     VARIABLE temp: STD_LOGIC_VECTOR(len-1 DOWNTO 0);
     SUBTYPE sw_range IS NATURAL range 0 TO len-1;
     VARIABLE sw: sw_range;
     VARIABLE temp_idx : INTEGER; --2.1.6.3
   BEGIN
     result := (others=>'0');
     result := arg1;
     sw := sdir MOD len;
     FOR i IN arg2'reverse_range LOOP
       EXIT WHEN sw = 0;
       IF signd2 AND i = arg2'LEFT THEN 
         sw := sub_int(len,sw); 
       END IF;
       -- temp := result(len-sw-1 DOWNTO 0) & result(len-1 DOWNTO len-sw)
       FOR i2 IN len-1 DOWNTO 0 LOOP
         --was: temp((i2+sw) MOD len) := result(i2);
         temp_idx := add_nat(i2,sw) MOD len;
         temp(temp_idx) := result(i2);
       END LOOP;
       result := mux_v(STD_LOGIC_VECTOR(concat_vect(result,temp)), arg2(i));
       sw := mod_natural(mult_natural(sw,2), len);
     END LOOP;
     RETURN result;
   END frot;

   FUNCTION frol(arg1: STD_LOGIC_VECTOR; arg2: UNSIGNED) RETURN STD_LOGIC_VECTOR IS
     BEGIN RETURN frot(arg1, STD_LOGIC_VECTOR(arg2), FALSE, 1); END;
   FUNCTION fror(arg1: STD_LOGIC_VECTOR; arg2: UNSIGNED) RETURN STD_LOGIC_VECTOR IS
     BEGIN RETURN frot(arg1, STD_LOGIC_VECTOR(arg2), FALSE, -1); END;
   FUNCTION frol(arg1: STD_LOGIC_VECTOR; arg2: SIGNED  ) RETURN STD_LOGIC_VECTOR IS
     BEGIN RETURN frot(arg1, STD_LOGIC_VECTOR(arg2), TRUE, 1); END;
   FUNCTION fror(arg1: STD_LOGIC_VECTOR; arg2: SIGNED  ) RETURN STD_LOGIC_VECTOR IS
     BEGIN RETURN frot(arg1, STD_LOGIC_VECTOR(arg2), TRUE, -1); END;

-----------------------------------------------------------------
-- indexing functions: LSB always has index 0
-----------------------------------------------------------------

   FUNCTION readindex(vec: STD_LOGIC_VECTOR; index: INTEGER                 ) RETURN STD_LOGIC IS
     CONSTANT len : INTEGER := vec'LENGTH;
     ALIAS    vec0: STD_LOGIC_VECTOR(len-1 DOWNTO 0) IS vec;
   BEGIN
     IF index >= len OR index < 0 THEN
       RETURN 'X';
     END IF;
     RETURN vec0(index);
   END;

   FUNCTION readslice(vec: STD_LOGIC_VECTOR; index: INTEGER; width: POSITIVE) RETURN STD_LOGIC_VECTOR IS
     CONSTANT len : INTEGER := vec'LENGTH;
     CONSTANT indexPwidthM1 : INTEGER := index+width-1; --2.1.6.3
     ALIAS    vec0: STD_LOGIC_VECTOR(len-1 DOWNTO 0) IS vec;
     CONSTANT xxx : STD_LOGIC_VECTOR(width-1 DOWNTO 0) := (others => 'X');
   BEGIN
     IF index+width > len OR index < 0 THEN
       RETURN xxx;
     END IF;
     RETURN vec0(indexPwidthM1 DOWNTO index);
   END;

   FUNCTION writeindex(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC       ; index: INTEGER) RETURN STD_LOGIC_VECTOR IS
     CONSTANT len : INTEGER := vec'LENGTH;
     VARIABLE vec0: STD_LOGIC_VECTOR(len-1 DOWNTO 0);
     CONSTANT xxx : STD_LOGIC_VECTOR(len-1 DOWNTO 0) := (others => 'X');
   BEGIN
     vec0 := vec;
     IF index >= len OR index < 0 THEN
       RETURN xxx;
     END IF;
     vec0(index) := dinput;
     RETURN vec0;
   END;

   FUNCTION n_bits(p: NATURAL) RETURN POSITIVE IS
     VARIABLE n_b : POSITIVE;
     VARIABLE p_v : NATURAL;
   BEGIN
     p_v := p;
     FOR i IN 1 TO 32 LOOP
       p_v := div_natural(p_v,2);
       n_b := i;
       EXIT WHEN (p_v = 0);
     END LOOP;
     RETURN n_b;
   END;


--   FUNCTION writeslice(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC_VECTOR; index: INTEGER) RETURN STD_LOGIC_VECTOR IS
--
--     CONSTANT vlen: INTEGER := vec'LENGTH;
--     CONSTANT ilen: INTEGER := dinput'LENGTH;
--     CONSTANT max_shift: INTEGER := vlen-ilen;
--     CONSTANT ones: UNSIGNED(ilen-1 DOWNTO 0) := (others => '1');
--     CONSTANT xxx : STD_LOGIC_VECTOR(vlen-1 DOWNTO 0) := (others => 'X');
--     VARIABLE shift : UNSIGNED(n_bits(max_shift)-1 DOWNTO 0);
--     VARIABLE vec0: STD_LOGIC_VECTOR(vlen-1 DOWNTO 0);
--     VARIABLE inp: UNSIGNED(vlen-1 DOWNTO 0);
--     VARIABLE mask: UNSIGNED(vlen-1 DOWNTO 0);
--   BEGIN
--     inp := (others => '0');
--     mask := (others => '0');
--
--     IF index > max_shift OR index < 0 THEN
--       RETURN xxx;
--     END IF;
--
--     shift := CONV_UNSIGNED(index, shift'LENGTH);
--     inp(ilen-1 DOWNTO 0) := UNSIGNED(dinput);
--     mask(ilen-1 DOWNTO 0) := ones;
--     inp := fshl(inp, shift, vlen);
--     mask := fshl(mask, shift, vlen);
--     vec0 := (vec and (not STD_LOGIC_VECTOR(mask))) or STD_LOGIC_VECTOR(inp);
--     RETURN vec0;
--   END;

   FUNCTION writeslice(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC_VECTOR; enable: STD_LOGIC_VECTOR; byte_width: INTEGER;  index: INTEGER) RETURN STD_LOGIC_VECTOR IS

     type enable_matrix is array (0 to enable'LENGTH-1 ) of std_logic_vector(byte_width-1 downto 0);
     CONSTANT vlen: INTEGER := vec'LENGTH;
     CONSTANT ilen: INTEGER := dinput'LENGTH;
     CONSTANT max_shift: INTEGER := vlen-ilen;
     CONSTANT ones: UNSIGNED(ilen-1 DOWNTO 0) := (others => '1');
     CONSTANT xxx : STD_LOGIC_VECTOR(vlen-1 DOWNTO 0) := (others => 'X');
     VARIABLE shift : UNSIGNED(n_bits(max_shift)-1 DOWNTO 0);
     VARIABLE vec0: STD_LOGIC_VECTOR(vlen-1 DOWNTO 0);
     VARIABLE inp: UNSIGNED(vlen-1 DOWNTO 0);
     VARIABLE mask: UNSIGNED(vlen-1 DOWNTO 0);
     VARIABLE mask2: UNSIGNED(vlen-1 DOWNTO 0);
     VARIABLE enables: enable_matrix;
     VARIABLE cat_enables: STD_LOGIC_VECTOR(ilen-1 DOWNTO 0 );
     VARIABLE lsbi : INTEGER;
     VARIABLE msbi : INTEGER;

   BEGIN
     cat_enables := (others => '0');
     lsbi := 0;
     msbi := byte_width-1;
     inp := (others => '0');
     mask := (others => '0');

     IF index > max_shift OR index < 0 THEN
       RETURN xxx;
     END IF;

     --initialize enables
     for i in 0 TO (enable'LENGTH-1) loop
       enables(i)  := (others => enable(i));
       cat_enables(msbi downto lsbi) := enables(i) ;
       lsbi := msbi+1;
       msbi := msbi+byte_width;
     end loop;


     shift := CONV_UNSIGNED(index, shift'LENGTH);
     inp(ilen-1 DOWNTO 0) := UNSIGNED(dinput);
     mask(ilen-1 DOWNTO 0) := UNSIGNED((STD_LOGIC_VECTOR(ones) AND cat_enables));
     inp := fshl(inp, shift, vlen);
     mask := fshl(mask, shift, vlen);
     vec0 := (vec and (not STD_LOGIC_VECTOR(mask))) or STD_LOGIC_VECTOR(inp);
     RETURN vec0;
   END;


   FUNCTION ceil_log2(size : NATURAL) return NATURAL is
     VARIABLE cnt : NATURAL;
     VARIABLE res : NATURAL;
   begin
     cnt := 1;
     res := 0;
     while (cnt < size) loop
       res := res + 1;
       cnt := 2 * cnt;
     end loop;
     return res;
   END;
   
   FUNCTION bits(size : NATURAL) return NATURAL is
   begin
     return ceil_log2(size);
   END;

   PROCEDURE csa(a, b, c: IN INTEGER; s, cout: OUT STD_LOGIC_VECTOR) IS
   BEGIN
     s    := conv_std_logic_vector(a, s'LENGTH) xor conv_std_logic_vector(b, s'LENGTH) xor conv_std_logic_vector(c, s'LENGTH);
     cout := ( (conv_std_logic_vector(a, cout'LENGTH) and conv_std_logic_vector(b, cout'LENGTH)) or (conv_std_logic_vector(a, cout'LENGTH) and conv_std_logic_vector(c, cout'LENGTH)) or (conv_std_logic_vector(b, cout'LENGTH) and conv_std_logic_vector(c, cout'LENGTH)) );
   END PROCEDURE csa;

   PROCEDURE csha(a, b: IN INTEGER; s, cout: OUT STD_LOGIC_VECTOR) IS
   BEGIN
     s    := conv_std_logic_vector(a, s'LENGTH) xor conv_std_logic_vector(b, s'LENGTH);
     cout := (conv_std_logic_vector(a, cout'LENGTH) and conv_std_logic_vector(b, cout'LENGTH));
   END PROCEDURE csha;

END funcs;

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_comps.vhd 
LIBRARY ieee;

USE ieee.std_logic_1164.all;

PACKAGE mgc_comps IS
 
FUNCTION ifeqsel(arg1, arg2, seleq, selne : INTEGER) RETURN INTEGER;
FUNCTION ceil_log2(size : NATURAL) return NATURAL;
 

COMPONENT mgc_not
  GENERIC (
    width  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    z: out std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_and
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_nand
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_or
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_nor
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_xor
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_xnor
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mux
  GENERIC (
    width  :  NATURAL;
    ctrlw  :  NATURAL;
    p2ctrlw : NATURAL := 0
  );
  PORT (
    a: in  std_logic_vector(width*(2**ctrlw) - 1 DOWNTO 0);
    c: in  std_logic_vector(ctrlw            - 1 DOWNTO 0);
    z: out std_logic_vector(width            - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mux1hot
  GENERIC (
    width  : NATURAL;
    ctrlw  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ctrlw - 1 DOWNTO 0);
    c: in  std_logic_vector(ctrlw       - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_reg_pos
  GENERIC (
    width  : NATURAL;
    has_a_rst : NATURAL;  -- 0 to 1
    a_rst_on  : NATURAL;  -- 0 to 1
    has_s_rst : NATURAL;  -- 0 to 1
    s_rst_on  : NATURAL;  -- 0 to 1
    has_enable : NATURAL; -- 0 to 1
    enable_on  : NATURAL  -- 0 to 1
  );
  PORT (
    clk: in  std_logic;
    d  : in  std_logic_vector(width-1 DOWNTO 0);
    z  : out std_logic_vector(width-1 DOWNTO 0);
    sync_rst_val : in std_logic_vector(width-1 DOWNTO 0);
    sync_rst : in std_logic;
    async_rst_val : in std_logic_vector(width-1 DOWNTO 0);
    async_rst : in std_logic;
    en : in std_logic
  );
END COMPONENT;

COMPONENT mgc_reg_neg
  GENERIC (
    width  : NATURAL;
    has_a_rst : NATURAL;  -- 0 to 1
    a_rst_on  : NATURAL;  -- 0 to 1
    has_s_rst : NATURAL;  -- 0 to 1
    s_rst_on  : NATURAL;   -- 0 to 1
    has_enable : NATURAL; -- 0 to 1
    enable_on  : NATURAL -- 0 to 1
  );
  PORT (
    clk: in  std_logic;
    d  : in  std_logic_vector(width-1 DOWNTO 0);
    z  : out std_logic_vector(width-1 DOWNTO 0);
    sync_rst_val : in std_logic_vector(width-1 DOWNTO 0);
    sync_rst : in std_logic;
    async_rst_val : in std_logic_vector(width-1 DOWNTO 0);
    async_rst : in std_logic;
    en : in std_logic
  );
END COMPONENT;

COMPONENT mgc_generic_reg
  GENERIC(
   width: natural := 8;
   ph_clk: integer range 0 to 1 := 1; -- clock polarity, 1=rising_edge
   ph_en: integer range 0 to 1 := 1;
   ph_a_rst: integer range 0 to 1 := 1;   --  0 to 1 IGNORED
   ph_s_rst: integer range 0 to 1 := 1;   --  0 to 1 IGNORED
   a_rst_used: integer range 0 to 1 := 1;
   s_rst_used: integer range 0 to 1 := 0;
   en_used: integer range 0 to 1 := 1
  );
  PORT(
   d: std_logic_vector(width-1 downto 0);
   clk: in std_logic;
   en: in std_logic;
   a_rst: in std_logic;
   s_rst: in std_logic;
   q: out std_logic_vector(width-1 downto 0)
  );
END COMPONENT;

COMPONENT mgc_equal
  GENERIC (
    width  : NATURAL
  );
  PORT (
    a : in  std_logic_vector(width-1 DOWNTO 0);
    b : in  std_logic_vector(width-1 DOWNTO 0);
    eq: out std_logic;
    ne: out std_logic
  );
END COMPONENT;

COMPONENT mgc_shift_l
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_r
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_bl
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_br
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_rot
  GENERIC (
    width  : NATURAL;
    width_s: NATURAL;
    signd_s: NATURAL;      -- 0:unsigned 1:signed
    sleft  : NATURAL;      -- 0:right 1:left;
    log2w  : NATURAL := 0; -- LOG2(width)
    l2wp2  : NATURAL := 0  --2**LOG2(width)
  );
  PORT (
    a : in  std_logic_vector(width  -1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width  -1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_add
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_sub
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_add_ci
  GENERIC (
    width_a : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width_a, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width_a, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width_a,width_b)-1 DOWNTO 0);
    c: in  std_logic_vector(0 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width_a,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_addc
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    c: in  std_logic_vector(0 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_add3
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_c : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_c : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    c: in  std_logic_vector(ifeqsel(width_c,0,width,width_c)-1 DOWNTO 0);
    d: in  std_logic_vector(0 DOWNTO 0);
    e: in  std_logic_vector(0 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_add_pipe
  GENERIC (
     width_a : natural := 16;
     signd_a : integer range 0 to 1 := 0;
     width_b : natural := 3;
     signd_b : integer range 0 to 1 := 0;
     width_z : natural := 18;
     ph_clk : integer range 0 to 1 := 1;
     ph_en : integer range 0 to 1 := 1;
     ph_a_rst : integer range 0 to 1 := 1;
     ph_s_rst : integer range 0 to 1 := 1;
     n_outreg : natural := 2;
     stages : natural := 2; -- Default value is minimum required value
     a_rst_used: integer range 0 to 1 := 1;
     s_rst_used: integer range 0 to 1 := 0;
     en_used: integer range 0 to 1 := 1
     );
  PORT(
     a: in std_logic_vector(width_a-1 downto 0);
     b: in std_logic_vector(width_b-1 downto 0);
     clk: in std_logic;
     en: in std_logic;
     a_rst: in std_logic;
     s_rst: in std_logic;
     z: out std_logic_vector(width_z-1 downto 0)
     );
END COMPONENT;

COMPONENT mgc_sub_pipe
  GENERIC (
     width_a : natural := 16;
     signd_a : integer range 0 to 1 := 0;
     width_b : natural := 3;
     signd_b : integer range 0 to 1 := 0;
     width_z : natural := 18;
     ph_clk : integer range 0 to 1 := 1;
     ph_en : integer range 0 to 1 := 1;
     ph_a_rst : integer range 0 to 1 := 1;
     ph_s_rst : integer range 0 to 1 := 1;
     n_outreg : natural := 2;
     stages : natural := 2; -- Default value is minimum required value
     a_rst_used: integer range 0 to 1 := 1;
     s_rst_used: integer range 0 to 1 := 0;
     en_used: integer range 0 to 1 := 1
     );
  PORT(
     a: in std_logic_vector(width_a-1 downto 0);
     b: in std_logic_vector(width_b-1 downto 0);
     clk: in std_logic;
     en: in std_logic;
     a_rst: in std_logic;
     s_rst: in std_logic;
     z: out std_logic_vector(width_z-1 downto 0)
     );
END COMPONENT;

COMPONENT mgc_addc_pipe
  GENERIC (
     width_a : natural := 16;
     signd_a : integer range 0 to 1 := 0;
     width_b : natural := 3;
     signd_b : integer range 0 to 1 := 0;
     width_z : natural := 18;
     ph_clk : integer range 0 to 1 := 1;
     ph_en : integer range 0 to 1 := 1;
     ph_a_rst : integer range 0 to 1 := 1;
     ph_s_rst : integer range 0 to 1 := 1;
     n_outreg : natural := 2;
     stages : natural := 2; -- Default value is minimum required value
     a_rst_used: integer range 0 to 1 := 1;
     s_rst_used: integer range 0 to 1 := 0;
     en_used: integer range 0 to 1 := 1
     );
  PORT(
     a: in std_logic_vector(width_a-1 downto 0);
     b: in std_logic_vector(width_b-1 downto 0);
     c: in std_logic_vector(0 downto 0);
     clk: in std_logic;
     en: in std_logic;
     a_rst: in std_logic;
     s_rst: in std_logic;
     z: out std_logic_vector(width_z-1 downto 0)
     );
END COMPONENT;

COMPONENT mgc_addsub
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    add: in  std_logic;
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_accu
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps-1 DOWNTO 0);
    z: out std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_abs
  GENERIC (
    width  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    z: out std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_z : NATURAL    -- <= width_a + width_b
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul_fast
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_z : NATURAL    -- <= width_a + width_b
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul_pipe
  GENERIC (
    width_a       : NATURAL;
    signd_a       : NATURAL;
    width_b       : NATURAL;
    signd_b       : NATURAL;
    width_z       : NATURAL; -- <= width_a + width_b
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 

  );
  PORT (
    a     : in  std_logic_vector(width_a-1 DOWNTO 0);
    b     : in  std_logic_vector(width_b-1 DOWNTO 0);
    clk   : in  std_logic;
    en    : in  std_logic;
    a_rst : in  std_logic;
    s_rst : in  std_logic;
    z     : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul2add1
  GENERIC (
    gentype : NATURAL;
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_b2 : NATURAL;
    signd_b2 : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_d2 : NATURAL;
    signd_d2 : NATURAL;
    width_e : NATURAL;
    signd_e : NATURAL;
    width_z : NATURAL;   -- <= max(width_a + width_b, width_c + width_d)+1
    isadd   : NATURAL;
    add_b2  : NATURAL;
    add_d2  : NATURAL
  );
  PORT (
    a   : in  std_logic_vector(width_a-1 DOWNTO 0);
    b   : in  std_logic_vector(width_b-1 DOWNTO 0);
    b2  : in  std_logic_vector(width_b2-1 DOWNTO 0);
    c   : in  std_logic_vector(width_c-1 DOWNTO 0);
    d   : in  std_logic_vector(width_d-1 DOWNTO 0);
    d2  : in  std_logic_vector(width_d2-1 DOWNTO 0);
    cst : in  std_logic_vector(width_e-1 DOWNTO 0);
    z   : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul2add1_pipe
  GENERIC (
    gentype : NATURAL;
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_b2 : NATURAL;
    signd_b2 : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_d2 : NATURAL;
    signd_d2 : NATURAL;
    width_e : NATURAL;
    signd_e : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c + width_d)+1
    isadd   : NATURAL;
    add_b2   : NATURAL;
    add_d2   : NATURAL;
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 
  );
  PORT (
    a     : in  std_logic_vector(width_a-1 DOWNTO 0);
    b     : in  std_logic_vector(width_b-1 DOWNTO 0);
    b2     : in  std_logic_vector(width_b2-1 DOWNTO 0);
    c     : in  std_logic_vector(width_c-1 DOWNTO 0);
    d     : in  std_logic_vector(width_d-1 DOWNTO 0);
    d2     : in  std_logic_vector(width_d2-1 DOWNTO 0);
    cst   : in  std_logic_vector(width_e-1 DOWNTO 0);
    clk   : in  std_logic;
    en    : in  std_logic;
    a_rst : in  std_logic;
    s_rst : in  std_logic;
    z     : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_muladd1
  -- operation is z = a * (b + d) + c + cst
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_cst : NATURAL;
    signd_cst : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c, width_cst)+1
    add_axb : NATURAL;
    add_c   : NATURAL;
    add_d   : NATURAL
  );
  PORT (
    a:   in  std_logic_vector(width_a-1 DOWNTO 0);
    b:   in  std_logic_vector(width_b-1 DOWNTO 0);
    c:   in  std_logic_vector(width_c-1 DOWNTO 0);
    cst: in  std_logic_vector(width_cst-1 DOWNTO 0);
    d:   in  std_logic_vector(width_d-1 DOWNTO 0);
    z:   out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_muladd1_pipe
  -- operation is z = a * (b + d) + c + cst
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_cst : NATURAL;
    signd_cst : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c, width_cst)+1
    add_axb : NATURAL;
    add_c   : NATURAL;
    add_d   : NATURAL;
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 
  );
  PORT (
    a     : in  std_logic_vector(width_a-1 DOWNTO 0);
    b     : in  std_logic_vector(width_b-1 DOWNTO 0);
    c     : in  std_logic_vector(width_c-1 DOWNTO 0);
    cst   : in  std_logic_vector(width_cst-1 DOWNTO 0);
    d     : in  std_logic_vector(width_d-1 DOWNTO 0);
    clk   : in  std_logic;
    en    : in  std_logic;
    a_rst : in  std_logic;
    s_rst : in  std_logic;
    z     : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mulacc_pipe
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c)+1
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 
  );
  PORT (
    a         : in  std_logic_vector(width_a-1 DOWNTO 0);
    b         : in  std_logic_vector(width_b-1 DOWNTO 0);
    c         : in  std_logic_vector(width_c-1 DOWNTO 0);
    load      : in  std_logic;
    datavalid : in  std_logic;
    clk       : in  std_logic;
    en        : in  std_logic;
    a_rst     : in  std_logic;
    s_rst     : in  std_logic;
    z         : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul2acc_pipe
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_e : NATURAL;
    signd_e : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c)+1
    add_cxd : NATURAL;
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 
  );
  PORT (
    a         : in  std_logic_vector(width_a-1 DOWNTO 0);
    b         : in  std_logic_vector(width_b-1 DOWNTO 0);
    c         : in  std_logic_vector(width_c-1 DOWNTO 0);
    d         : in  std_logic_vector(width_d-1 DOWNTO 0);
    e         : in  std_logic_vector(width_e-1 DOWNTO 0);
    load      : in  std_logic;
    datavalid : in  std_logic;
    clk       : in  std_logic;
    en        : in  std_logic;
    a_rst     : in  std_logic;
    s_rst     : in  std_logic;
    z         : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_div
  GENERIC (
    width_a : NATURAL;
    width_b : NATURAL;
    signd   : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_a-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mod
  GENERIC (
    width_a : NATURAL;
    width_b : NATURAL;
    signd   : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_b-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_rem
  GENERIC (
    width_a : NATURAL;
    width_b : NATURAL;
    signd   : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_b-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_csa
  GENERIC (
     width : NATURAL
  );
  PORT (
     a: in std_logic_vector(width-1 downto 0);
     b: in std_logic_vector(width-1 downto 0);
     c: in std_logic_vector(width-1 downto 0);
     s: out std_logic_vector(width-1 downto 0);
     cout: out std_logic_vector(width-1 downto 0)
  );
END COMPONENT;

COMPONENT mgc_csha
  GENERIC (
     width : NATURAL
  );
  PORT (
     a: in std_logic_vector(width-1 downto 0);
     b: in std_logic_vector(width-1 downto 0);
     s: out std_logic_vector(width-1 downto 0);
     cout: out std_logic_vector(width-1 downto 0)
  );
END COMPONENT;

COMPONENT mgc_rom
    GENERIC (
      rom_id : natural := 1;
      size : natural := 33;
      width : natural := 32
      );
    PORT (
      data_in : std_logic_vector((size*width)-1 downto 0);
      addr : std_logic_vector(ceil_log2(size)-1 downto 0);
      data_out : out std_logic_vector(width-1 downto 0)
    );
END COMPONENT;

END mgc_comps;

PACKAGE BODY mgc_comps IS
 
   FUNCTION ceil_log2(size : NATURAL) return NATURAL is
     VARIABLE cnt : NATURAL;
     VARIABLE res : NATURAL;
   begin
     cnt := 1;
     res := 0;
     while (cnt < size) loop
       res := res + 1;
       cnt := 2 * cnt;
     end loop;
     return res;
   END;

   FUNCTION ifeqsel(arg1, arg2, seleq, selne : INTEGER) RETURN INTEGER IS
   BEGIN
     IF(arg1 = arg2) THEN
       RETURN(seleq) ;
     ELSE
       RETURN(selne) ;
     END IF;
   END;
 
END mgc_comps;

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_rem_beh.vhd 

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY mgc_rem IS
  GENERIC (
    width_a : NATURAL;
    width_b : NATURAL;
    signd   : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_b-1 DOWNTO 0)
  );
END mgc_rem;

LIBRARY ieee;

USE ieee.std_logic_arith.all;

USE work.funcs.all;

ARCHITECTURE beh OF mgc_rem IS
BEGIN
  z <= std_logic_vector(unsigned(a) rem unsigned(b)) WHEN signd = 0 ELSE
       std_logic_vector(  signed(a) rem   signed(b));
END beh;

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_div_beh.vhd 

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY mgc_div IS
  GENERIC (
    width_a : NATURAL;
    width_b : NATURAL;
    signd   : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_a-1 DOWNTO 0)
  );
END mgc_div;

LIBRARY ieee;

USE ieee.std_logic_arith.all;

USE work.funcs.all;

ARCHITECTURE beh OF mgc_div IS
BEGIN
  z <= std_logic_vector(unsigned(a) / unsigned(b)) WHEN signd = 0 ELSE
       std_logic_vector(  signed(a) /   signed(b));
END beh;

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_shift_comps_v5.vhd 
LIBRARY ieee;

USE ieee.std_logic_1164.all;

PACKAGE mgc_shift_comps_v5 IS

COMPONENT mgc_shift_l_v5
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_r_v5
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_bl_v5
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_br_v5
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

END mgc_shift_comps_v5;

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_shift_l_beh_v5.vhd 
LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY mgc_shift_l_v5 IS
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END mgc_shift_l_v5;

LIBRARY ieee;

USE ieee.std_logic_arith.all;

ARCHITECTURE beh OF mgc_shift_l_v5 IS

  FUNCTION maximum (arg1,arg2: INTEGER) RETURN INTEGER IS
  BEGIN
    IF(arg1 > arg2) THEN
      RETURN(arg1) ;
    ELSE
      RETURN(arg2) ;
    END IF;
  END;

  FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
    CONSTANT ilen: INTEGER := arg1'LENGTH;
    CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
    CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
    CONSTANT len: INTEGER := maximum(ilen, olen);
    VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
  BEGIN
    result := (others => sbit);
    result(ilenub DOWNTO 0) := arg1;
    result := shl(result, arg2);
    RETURN result(olenM1 DOWNTO 0);
  END;

  FUNCTION fshl_stdar(arg1: SIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
    CONSTANT ilen: INTEGER := arg1'LENGTH;
    CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
    CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
    CONSTANT len: INTEGER := maximum(ilen, olen);
    VARIABLE result: SIGNED(len-1 DOWNTO 0);
  BEGIN
    result := (others => sbit);
    result(ilenub DOWNTO 0) := arg1;
    result := shl(SIGNED(result), arg2);
    RETURN result(olenM1 DOWNTO 0);
  END;

  FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE)
  RETURN UNSIGNED IS
  BEGIN
    RETURN fshl_stdar(arg1, arg2, '0', olen);
  END;

  FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE)
  RETURN SIGNED IS
  BEGIN
    RETURN fshl_stdar(arg1, arg2, arg1(arg1'LEFT), olen);
  END;

BEGIN
UNSGNED:  IF signd_a = 0 GENERATE
    z <= std_logic_vector(fshl_stdar(unsigned(a), unsigned(s), width_z));
  END GENERATE;
SGNED:  IF signd_a /= 0 GENERATE
    z <= std_logic_vector(fshl_stdar(  signed(a), unsigned(s), width_z));
  END GENERATE;
END beh;

--------> ./rtl.vhdl 
-- ----------------------------------------------------------------------
--  HLS HDL:        VHDL Netlister
--  HLS Version:    10.5c/896140 Production Release
--  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
-- 
--  Generated by:   yl7897@newnano.poly.edu
--  Generated date: Thu Jul  1 13:31:47 2021
-- ----------------------------------------------------------------------

-- 
-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_19_8_64_256_256_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_19_8_64_256_256_64_1_gen
    IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_19_8_64_256_256_64_1_gen;

ARCHITECTURE v44 OF inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_19_8_64_256_256_64_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v44;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_18_8_64_256_256_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_18_8_64_256_256_64_1_gen
    IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_18_8_64_256_256_64_1_gen;

ARCHITECTURE v44 OF inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_18_8_64_256_256_64_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v44;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_17_8_64_256_256_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_17_8_64_256_256_64_1_gen
    IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_17_8_64_256_256_64_1_gen;

ARCHITECTURE v44 OF inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_17_8_64_256_256_64_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v44;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_16_8_64_256_256_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_16_8_64_256_256_64_1_gen
    IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_16_8_64_256_256_64_1_gen;

ARCHITECTURE v44 OF inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_16_8_64_256_256_64_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v44;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_15_8_64_256_256_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_15_8_64_256_256_64_1_gen
    IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_15_8_64_256_256_64_1_gen;

ARCHITECTURE v44 OF inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_15_8_64_256_256_64_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v44;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_14_8_64_256_256_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_14_8_64_256_256_64_1_gen
    IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_14_8_64_256_256_64_1_gen;

ARCHITECTURE v44 OF inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_14_8_64_256_256_64_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v44;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_13_8_64_256_256_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_13_8_64_256_256_64_1_gen
    IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_13_8_64_256_256_64_1_gen;

ARCHITECTURE v44 OF inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_13_8_64_256_256_64_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v44;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_12_8_64_256_256_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_12_8_64_256_256_64_1_gen
    IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_12_8_64_256_256_64_1_gen;

ARCHITECTURE v44 OF inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_12_8_64_256_256_64_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v44;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_11_8_64_256_256_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_11_8_64_256_256_64_1_gen
    IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_11_8_64_256_256_64_1_gen;

ARCHITECTURE v44 OF inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_11_8_64_256_256_64_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v44;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_10_8_64_256_256_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_10_8_64_256_256_64_1_gen
    IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_10_8_64_256_256_64_1_gen;

ARCHITECTURE v44 OF inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_10_8_64_256_256_64_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v44;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_9_8_64_256_256_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_9_8_64_256_256_64_1_gen
    IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_9_8_64_256_256_64_1_gen;

ARCHITECTURE v44 OF inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_9_8_64_256_256_64_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v44;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_8_8_64_256_256_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_8_8_64_256_256_64_1_gen
    IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_8_8_64_256_256_64_1_gen;

ARCHITECTURE v44 OF inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_8_8_64_256_256_64_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v44;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_7_8_64_256_256_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_7_8_64_256_256_64_1_gen
    IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_7_8_64_256_256_64_1_gen;

ARCHITECTURE v44 OF inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_7_8_64_256_256_64_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v44;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_6_8_64_256_256_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_6_8_64_256_256_64_1_gen
    IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_6_8_64_256_256_64_1_gen;

ARCHITECTURE v44 OF inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_6_8_64_256_256_64_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v44;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_5_8_64_256_256_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_5_8_64_256_256_64_1_gen
    IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_5_8_64_256_256_64_1_gen;

ARCHITECTURE v44 OF inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_5_8_64_256_256_64_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v44;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_4_8_64_256_256_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_4_8_64_256_256_64_1_gen
    IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_4_8_64_256_256_64_1_gen;

ARCHITECTURE v44 OF inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_4_8_64_256_256_64_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v44;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT_core_core_fsm
--  FSM Module
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT_core_core_fsm IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    fsm_output : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
    STAGE_LOOP_C_8_tr0 : IN STD_LOGIC;
    modExp_while_C_38_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_1_tr0 : IN STD_LOGIC;
    COMP_LOOP_1_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_64_tr0 : IN STD_LOGIC;
    COMP_LOOP_2_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_128_tr0 : IN STD_LOGIC;
    COMP_LOOP_3_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_192_tr0 : IN STD_LOGIC;
    COMP_LOOP_4_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_256_tr0 : IN STD_LOGIC;
    COMP_LOOP_5_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_320_tr0 : IN STD_LOGIC;
    COMP_LOOP_6_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_384_tr0 : IN STD_LOGIC;
    COMP_LOOP_7_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_448_tr0 : IN STD_LOGIC;
    COMP_LOOP_8_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_512_tr0 : IN STD_LOGIC;
    COMP_LOOP_9_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_576_tr0 : IN STD_LOGIC;
    COMP_LOOP_10_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_640_tr0 : IN STD_LOGIC;
    COMP_LOOP_11_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_704_tr0 : IN STD_LOGIC;
    COMP_LOOP_12_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_768_tr0 : IN STD_LOGIC;
    COMP_LOOP_13_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_832_tr0 : IN STD_LOGIC;
    COMP_LOOP_14_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_896_tr0 : IN STD_LOGIC;
    COMP_LOOP_15_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_960_tr0 : IN STD_LOGIC;
    COMP_LOOP_16_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_1024_tr0 : IN STD_LOGIC;
    VEC_LOOP_C_0_tr0 : IN STD_LOGIC;
    STAGE_LOOP_C_9_tr0 : IN STD_LOGIC
  );
END inPlaceNTT_DIT_core_core_fsm;

ARCHITECTURE v44 OF inPlaceNTT_DIT_core_core_fsm IS
  -- Default Constants

  -- FSM State Type Declaration for inPlaceNTT_DIT_core_core_fsm_1
  TYPE inPlaceNTT_DIT_core_core_fsm_1_ST IS (main_C_0, STAGE_LOOP_C_0, STAGE_LOOP_C_1,
      STAGE_LOOP_C_2, STAGE_LOOP_C_3, STAGE_LOOP_C_4, STAGE_LOOP_C_5, STAGE_LOOP_C_6,
      STAGE_LOOP_C_7, STAGE_LOOP_C_8, modExp_while_C_0, modExp_while_C_1, modExp_while_C_2,
      modExp_while_C_3, modExp_while_C_4, modExp_while_C_5, modExp_while_C_6, modExp_while_C_7,
      modExp_while_C_8, modExp_while_C_9, modExp_while_C_10, modExp_while_C_11, modExp_while_C_12,
      modExp_while_C_13, modExp_while_C_14, modExp_while_C_15, modExp_while_C_16,
      modExp_while_C_17, modExp_while_C_18, modExp_while_C_19, modExp_while_C_20,
      modExp_while_C_21, modExp_while_C_22, modExp_while_C_23, modExp_while_C_24,
      modExp_while_C_25, modExp_while_C_26, modExp_while_C_27, modExp_while_C_28,
      modExp_while_C_29, modExp_while_C_30, modExp_while_C_31, modExp_while_C_32,
      modExp_while_C_33, modExp_while_C_34, modExp_while_C_35, modExp_while_C_36,
      modExp_while_C_37, modExp_while_C_38, COMP_LOOP_C_0, COMP_LOOP_C_1, COMP_LOOP_1_modExp_1_while_C_0,
      COMP_LOOP_1_modExp_1_while_C_1, COMP_LOOP_1_modExp_1_while_C_2, COMP_LOOP_1_modExp_1_while_C_3,
      COMP_LOOP_1_modExp_1_while_C_4, COMP_LOOP_1_modExp_1_while_C_5, COMP_LOOP_1_modExp_1_while_C_6,
      COMP_LOOP_1_modExp_1_while_C_7, COMP_LOOP_1_modExp_1_while_C_8, COMP_LOOP_1_modExp_1_while_C_9,
      COMP_LOOP_1_modExp_1_while_C_10, COMP_LOOP_1_modExp_1_while_C_11, COMP_LOOP_1_modExp_1_while_C_12,
      COMP_LOOP_1_modExp_1_while_C_13, COMP_LOOP_1_modExp_1_while_C_14, COMP_LOOP_1_modExp_1_while_C_15,
      COMP_LOOP_1_modExp_1_while_C_16, COMP_LOOP_1_modExp_1_while_C_17, COMP_LOOP_1_modExp_1_while_C_18,
      COMP_LOOP_1_modExp_1_while_C_19, COMP_LOOP_1_modExp_1_while_C_20, COMP_LOOP_1_modExp_1_while_C_21,
      COMP_LOOP_1_modExp_1_while_C_22, COMP_LOOP_1_modExp_1_while_C_23, COMP_LOOP_1_modExp_1_while_C_24,
      COMP_LOOP_1_modExp_1_while_C_25, COMP_LOOP_1_modExp_1_while_C_26, COMP_LOOP_1_modExp_1_while_C_27,
      COMP_LOOP_1_modExp_1_while_C_28, COMP_LOOP_1_modExp_1_while_C_29, COMP_LOOP_1_modExp_1_while_C_30,
      COMP_LOOP_1_modExp_1_while_C_31, COMP_LOOP_1_modExp_1_while_C_32, COMP_LOOP_1_modExp_1_while_C_33,
      COMP_LOOP_1_modExp_1_while_C_34, COMP_LOOP_1_modExp_1_while_C_35, COMP_LOOP_1_modExp_1_while_C_36,
      COMP_LOOP_1_modExp_1_while_C_37, COMP_LOOP_1_modExp_1_while_C_38, COMP_LOOP_C_2,
      COMP_LOOP_C_3, COMP_LOOP_C_4, COMP_LOOP_C_5, COMP_LOOP_C_6, COMP_LOOP_C_7,
      COMP_LOOP_C_8, COMP_LOOP_C_9, COMP_LOOP_C_10, COMP_LOOP_C_11, COMP_LOOP_C_12,
      COMP_LOOP_C_13, COMP_LOOP_C_14, COMP_LOOP_C_15, COMP_LOOP_C_16, COMP_LOOP_C_17,
      COMP_LOOP_C_18, COMP_LOOP_C_19, COMP_LOOP_C_20, COMP_LOOP_C_21, COMP_LOOP_C_22,
      COMP_LOOP_C_23, COMP_LOOP_C_24, COMP_LOOP_C_25, COMP_LOOP_C_26, COMP_LOOP_C_27,
      COMP_LOOP_C_28, COMP_LOOP_C_29, COMP_LOOP_C_30, COMP_LOOP_C_31, COMP_LOOP_C_32,
      COMP_LOOP_C_33, COMP_LOOP_C_34, COMP_LOOP_C_35, COMP_LOOP_C_36, COMP_LOOP_C_37,
      COMP_LOOP_C_38, COMP_LOOP_C_39, COMP_LOOP_C_40, COMP_LOOP_C_41, COMP_LOOP_C_42,
      COMP_LOOP_C_43, COMP_LOOP_C_44, COMP_LOOP_C_45, COMP_LOOP_C_46, COMP_LOOP_C_47,
      COMP_LOOP_C_48, COMP_LOOP_C_49, COMP_LOOP_C_50, COMP_LOOP_C_51, COMP_LOOP_C_52,
      COMP_LOOP_C_53, COMP_LOOP_C_54, COMP_LOOP_C_55, COMP_LOOP_C_56, COMP_LOOP_C_57,
      COMP_LOOP_C_58, COMP_LOOP_C_59, COMP_LOOP_C_60, COMP_LOOP_C_61, COMP_LOOP_C_62,
      COMP_LOOP_C_63, COMP_LOOP_C_64, COMP_LOOP_C_65, COMP_LOOP_2_modExp_1_while_C_0,
      COMP_LOOP_2_modExp_1_while_C_1, COMP_LOOP_2_modExp_1_while_C_2, COMP_LOOP_2_modExp_1_while_C_3,
      COMP_LOOP_2_modExp_1_while_C_4, COMP_LOOP_2_modExp_1_while_C_5, COMP_LOOP_2_modExp_1_while_C_6,
      COMP_LOOP_2_modExp_1_while_C_7, COMP_LOOP_2_modExp_1_while_C_8, COMP_LOOP_2_modExp_1_while_C_9,
      COMP_LOOP_2_modExp_1_while_C_10, COMP_LOOP_2_modExp_1_while_C_11, COMP_LOOP_2_modExp_1_while_C_12,
      COMP_LOOP_2_modExp_1_while_C_13, COMP_LOOP_2_modExp_1_while_C_14, COMP_LOOP_2_modExp_1_while_C_15,
      COMP_LOOP_2_modExp_1_while_C_16, COMP_LOOP_2_modExp_1_while_C_17, COMP_LOOP_2_modExp_1_while_C_18,
      COMP_LOOP_2_modExp_1_while_C_19, COMP_LOOP_2_modExp_1_while_C_20, COMP_LOOP_2_modExp_1_while_C_21,
      COMP_LOOP_2_modExp_1_while_C_22, COMP_LOOP_2_modExp_1_while_C_23, COMP_LOOP_2_modExp_1_while_C_24,
      COMP_LOOP_2_modExp_1_while_C_25, COMP_LOOP_2_modExp_1_while_C_26, COMP_LOOP_2_modExp_1_while_C_27,
      COMP_LOOP_2_modExp_1_while_C_28, COMP_LOOP_2_modExp_1_while_C_29, COMP_LOOP_2_modExp_1_while_C_30,
      COMP_LOOP_2_modExp_1_while_C_31, COMP_LOOP_2_modExp_1_while_C_32, COMP_LOOP_2_modExp_1_while_C_33,
      COMP_LOOP_2_modExp_1_while_C_34, COMP_LOOP_2_modExp_1_while_C_35, COMP_LOOP_2_modExp_1_while_C_36,
      COMP_LOOP_2_modExp_1_while_C_37, COMP_LOOP_2_modExp_1_while_C_38, COMP_LOOP_C_66,
      COMP_LOOP_C_67, COMP_LOOP_C_68, COMP_LOOP_C_69, COMP_LOOP_C_70, COMP_LOOP_C_71,
      COMP_LOOP_C_72, COMP_LOOP_C_73, COMP_LOOP_C_74, COMP_LOOP_C_75, COMP_LOOP_C_76,
      COMP_LOOP_C_77, COMP_LOOP_C_78, COMP_LOOP_C_79, COMP_LOOP_C_80, COMP_LOOP_C_81,
      COMP_LOOP_C_82, COMP_LOOP_C_83, COMP_LOOP_C_84, COMP_LOOP_C_85, COMP_LOOP_C_86,
      COMP_LOOP_C_87, COMP_LOOP_C_88, COMP_LOOP_C_89, COMP_LOOP_C_90, COMP_LOOP_C_91,
      COMP_LOOP_C_92, COMP_LOOP_C_93, COMP_LOOP_C_94, COMP_LOOP_C_95, COMP_LOOP_C_96,
      COMP_LOOP_C_97, COMP_LOOP_C_98, COMP_LOOP_C_99, COMP_LOOP_C_100, COMP_LOOP_C_101,
      COMP_LOOP_C_102, COMP_LOOP_C_103, COMP_LOOP_C_104, COMP_LOOP_C_105, COMP_LOOP_C_106,
      COMP_LOOP_C_107, COMP_LOOP_C_108, COMP_LOOP_C_109, COMP_LOOP_C_110, COMP_LOOP_C_111,
      COMP_LOOP_C_112, COMP_LOOP_C_113, COMP_LOOP_C_114, COMP_LOOP_C_115, COMP_LOOP_C_116,
      COMP_LOOP_C_117, COMP_LOOP_C_118, COMP_LOOP_C_119, COMP_LOOP_C_120, COMP_LOOP_C_121,
      COMP_LOOP_C_122, COMP_LOOP_C_123, COMP_LOOP_C_124, COMP_LOOP_C_125, COMP_LOOP_C_126,
      COMP_LOOP_C_127, COMP_LOOP_C_128, COMP_LOOP_C_129, COMP_LOOP_3_modExp_1_while_C_0,
      COMP_LOOP_3_modExp_1_while_C_1, COMP_LOOP_3_modExp_1_while_C_2, COMP_LOOP_3_modExp_1_while_C_3,
      COMP_LOOP_3_modExp_1_while_C_4, COMP_LOOP_3_modExp_1_while_C_5, COMP_LOOP_3_modExp_1_while_C_6,
      COMP_LOOP_3_modExp_1_while_C_7, COMP_LOOP_3_modExp_1_while_C_8, COMP_LOOP_3_modExp_1_while_C_9,
      COMP_LOOP_3_modExp_1_while_C_10, COMP_LOOP_3_modExp_1_while_C_11, COMP_LOOP_3_modExp_1_while_C_12,
      COMP_LOOP_3_modExp_1_while_C_13, COMP_LOOP_3_modExp_1_while_C_14, COMP_LOOP_3_modExp_1_while_C_15,
      COMP_LOOP_3_modExp_1_while_C_16, COMP_LOOP_3_modExp_1_while_C_17, COMP_LOOP_3_modExp_1_while_C_18,
      COMP_LOOP_3_modExp_1_while_C_19, COMP_LOOP_3_modExp_1_while_C_20, COMP_LOOP_3_modExp_1_while_C_21,
      COMP_LOOP_3_modExp_1_while_C_22, COMP_LOOP_3_modExp_1_while_C_23, COMP_LOOP_3_modExp_1_while_C_24,
      COMP_LOOP_3_modExp_1_while_C_25, COMP_LOOP_3_modExp_1_while_C_26, COMP_LOOP_3_modExp_1_while_C_27,
      COMP_LOOP_3_modExp_1_while_C_28, COMP_LOOP_3_modExp_1_while_C_29, COMP_LOOP_3_modExp_1_while_C_30,
      COMP_LOOP_3_modExp_1_while_C_31, COMP_LOOP_3_modExp_1_while_C_32, COMP_LOOP_3_modExp_1_while_C_33,
      COMP_LOOP_3_modExp_1_while_C_34, COMP_LOOP_3_modExp_1_while_C_35, COMP_LOOP_3_modExp_1_while_C_36,
      COMP_LOOP_3_modExp_1_while_C_37, COMP_LOOP_3_modExp_1_while_C_38, COMP_LOOP_C_130,
      COMP_LOOP_C_131, COMP_LOOP_C_132, COMP_LOOP_C_133, COMP_LOOP_C_134, COMP_LOOP_C_135,
      COMP_LOOP_C_136, COMP_LOOP_C_137, COMP_LOOP_C_138, COMP_LOOP_C_139, COMP_LOOP_C_140,
      COMP_LOOP_C_141, COMP_LOOP_C_142, COMP_LOOP_C_143, COMP_LOOP_C_144, COMP_LOOP_C_145,
      COMP_LOOP_C_146, COMP_LOOP_C_147, COMP_LOOP_C_148, COMP_LOOP_C_149, COMP_LOOP_C_150,
      COMP_LOOP_C_151, COMP_LOOP_C_152, COMP_LOOP_C_153, COMP_LOOP_C_154, COMP_LOOP_C_155,
      COMP_LOOP_C_156, COMP_LOOP_C_157, COMP_LOOP_C_158, COMP_LOOP_C_159, COMP_LOOP_C_160,
      COMP_LOOP_C_161, COMP_LOOP_C_162, COMP_LOOP_C_163, COMP_LOOP_C_164, COMP_LOOP_C_165,
      COMP_LOOP_C_166, COMP_LOOP_C_167, COMP_LOOP_C_168, COMP_LOOP_C_169, COMP_LOOP_C_170,
      COMP_LOOP_C_171, COMP_LOOP_C_172, COMP_LOOP_C_173, COMP_LOOP_C_174, COMP_LOOP_C_175,
      COMP_LOOP_C_176, COMP_LOOP_C_177, COMP_LOOP_C_178, COMP_LOOP_C_179, COMP_LOOP_C_180,
      COMP_LOOP_C_181, COMP_LOOP_C_182, COMP_LOOP_C_183, COMP_LOOP_C_184, COMP_LOOP_C_185,
      COMP_LOOP_C_186, COMP_LOOP_C_187, COMP_LOOP_C_188, COMP_LOOP_C_189, COMP_LOOP_C_190,
      COMP_LOOP_C_191, COMP_LOOP_C_192, COMP_LOOP_C_193, COMP_LOOP_4_modExp_1_while_C_0,
      COMP_LOOP_4_modExp_1_while_C_1, COMP_LOOP_4_modExp_1_while_C_2, COMP_LOOP_4_modExp_1_while_C_3,
      COMP_LOOP_4_modExp_1_while_C_4, COMP_LOOP_4_modExp_1_while_C_5, COMP_LOOP_4_modExp_1_while_C_6,
      COMP_LOOP_4_modExp_1_while_C_7, COMP_LOOP_4_modExp_1_while_C_8, COMP_LOOP_4_modExp_1_while_C_9,
      COMP_LOOP_4_modExp_1_while_C_10, COMP_LOOP_4_modExp_1_while_C_11, COMP_LOOP_4_modExp_1_while_C_12,
      COMP_LOOP_4_modExp_1_while_C_13, COMP_LOOP_4_modExp_1_while_C_14, COMP_LOOP_4_modExp_1_while_C_15,
      COMP_LOOP_4_modExp_1_while_C_16, COMP_LOOP_4_modExp_1_while_C_17, COMP_LOOP_4_modExp_1_while_C_18,
      COMP_LOOP_4_modExp_1_while_C_19, COMP_LOOP_4_modExp_1_while_C_20, COMP_LOOP_4_modExp_1_while_C_21,
      COMP_LOOP_4_modExp_1_while_C_22, COMP_LOOP_4_modExp_1_while_C_23, COMP_LOOP_4_modExp_1_while_C_24,
      COMP_LOOP_4_modExp_1_while_C_25, COMP_LOOP_4_modExp_1_while_C_26, COMP_LOOP_4_modExp_1_while_C_27,
      COMP_LOOP_4_modExp_1_while_C_28, COMP_LOOP_4_modExp_1_while_C_29, COMP_LOOP_4_modExp_1_while_C_30,
      COMP_LOOP_4_modExp_1_while_C_31, COMP_LOOP_4_modExp_1_while_C_32, COMP_LOOP_4_modExp_1_while_C_33,
      COMP_LOOP_4_modExp_1_while_C_34, COMP_LOOP_4_modExp_1_while_C_35, COMP_LOOP_4_modExp_1_while_C_36,
      COMP_LOOP_4_modExp_1_while_C_37, COMP_LOOP_4_modExp_1_while_C_38, COMP_LOOP_C_194,
      COMP_LOOP_C_195, COMP_LOOP_C_196, COMP_LOOP_C_197, COMP_LOOP_C_198, COMP_LOOP_C_199,
      COMP_LOOP_C_200, COMP_LOOP_C_201, COMP_LOOP_C_202, COMP_LOOP_C_203, COMP_LOOP_C_204,
      COMP_LOOP_C_205, COMP_LOOP_C_206, COMP_LOOP_C_207, COMP_LOOP_C_208, COMP_LOOP_C_209,
      COMP_LOOP_C_210, COMP_LOOP_C_211, COMP_LOOP_C_212, COMP_LOOP_C_213, COMP_LOOP_C_214,
      COMP_LOOP_C_215, COMP_LOOP_C_216, COMP_LOOP_C_217, COMP_LOOP_C_218, COMP_LOOP_C_219,
      COMP_LOOP_C_220, COMP_LOOP_C_221, COMP_LOOP_C_222, COMP_LOOP_C_223, COMP_LOOP_C_224,
      COMP_LOOP_C_225, COMP_LOOP_C_226, COMP_LOOP_C_227, COMP_LOOP_C_228, COMP_LOOP_C_229,
      COMP_LOOP_C_230, COMP_LOOP_C_231, COMP_LOOP_C_232, COMP_LOOP_C_233, COMP_LOOP_C_234,
      COMP_LOOP_C_235, COMP_LOOP_C_236, COMP_LOOP_C_237, COMP_LOOP_C_238, COMP_LOOP_C_239,
      COMP_LOOP_C_240, COMP_LOOP_C_241, COMP_LOOP_C_242, COMP_LOOP_C_243, COMP_LOOP_C_244,
      COMP_LOOP_C_245, COMP_LOOP_C_246, COMP_LOOP_C_247, COMP_LOOP_C_248, COMP_LOOP_C_249,
      COMP_LOOP_C_250, COMP_LOOP_C_251, COMP_LOOP_C_252, COMP_LOOP_C_253, COMP_LOOP_C_254,
      COMP_LOOP_C_255, COMP_LOOP_C_256, COMP_LOOP_C_257, COMP_LOOP_5_modExp_1_while_C_0,
      COMP_LOOP_5_modExp_1_while_C_1, COMP_LOOP_5_modExp_1_while_C_2, COMP_LOOP_5_modExp_1_while_C_3,
      COMP_LOOP_5_modExp_1_while_C_4, COMP_LOOP_5_modExp_1_while_C_5, COMP_LOOP_5_modExp_1_while_C_6,
      COMP_LOOP_5_modExp_1_while_C_7, COMP_LOOP_5_modExp_1_while_C_8, COMP_LOOP_5_modExp_1_while_C_9,
      COMP_LOOP_5_modExp_1_while_C_10, COMP_LOOP_5_modExp_1_while_C_11, COMP_LOOP_5_modExp_1_while_C_12,
      COMP_LOOP_5_modExp_1_while_C_13, COMP_LOOP_5_modExp_1_while_C_14, COMP_LOOP_5_modExp_1_while_C_15,
      COMP_LOOP_5_modExp_1_while_C_16, COMP_LOOP_5_modExp_1_while_C_17, COMP_LOOP_5_modExp_1_while_C_18,
      COMP_LOOP_5_modExp_1_while_C_19, COMP_LOOP_5_modExp_1_while_C_20, COMP_LOOP_5_modExp_1_while_C_21,
      COMP_LOOP_5_modExp_1_while_C_22, COMP_LOOP_5_modExp_1_while_C_23, COMP_LOOP_5_modExp_1_while_C_24,
      COMP_LOOP_5_modExp_1_while_C_25, COMP_LOOP_5_modExp_1_while_C_26, COMP_LOOP_5_modExp_1_while_C_27,
      COMP_LOOP_5_modExp_1_while_C_28, COMP_LOOP_5_modExp_1_while_C_29, COMP_LOOP_5_modExp_1_while_C_30,
      COMP_LOOP_5_modExp_1_while_C_31, COMP_LOOP_5_modExp_1_while_C_32, COMP_LOOP_5_modExp_1_while_C_33,
      COMP_LOOP_5_modExp_1_while_C_34, COMP_LOOP_5_modExp_1_while_C_35, COMP_LOOP_5_modExp_1_while_C_36,
      COMP_LOOP_5_modExp_1_while_C_37, COMP_LOOP_5_modExp_1_while_C_38, COMP_LOOP_C_258,
      COMP_LOOP_C_259, COMP_LOOP_C_260, COMP_LOOP_C_261, COMP_LOOP_C_262, COMP_LOOP_C_263,
      COMP_LOOP_C_264, COMP_LOOP_C_265, COMP_LOOP_C_266, COMP_LOOP_C_267, COMP_LOOP_C_268,
      COMP_LOOP_C_269, COMP_LOOP_C_270, COMP_LOOP_C_271, COMP_LOOP_C_272, COMP_LOOP_C_273,
      COMP_LOOP_C_274, COMP_LOOP_C_275, COMP_LOOP_C_276, COMP_LOOP_C_277, COMP_LOOP_C_278,
      COMP_LOOP_C_279, COMP_LOOP_C_280, COMP_LOOP_C_281, COMP_LOOP_C_282, COMP_LOOP_C_283,
      COMP_LOOP_C_284, COMP_LOOP_C_285, COMP_LOOP_C_286, COMP_LOOP_C_287, COMP_LOOP_C_288,
      COMP_LOOP_C_289, COMP_LOOP_C_290, COMP_LOOP_C_291, COMP_LOOP_C_292, COMP_LOOP_C_293,
      COMP_LOOP_C_294, COMP_LOOP_C_295, COMP_LOOP_C_296, COMP_LOOP_C_297, COMP_LOOP_C_298,
      COMP_LOOP_C_299, COMP_LOOP_C_300, COMP_LOOP_C_301, COMP_LOOP_C_302, COMP_LOOP_C_303,
      COMP_LOOP_C_304, COMP_LOOP_C_305, COMP_LOOP_C_306, COMP_LOOP_C_307, COMP_LOOP_C_308,
      COMP_LOOP_C_309, COMP_LOOP_C_310, COMP_LOOP_C_311, COMP_LOOP_C_312, COMP_LOOP_C_313,
      COMP_LOOP_C_314, COMP_LOOP_C_315, COMP_LOOP_C_316, COMP_LOOP_C_317, COMP_LOOP_C_318,
      COMP_LOOP_C_319, COMP_LOOP_C_320, COMP_LOOP_C_321, COMP_LOOP_6_modExp_1_while_C_0,
      COMP_LOOP_6_modExp_1_while_C_1, COMP_LOOP_6_modExp_1_while_C_2, COMP_LOOP_6_modExp_1_while_C_3,
      COMP_LOOP_6_modExp_1_while_C_4, COMP_LOOP_6_modExp_1_while_C_5, COMP_LOOP_6_modExp_1_while_C_6,
      COMP_LOOP_6_modExp_1_while_C_7, COMP_LOOP_6_modExp_1_while_C_8, COMP_LOOP_6_modExp_1_while_C_9,
      COMP_LOOP_6_modExp_1_while_C_10, COMP_LOOP_6_modExp_1_while_C_11, COMP_LOOP_6_modExp_1_while_C_12,
      COMP_LOOP_6_modExp_1_while_C_13, COMP_LOOP_6_modExp_1_while_C_14, COMP_LOOP_6_modExp_1_while_C_15,
      COMP_LOOP_6_modExp_1_while_C_16, COMP_LOOP_6_modExp_1_while_C_17, COMP_LOOP_6_modExp_1_while_C_18,
      COMP_LOOP_6_modExp_1_while_C_19, COMP_LOOP_6_modExp_1_while_C_20, COMP_LOOP_6_modExp_1_while_C_21,
      COMP_LOOP_6_modExp_1_while_C_22, COMP_LOOP_6_modExp_1_while_C_23, COMP_LOOP_6_modExp_1_while_C_24,
      COMP_LOOP_6_modExp_1_while_C_25, COMP_LOOP_6_modExp_1_while_C_26, COMP_LOOP_6_modExp_1_while_C_27,
      COMP_LOOP_6_modExp_1_while_C_28, COMP_LOOP_6_modExp_1_while_C_29, COMP_LOOP_6_modExp_1_while_C_30,
      COMP_LOOP_6_modExp_1_while_C_31, COMP_LOOP_6_modExp_1_while_C_32, COMP_LOOP_6_modExp_1_while_C_33,
      COMP_LOOP_6_modExp_1_while_C_34, COMP_LOOP_6_modExp_1_while_C_35, COMP_LOOP_6_modExp_1_while_C_36,
      COMP_LOOP_6_modExp_1_while_C_37, COMP_LOOP_6_modExp_1_while_C_38, COMP_LOOP_C_322,
      COMP_LOOP_C_323, COMP_LOOP_C_324, COMP_LOOP_C_325, COMP_LOOP_C_326, COMP_LOOP_C_327,
      COMP_LOOP_C_328, COMP_LOOP_C_329, COMP_LOOP_C_330, COMP_LOOP_C_331, COMP_LOOP_C_332,
      COMP_LOOP_C_333, COMP_LOOP_C_334, COMP_LOOP_C_335, COMP_LOOP_C_336, COMP_LOOP_C_337,
      COMP_LOOP_C_338, COMP_LOOP_C_339, COMP_LOOP_C_340, COMP_LOOP_C_341, COMP_LOOP_C_342,
      COMP_LOOP_C_343, COMP_LOOP_C_344, COMP_LOOP_C_345, COMP_LOOP_C_346, COMP_LOOP_C_347,
      COMP_LOOP_C_348, COMP_LOOP_C_349, COMP_LOOP_C_350, COMP_LOOP_C_351, COMP_LOOP_C_352,
      COMP_LOOP_C_353, COMP_LOOP_C_354, COMP_LOOP_C_355, COMP_LOOP_C_356, COMP_LOOP_C_357,
      COMP_LOOP_C_358, COMP_LOOP_C_359, COMP_LOOP_C_360, COMP_LOOP_C_361, COMP_LOOP_C_362,
      COMP_LOOP_C_363, COMP_LOOP_C_364, COMP_LOOP_C_365, COMP_LOOP_C_366, COMP_LOOP_C_367,
      COMP_LOOP_C_368, COMP_LOOP_C_369, COMP_LOOP_C_370, COMP_LOOP_C_371, COMP_LOOP_C_372,
      COMP_LOOP_C_373, COMP_LOOP_C_374, COMP_LOOP_C_375, COMP_LOOP_C_376, COMP_LOOP_C_377,
      COMP_LOOP_C_378, COMP_LOOP_C_379, COMP_LOOP_C_380, COMP_LOOP_C_381, COMP_LOOP_C_382,
      COMP_LOOP_C_383, COMP_LOOP_C_384, COMP_LOOP_C_385, COMP_LOOP_7_modExp_1_while_C_0,
      COMP_LOOP_7_modExp_1_while_C_1, COMP_LOOP_7_modExp_1_while_C_2, COMP_LOOP_7_modExp_1_while_C_3,
      COMP_LOOP_7_modExp_1_while_C_4, COMP_LOOP_7_modExp_1_while_C_5, COMP_LOOP_7_modExp_1_while_C_6,
      COMP_LOOP_7_modExp_1_while_C_7, COMP_LOOP_7_modExp_1_while_C_8, COMP_LOOP_7_modExp_1_while_C_9,
      COMP_LOOP_7_modExp_1_while_C_10, COMP_LOOP_7_modExp_1_while_C_11, COMP_LOOP_7_modExp_1_while_C_12,
      COMP_LOOP_7_modExp_1_while_C_13, COMP_LOOP_7_modExp_1_while_C_14, COMP_LOOP_7_modExp_1_while_C_15,
      COMP_LOOP_7_modExp_1_while_C_16, COMP_LOOP_7_modExp_1_while_C_17, COMP_LOOP_7_modExp_1_while_C_18,
      COMP_LOOP_7_modExp_1_while_C_19, COMP_LOOP_7_modExp_1_while_C_20, COMP_LOOP_7_modExp_1_while_C_21,
      COMP_LOOP_7_modExp_1_while_C_22, COMP_LOOP_7_modExp_1_while_C_23, COMP_LOOP_7_modExp_1_while_C_24,
      COMP_LOOP_7_modExp_1_while_C_25, COMP_LOOP_7_modExp_1_while_C_26, COMP_LOOP_7_modExp_1_while_C_27,
      COMP_LOOP_7_modExp_1_while_C_28, COMP_LOOP_7_modExp_1_while_C_29, COMP_LOOP_7_modExp_1_while_C_30,
      COMP_LOOP_7_modExp_1_while_C_31, COMP_LOOP_7_modExp_1_while_C_32, COMP_LOOP_7_modExp_1_while_C_33,
      COMP_LOOP_7_modExp_1_while_C_34, COMP_LOOP_7_modExp_1_while_C_35, COMP_LOOP_7_modExp_1_while_C_36,
      COMP_LOOP_7_modExp_1_while_C_37, COMP_LOOP_7_modExp_1_while_C_38, COMP_LOOP_C_386,
      COMP_LOOP_C_387, COMP_LOOP_C_388, COMP_LOOP_C_389, COMP_LOOP_C_390, COMP_LOOP_C_391,
      COMP_LOOP_C_392, COMP_LOOP_C_393, COMP_LOOP_C_394, COMP_LOOP_C_395, COMP_LOOP_C_396,
      COMP_LOOP_C_397, COMP_LOOP_C_398, COMP_LOOP_C_399, COMP_LOOP_C_400, COMP_LOOP_C_401,
      COMP_LOOP_C_402, COMP_LOOP_C_403, COMP_LOOP_C_404, COMP_LOOP_C_405, COMP_LOOP_C_406,
      COMP_LOOP_C_407, COMP_LOOP_C_408, COMP_LOOP_C_409, COMP_LOOP_C_410, COMP_LOOP_C_411,
      COMP_LOOP_C_412, COMP_LOOP_C_413, COMP_LOOP_C_414, COMP_LOOP_C_415, COMP_LOOP_C_416,
      COMP_LOOP_C_417, COMP_LOOP_C_418, COMP_LOOP_C_419, COMP_LOOP_C_420, COMP_LOOP_C_421,
      COMP_LOOP_C_422, COMP_LOOP_C_423, COMP_LOOP_C_424, COMP_LOOP_C_425, COMP_LOOP_C_426,
      COMP_LOOP_C_427, COMP_LOOP_C_428, COMP_LOOP_C_429, COMP_LOOP_C_430, COMP_LOOP_C_431,
      COMP_LOOP_C_432, COMP_LOOP_C_433, COMP_LOOP_C_434, COMP_LOOP_C_435, COMP_LOOP_C_436,
      COMP_LOOP_C_437, COMP_LOOP_C_438, COMP_LOOP_C_439, COMP_LOOP_C_440, COMP_LOOP_C_441,
      COMP_LOOP_C_442, COMP_LOOP_C_443, COMP_LOOP_C_444, COMP_LOOP_C_445, COMP_LOOP_C_446,
      COMP_LOOP_C_447, COMP_LOOP_C_448, COMP_LOOP_C_449, COMP_LOOP_8_modExp_1_while_C_0,
      COMP_LOOP_8_modExp_1_while_C_1, COMP_LOOP_8_modExp_1_while_C_2, COMP_LOOP_8_modExp_1_while_C_3,
      COMP_LOOP_8_modExp_1_while_C_4, COMP_LOOP_8_modExp_1_while_C_5, COMP_LOOP_8_modExp_1_while_C_6,
      COMP_LOOP_8_modExp_1_while_C_7, COMP_LOOP_8_modExp_1_while_C_8, COMP_LOOP_8_modExp_1_while_C_9,
      COMP_LOOP_8_modExp_1_while_C_10, COMP_LOOP_8_modExp_1_while_C_11, COMP_LOOP_8_modExp_1_while_C_12,
      COMP_LOOP_8_modExp_1_while_C_13, COMP_LOOP_8_modExp_1_while_C_14, COMP_LOOP_8_modExp_1_while_C_15,
      COMP_LOOP_8_modExp_1_while_C_16, COMP_LOOP_8_modExp_1_while_C_17, COMP_LOOP_8_modExp_1_while_C_18,
      COMP_LOOP_8_modExp_1_while_C_19, COMP_LOOP_8_modExp_1_while_C_20, COMP_LOOP_8_modExp_1_while_C_21,
      COMP_LOOP_8_modExp_1_while_C_22, COMP_LOOP_8_modExp_1_while_C_23, COMP_LOOP_8_modExp_1_while_C_24,
      COMP_LOOP_8_modExp_1_while_C_25, COMP_LOOP_8_modExp_1_while_C_26, COMP_LOOP_8_modExp_1_while_C_27,
      COMP_LOOP_8_modExp_1_while_C_28, COMP_LOOP_8_modExp_1_while_C_29, COMP_LOOP_8_modExp_1_while_C_30,
      COMP_LOOP_8_modExp_1_while_C_31, COMP_LOOP_8_modExp_1_while_C_32, COMP_LOOP_8_modExp_1_while_C_33,
      COMP_LOOP_8_modExp_1_while_C_34, COMP_LOOP_8_modExp_1_while_C_35, COMP_LOOP_8_modExp_1_while_C_36,
      COMP_LOOP_8_modExp_1_while_C_37, COMP_LOOP_8_modExp_1_while_C_38, COMP_LOOP_C_450,
      COMP_LOOP_C_451, COMP_LOOP_C_452, COMP_LOOP_C_453, COMP_LOOP_C_454, COMP_LOOP_C_455,
      COMP_LOOP_C_456, COMP_LOOP_C_457, COMP_LOOP_C_458, COMP_LOOP_C_459, COMP_LOOP_C_460,
      COMP_LOOP_C_461, COMP_LOOP_C_462, COMP_LOOP_C_463, COMP_LOOP_C_464, COMP_LOOP_C_465,
      COMP_LOOP_C_466, COMP_LOOP_C_467, COMP_LOOP_C_468, COMP_LOOP_C_469, COMP_LOOP_C_470,
      COMP_LOOP_C_471, COMP_LOOP_C_472, COMP_LOOP_C_473, COMP_LOOP_C_474, COMP_LOOP_C_475,
      COMP_LOOP_C_476, COMP_LOOP_C_477, COMP_LOOP_C_478, COMP_LOOP_C_479, COMP_LOOP_C_480,
      COMP_LOOP_C_481, COMP_LOOP_C_482, COMP_LOOP_C_483, COMP_LOOP_C_484, COMP_LOOP_C_485,
      COMP_LOOP_C_486, COMP_LOOP_C_487, COMP_LOOP_C_488, COMP_LOOP_C_489, COMP_LOOP_C_490,
      COMP_LOOP_C_491, COMP_LOOP_C_492, COMP_LOOP_C_493, COMP_LOOP_C_494, COMP_LOOP_C_495,
      COMP_LOOP_C_496, COMP_LOOP_C_497, COMP_LOOP_C_498, COMP_LOOP_C_499, COMP_LOOP_C_500,
      COMP_LOOP_C_501, COMP_LOOP_C_502, COMP_LOOP_C_503, COMP_LOOP_C_504, COMP_LOOP_C_505,
      COMP_LOOP_C_506, COMP_LOOP_C_507, COMP_LOOP_C_508, COMP_LOOP_C_509, COMP_LOOP_C_510,
      COMP_LOOP_C_511, COMP_LOOP_C_512, COMP_LOOP_C_513, COMP_LOOP_9_modExp_1_while_C_0,
      COMP_LOOP_9_modExp_1_while_C_1, COMP_LOOP_9_modExp_1_while_C_2, COMP_LOOP_9_modExp_1_while_C_3,
      COMP_LOOP_9_modExp_1_while_C_4, COMP_LOOP_9_modExp_1_while_C_5, COMP_LOOP_9_modExp_1_while_C_6,
      COMP_LOOP_9_modExp_1_while_C_7, COMP_LOOP_9_modExp_1_while_C_8, COMP_LOOP_9_modExp_1_while_C_9,
      COMP_LOOP_9_modExp_1_while_C_10, COMP_LOOP_9_modExp_1_while_C_11, COMP_LOOP_9_modExp_1_while_C_12,
      COMP_LOOP_9_modExp_1_while_C_13, COMP_LOOP_9_modExp_1_while_C_14, COMP_LOOP_9_modExp_1_while_C_15,
      COMP_LOOP_9_modExp_1_while_C_16, COMP_LOOP_9_modExp_1_while_C_17, COMP_LOOP_9_modExp_1_while_C_18,
      COMP_LOOP_9_modExp_1_while_C_19, COMP_LOOP_9_modExp_1_while_C_20, COMP_LOOP_9_modExp_1_while_C_21,
      COMP_LOOP_9_modExp_1_while_C_22, COMP_LOOP_9_modExp_1_while_C_23, COMP_LOOP_9_modExp_1_while_C_24,
      COMP_LOOP_9_modExp_1_while_C_25, COMP_LOOP_9_modExp_1_while_C_26, COMP_LOOP_9_modExp_1_while_C_27,
      COMP_LOOP_9_modExp_1_while_C_28, COMP_LOOP_9_modExp_1_while_C_29, COMP_LOOP_9_modExp_1_while_C_30,
      COMP_LOOP_9_modExp_1_while_C_31, COMP_LOOP_9_modExp_1_while_C_32, COMP_LOOP_9_modExp_1_while_C_33,
      COMP_LOOP_9_modExp_1_while_C_34, COMP_LOOP_9_modExp_1_while_C_35, COMP_LOOP_9_modExp_1_while_C_36,
      COMP_LOOP_9_modExp_1_while_C_37, COMP_LOOP_9_modExp_1_while_C_38, COMP_LOOP_C_514,
      COMP_LOOP_C_515, COMP_LOOP_C_516, COMP_LOOP_C_517, COMP_LOOP_C_518, COMP_LOOP_C_519,
      COMP_LOOP_C_520, COMP_LOOP_C_521, COMP_LOOP_C_522, COMP_LOOP_C_523, COMP_LOOP_C_524,
      COMP_LOOP_C_525, COMP_LOOP_C_526, COMP_LOOP_C_527, COMP_LOOP_C_528, COMP_LOOP_C_529,
      COMP_LOOP_C_530, COMP_LOOP_C_531, COMP_LOOP_C_532, COMP_LOOP_C_533, COMP_LOOP_C_534,
      COMP_LOOP_C_535, COMP_LOOP_C_536, COMP_LOOP_C_537, COMP_LOOP_C_538, COMP_LOOP_C_539,
      COMP_LOOP_C_540, COMP_LOOP_C_541, COMP_LOOP_C_542, COMP_LOOP_C_543, COMP_LOOP_C_544,
      COMP_LOOP_C_545, COMP_LOOP_C_546, COMP_LOOP_C_547, COMP_LOOP_C_548, COMP_LOOP_C_549,
      COMP_LOOP_C_550, COMP_LOOP_C_551, COMP_LOOP_C_552, COMP_LOOP_C_553, COMP_LOOP_C_554,
      COMP_LOOP_C_555, COMP_LOOP_C_556, COMP_LOOP_C_557, COMP_LOOP_C_558, COMP_LOOP_C_559,
      COMP_LOOP_C_560, COMP_LOOP_C_561, COMP_LOOP_C_562, COMP_LOOP_C_563, COMP_LOOP_C_564,
      COMP_LOOP_C_565, COMP_LOOP_C_566, COMP_LOOP_C_567, COMP_LOOP_C_568, COMP_LOOP_C_569,
      COMP_LOOP_C_570, COMP_LOOP_C_571, COMP_LOOP_C_572, COMP_LOOP_C_573, COMP_LOOP_C_574,
      COMP_LOOP_C_575, COMP_LOOP_C_576, COMP_LOOP_C_577, COMP_LOOP_10_modExp_1_while_C_0,
      COMP_LOOP_10_modExp_1_while_C_1, COMP_LOOP_10_modExp_1_while_C_2, COMP_LOOP_10_modExp_1_while_C_3,
      COMP_LOOP_10_modExp_1_while_C_4, COMP_LOOP_10_modExp_1_while_C_5, COMP_LOOP_10_modExp_1_while_C_6,
      COMP_LOOP_10_modExp_1_while_C_7, COMP_LOOP_10_modExp_1_while_C_8, COMP_LOOP_10_modExp_1_while_C_9,
      COMP_LOOP_10_modExp_1_while_C_10, COMP_LOOP_10_modExp_1_while_C_11, COMP_LOOP_10_modExp_1_while_C_12,
      COMP_LOOP_10_modExp_1_while_C_13, COMP_LOOP_10_modExp_1_while_C_14, COMP_LOOP_10_modExp_1_while_C_15,
      COMP_LOOP_10_modExp_1_while_C_16, COMP_LOOP_10_modExp_1_while_C_17, COMP_LOOP_10_modExp_1_while_C_18,
      COMP_LOOP_10_modExp_1_while_C_19, COMP_LOOP_10_modExp_1_while_C_20, COMP_LOOP_10_modExp_1_while_C_21,
      COMP_LOOP_10_modExp_1_while_C_22, COMP_LOOP_10_modExp_1_while_C_23, COMP_LOOP_10_modExp_1_while_C_24,
      COMP_LOOP_10_modExp_1_while_C_25, COMP_LOOP_10_modExp_1_while_C_26, COMP_LOOP_10_modExp_1_while_C_27,
      COMP_LOOP_10_modExp_1_while_C_28, COMP_LOOP_10_modExp_1_while_C_29, COMP_LOOP_10_modExp_1_while_C_30,
      COMP_LOOP_10_modExp_1_while_C_31, COMP_LOOP_10_modExp_1_while_C_32, COMP_LOOP_10_modExp_1_while_C_33,
      COMP_LOOP_10_modExp_1_while_C_34, COMP_LOOP_10_modExp_1_while_C_35, COMP_LOOP_10_modExp_1_while_C_36,
      COMP_LOOP_10_modExp_1_while_C_37, COMP_LOOP_10_modExp_1_while_C_38, COMP_LOOP_C_578,
      COMP_LOOP_C_579, COMP_LOOP_C_580, COMP_LOOP_C_581, COMP_LOOP_C_582, COMP_LOOP_C_583,
      COMP_LOOP_C_584, COMP_LOOP_C_585, COMP_LOOP_C_586, COMP_LOOP_C_587, COMP_LOOP_C_588,
      COMP_LOOP_C_589, COMP_LOOP_C_590, COMP_LOOP_C_591, COMP_LOOP_C_592, COMP_LOOP_C_593,
      COMP_LOOP_C_594, COMP_LOOP_C_595, COMP_LOOP_C_596, COMP_LOOP_C_597, COMP_LOOP_C_598,
      COMP_LOOP_C_599, COMP_LOOP_C_600, COMP_LOOP_C_601, COMP_LOOP_C_602, COMP_LOOP_C_603,
      COMP_LOOP_C_604, COMP_LOOP_C_605, COMP_LOOP_C_606, COMP_LOOP_C_607, COMP_LOOP_C_608,
      COMP_LOOP_C_609, COMP_LOOP_C_610, COMP_LOOP_C_611, COMP_LOOP_C_612, COMP_LOOP_C_613,
      COMP_LOOP_C_614, COMP_LOOP_C_615, COMP_LOOP_C_616, COMP_LOOP_C_617, COMP_LOOP_C_618,
      COMP_LOOP_C_619, COMP_LOOP_C_620, COMP_LOOP_C_621, COMP_LOOP_C_622, COMP_LOOP_C_623,
      COMP_LOOP_C_624, COMP_LOOP_C_625, COMP_LOOP_C_626, COMP_LOOP_C_627, COMP_LOOP_C_628,
      COMP_LOOP_C_629, COMP_LOOP_C_630, COMP_LOOP_C_631, COMP_LOOP_C_632, COMP_LOOP_C_633,
      COMP_LOOP_C_634, COMP_LOOP_C_635, COMP_LOOP_C_636, COMP_LOOP_C_637, COMP_LOOP_C_638,
      COMP_LOOP_C_639, COMP_LOOP_C_640, COMP_LOOP_C_641, COMP_LOOP_11_modExp_1_while_C_0,
      COMP_LOOP_11_modExp_1_while_C_1, COMP_LOOP_11_modExp_1_while_C_2, COMP_LOOP_11_modExp_1_while_C_3,
      COMP_LOOP_11_modExp_1_while_C_4, COMP_LOOP_11_modExp_1_while_C_5, COMP_LOOP_11_modExp_1_while_C_6,
      COMP_LOOP_11_modExp_1_while_C_7, COMP_LOOP_11_modExp_1_while_C_8, COMP_LOOP_11_modExp_1_while_C_9,
      COMP_LOOP_11_modExp_1_while_C_10, COMP_LOOP_11_modExp_1_while_C_11, COMP_LOOP_11_modExp_1_while_C_12,
      COMP_LOOP_11_modExp_1_while_C_13, COMP_LOOP_11_modExp_1_while_C_14, COMP_LOOP_11_modExp_1_while_C_15,
      COMP_LOOP_11_modExp_1_while_C_16, COMP_LOOP_11_modExp_1_while_C_17, COMP_LOOP_11_modExp_1_while_C_18,
      COMP_LOOP_11_modExp_1_while_C_19, COMP_LOOP_11_modExp_1_while_C_20, COMP_LOOP_11_modExp_1_while_C_21,
      COMP_LOOP_11_modExp_1_while_C_22, COMP_LOOP_11_modExp_1_while_C_23, COMP_LOOP_11_modExp_1_while_C_24,
      COMP_LOOP_11_modExp_1_while_C_25, COMP_LOOP_11_modExp_1_while_C_26, COMP_LOOP_11_modExp_1_while_C_27,
      COMP_LOOP_11_modExp_1_while_C_28, COMP_LOOP_11_modExp_1_while_C_29, COMP_LOOP_11_modExp_1_while_C_30,
      COMP_LOOP_11_modExp_1_while_C_31, COMP_LOOP_11_modExp_1_while_C_32, COMP_LOOP_11_modExp_1_while_C_33,
      COMP_LOOP_11_modExp_1_while_C_34, COMP_LOOP_11_modExp_1_while_C_35, COMP_LOOP_11_modExp_1_while_C_36,
      COMP_LOOP_11_modExp_1_while_C_37, COMP_LOOP_11_modExp_1_while_C_38, COMP_LOOP_C_642,
      COMP_LOOP_C_643, COMP_LOOP_C_644, COMP_LOOP_C_645, COMP_LOOP_C_646, COMP_LOOP_C_647,
      COMP_LOOP_C_648, COMP_LOOP_C_649, COMP_LOOP_C_650, COMP_LOOP_C_651, COMP_LOOP_C_652,
      COMP_LOOP_C_653, COMP_LOOP_C_654, COMP_LOOP_C_655, COMP_LOOP_C_656, COMP_LOOP_C_657,
      COMP_LOOP_C_658, COMP_LOOP_C_659, COMP_LOOP_C_660, COMP_LOOP_C_661, COMP_LOOP_C_662,
      COMP_LOOP_C_663, COMP_LOOP_C_664, COMP_LOOP_C_665, COMP_LOOP_C_666, COMP_LOOP_C_667,
      COMP_LOOP_C_668, COMP_LOOP_C_669, COMP_LOOP_C_670, COMP_LOOP_C_671, COMP_LOOP_C_672,
      COMP_LOOP_C_673, COMP_LOOP_C_674, COMP_LOOP_C_675, COMP_LOOP_C_676, COMP_LOOP_C_677,
      COMP_LOOP_C_678, COMP_LOOP_C_679, COMP_LOOP_C_680, COMP_LOOP_C_681, COMP_LOOP_C_682,
      COMP_LOOP_C_683, COMP_LOOP_C_684, COMP_LOOP_C_685, COMP_LOOP_C_686, COMP_LOOP_C_687,
      COMP_LOOP_C_688, COMP_LOOP_C_689, COMP_LOOP_C_690, COMP_LOOP_C_691, COMP_LOOP_C_692,
      COMP_LOOP_C_693, COMP_LOOP_C_694, COMP_LOOP_C_695, COMP_LOOP_C_696, COMP_LOOP_C_697,
      COMP_LOOP_C_698, COMP_LOOP_C_699, COMP_LOOP_C_700, COMP_LOOP_C_701, COMP_LOOP_C_702,
      COMP_LOOP_C_703, COMP_LOOP_C_704, COMP_LOOP_C_705, COMP_LOOP_12_modExp_1_while_C_0,
      COMP_LOOP_12_modExp_1_while_C_1, COMP_LOOP_12_modExp_1_while_C_2, COMP_LOOP_12_modExp_1_while_C_3,
      COMP_LOOP_12_modExp_1_while_C_4, COMP_LOOP_12_modExp_1_while_C_5, COMP_LOOP_12_modExp_1_while_C_6,
      COMP_LOOP_12_modExp_1_while_C_7, COMP_LOOP_12_modExp_1_while_C_8, COMP_LOOP_12_modExp_1_while_C_9,
      COMP_LOOP_12_modExp_1_while_C_10, COMP_LOOP_12_modExp_1_while_C_11, COMP_LOOP_12_modExp_1_while_C_12,
      COMP_LOOP_12_modExp_1_while_C_13, COMP_LOOP_12_modExp_1_while_C_14, COMP_LOOP_12_modExp_1_while_C_15,
      COMP_LOOP_12_modExp_1_while_C_16, COMP_LOOP_12_modExp_1_while_C_17, COMP_LOOP_12_modExp_1_while_C_18,
      COMP_LOOP_12_modExp_1_while_C_19, COMP_LOOP_12_modExp_1_while_C_20, COMP_LOOP_12_modExp_1_while_C_21,
      COMP_LOOP_12_modExp_1_while_C_22, COMP_LOOP_12_modExp_1_while_C_23, COMP_LOOP_12_modExp_1_while_C_24,
      COMP_LOOP_12_modExp_1_while_C_25, COMP_LOOP_12_modExp_1_while_C_26, COMP_LOOP_12_modExp_1_while_C_27,
      COMP_LOOP_12_modExp_1_while_C_28, COMP_LOOP_12_modExp_1_while_C_29, COMP_LOOP_12_modExp_1_while_C_30,
      COMP_LOOP_12_modExp_1_while_C_31, COMP_LOOP_12_modExp_1_while_C_32, COMP_LOOP_12_modExp_1_while_C_33,
      COMP_LOOP_12_modExp_1_while_C_34, COMP_LOOP_12_modExp_1_while_C_35, COMP_LOOP_12_modExp_1_while_C_36,
      COMP_LOOP_12_modExp_1_while_C_37, COMP_LOOP_12_modExp_1_while_C_38, COMP_LOOP_C_706,
      COMP_LOOP_C_707, COMP_LOOP_C_708, COMP_LOOP_C_709, COMP_LOOP_C_710, COMP_LOOP_C_711,
      COMP_LOOP_C_712, COMP_LOOP_C_713, COMP_LOOP_C_714, COMP_LOOP_C_715, COMP_LOOP_C_716,
      COMP_LOOP_C_717, COMP_LOOP_C_718, COMP_LOOP_C_719, COMP_LOOP_C_720, COMP_LOOP_C_721,
      COMP_LOOP_C_722, COMP_LOOP_C_723, COMP_LOOP_C_724, COMP_LOOP_C_725, COMP_LOOP_C_726,
      COMP_LOOP_C_727, COMP_LOOP_C_728, COMP_LOOP_C_729, COMP_LOOP_C_730, COMP_LOOP_C_731,
      COMP_LOOP_C_732, COMP_LOOP_C_733, COMP_LOOP_C_734, COMP_LOOP_C_735, COMP_LOOP_C_736,
      COMP_LOOP_C_737, COMP_LOOP_C_738, COMP_LOOP_C_739, COMP_LOOP_C_740, COMP_LOOP_C_741,
      COMP_LOOP_C_742, COMP_LOOP_C_743, COMP_LOOP_C_744, COMP_LOOP_C_745, COMP_LOOP_C_746,
      COMP_LOOP_C_747, COMP_LOOP_C_748, COMP_LOOP_C_749, COMP_LOOP_C_750, COMP_LOOP_C_751,
      COMP_LOOP_C_752, COMP_LOOP_C_753, COMP_LOOP_C_754, COMP_LOOP_C_755, COMP_LOOP_C_756,
      COMP_LOOP_C_757, COMP_LOOP_C_758, COMP_LOOP_C_759, COMP_LOOP_C_760, COMP_LOOP_C_761,
      COMP_LOOP_C_762, COMP_LOOP_C_763, COMP_LOOP_C_764, COMP_LOOP_C_765, COMP_LOOP_C_766,
      COMP_LOOP_C_767, COMP_LOOP_C_768, COMP_LOOP_C_769, COMP_LOOP_13_modExp_1_while_C_0,
      COMP_LOOP_13_modExp_1_while_C_1, COMP_LOOP_13_modExp_1_while_C_2, COMP_LOOP_13_modExp_1_while_C_3,
      COMP_LOOP_13_modExp_1_while_C_4, COMP_LOOP_13_modExp_1_while_C_5, COMP_LOOP_13_modExp_1_while_C_6,
      COMP_LOOP_13_modExp_1_while_C_7, COMP_LOOP_13_modExp_1_while_C_8, COMP_LOOP_13_modExp_1_while_C_9,
      COMP_LOOP_13_modExp_1_while_C_10, COMP_LOOP_13_modExp_1_while_C_11, COMP_LOOP_13_modExp_1_while_C_12,
      COMP_LOOP_13_modExp_1_while_C_13, COMP_LOOP_13_modExp_1_while_C_14, COMP_LOOP_13_modExp_1_while_C_15,
      COMP_LOOP_13_modExp_1_while_C_16, COMP_LOOP_13_modExp_1_while_C_17, COMP_LOOP_13_modExp_1_while_C_18,
      COMP_LOOP_13_modExp_1_while_C_19, COMP_LOOP_13_modExp_1_while_C_20, COMP_LOOP_13_modExp_1_while_C_21,
      COMP_LOOP_13_modExp_1_while_C_22, COMP_LOOP_13_modExp_1_while_C_23, COMP_LOOP_13_modExp_1_while_C_24,
      COMP_LOOP_13_modExp_1_while_C_25, COMP_LOOP_13_modExp_1_while_C_26, COMP_LOOP_13_modExp_1_while_C_27,
      COMP_LOOP_13_modExp_1_while_C_28, COMP_LOOP_13_modExp_1_while_C_29, COMP_LOOP_13_modExp_1_while_C_30,
      COMP_LOOP_13_modExp_1_while_C_31, COMP_LOOP_13_modExp_1_while_C_32, COMP_LOOP_13_modExp_1_while_C_33,
      COMP_LOOP_13_modExp_1_while_C_34, COMP_LOOP_13_modExp_1_while_C_35, COMP_LOOP_13_modExp_1_while_C_36,
      COMP_LOOP_13_modExp_1_while_C_37, COMP_LOOP_13_modExp_1_while_C_38, COMP_LOOP_C_770,
      COMP_LOOP_C_771, COMP_LOOP_C_772, COMP_LOOP_C_773, COMP_LOOP_C_774, COMP_LOOP_C_775,
      COMP_LOOP_C_776, COMP_LOOP_C_777, COMP_LOOP_C_778, COMP_LOOP_C_779, COMP_LOOP_C_780,
      COMP_LOOP_C_781, COMP_LOOP_C_782, COMP_LOOP_C_783, COMP_LOOP_C_784, COMP_LOOP_C_785,
      COMP_LOOP_C_786, COMP_LOOP_C_787, COMP_LOOP_C_788, COMP_LOOP_C_789, COMP_LOOP_C_790,
      COMP_LOOP_C_791, COMP_LOOP_C_792, COMP_LOOP_C_793, COMP_LOOP_C_794, COMP_LOOP_C_795,
      COMP_LOOP_C_796, COMP_LOOP_C_797, COMP_LOOP_C_798, COMP_LOOP_C_799, COMP_LOOP_C_800,
      COMP_LOOP_C_801, COMP_LOOP_C_802, COMP_LOOP_C_803, COMP_LOOP_C_804, COMP_LOOP_C_805,
      COMP_LOOP_C_806, COMP_LOOP_C_807, COMP_LOOP_C_808, COMP_LOOP_C_809, COMP_LOOP_C_810,
      COMP_LOOP_C_811, COMP_LOOP_C_812, COMP_LOOP_C_813, COMP_LOOP_C_814, COMP_LOOP_C_815,
      COMP_LOOP_C_816, COMP_LOOP_C_817, COMP_LOOP_C_818, COMP_LOOP_C_819, COMP_LOOP_C_820,
      COMP_LOOP_C_821, COMP_LOOP_C_822, COMP_LOOP_C_823, COMP_LOOP_C_824, COMP_LOOP_C_825,
      COMP_LOOP_C_826, COMP_LOOP_C_827, COMP_LOOP_C_828, COMP_LOOP_C_829, COMP_LOOP_C_830,
      COMP_LOOP_C_831, COMP_LOOP_C_832, COMP_LOOP_C_833, COMP_LOOP_14_modExp_1_while_C_0,
      COMP_LOOP_14_modExp_1_while_C_1, COMP_LOOP_14_modExp_1_while_C_2, COMP_LOOP_14_modExp_1_while_C_3,
      COMP_LOOP_14_modExp_1_while_C_4, COMP_LOOP_14_modExp_1_while_C_5, COMP_LOOP_14_modExp_1_while_C_6,
      COMP_LOOP_14_modExp_1_while_C_7, COMP_LOOP_14_modExp_1_while_C_8, COMP_LOOP_14_modExp_1_while_C_9,
      COMP_LOOP_14_modExp_1_while_C_10, COMP_LOOP_14_modExp_1_while_C_11, COMP_LOOP_14_modExp_1_while_C_12,
      COMP_LOOP_14_modExp_1_while_C_13, COMP_LOOP_14_modExp_1_while_C_14, COMP_LOOP_14_modExp_1_while_C_15,
      COMP_LOOP_14_modExp_1_while_C_16, COMP_LOOP_14_modExp_1_while_C_17, COMP_LOOP_14_modExp_1_while_C_18,
      COMP_LOOP_14_modExp_1_while_C_19, COMP_LOOP_14_modExp_1_while_C_20, COMP_LOOP_14_modExp_1_while_C_21,
      COMP_LOOP_14_modExp_1_while_C_22, COMP_LOOP_14_modExp_1_while_C_23, COMP_LOOP_14_modExp_1_while_C_24,
      COMP_LOOP_14_modExp_1_while_C_25, COMP_LOOP_14_modExp_1_while_C_26, COMP_LOOP_14_modExp_1_while_C_27,
      COMP_LOOP_14_modExp_1_while_C_28, COMP_LOOP_14_modExp_1_while_C_29, COMP_LOOP_14_modExp_1_while_C_30,
      COMP_LOOP_14_modExp_1_while_C_31, COMP_LOOP_14_modExp_1_while_C_32, COMP_LOOP_14_modExp_1_while_C_33,
      COMP_LOOP_14_modExp_1_while_C_34, COMP_LOOP_14_modExp_1_while_C_35, COMP_LOOP_14_modExp_1_while_C_36,
      COMP_LOOP_14_modExp_1_while_C_37, COMP_LOOP_14_modExp_1_while_C_38, COMP_LOOP_C_834,
      COMP_LOOP_C_835, COMP_LOOP_C_836, COMP_LOOP_C_837, COMP_LOOP_C_838, COMP_LOOP_C_839,
      COMP_LOOP_C_840, COMP_LOOP_C_841, COMP_LOOP_C_842, COMP_LOOP_C_843, COMP_LOOP_C_844,
      COMP_LOOP_C_845, COMP_LOOP_C_846, COMP_LOOP_C_847, COMP_LOOP_C_848, COMP_LOOP_C_849,
      COMP_LOOP_C_850, COMP_LOOP_C_851, COMP_LOOP_C_852, COMP_LOOP_C_853, COMP_LOOP_C_854,
      COMP_LOOP_C_855, COMP_LOOP_C_856, COMP_LOOP_C_857, COMP_LOOP_C_858, COMP_LOOP_C_859,
      COMP_LOOP_C_860, COMP_LOOP_C_861, COMP_LOOP_C_862, COMP_LOOP_C_863, COMP_LOOP_C_864,
      COMP_LOOP_C_865, COMP_LOOP_C_866, COMP_LOOP_C_867, COMP_LOOP_C_868, COMP_LOOP_C_869,
      COMP_LOOP_C_870, COMP_LOOP_C_871, COMP_LOOP_C_872, COMP_LOOP_C_873, COMP_LOOP_C_874,
      COMP_LOOP_C_875, COMP_LOOP_C_876, COMP_LOOP_C_877, COMP_LOOP_C_878, COMP_LOOP_C_879,
      COMP_LOOP_C_880, COMP_LOOP_C_881, COMP_LOOP_C_882, COMP_LOOP_C_883, COMP_LOOP_C_884,
      COMP_LOOP_C_885, COMP_LOOP_C_886, COMP_LOOP_C_887, COMP_LOOP_C_888, COMP_LOOP_C_889,
      COMP_LOOP_C_890, COMP_LOOP_C_891, COMP_LOOP_C_892, COMP_LOOP_C_893, COMP_LOOP_C_894,
      COMP_LOOP_C_895, COMP_LOOP_C_896, COMP_LOOP_C_897, COMP_LOOP_15_modExp_1_while_C_0,
      COMP_LOOP_15_modExp_1_while_C_1, COMP_LOOP_15_modExp_1_while_C_2, COMP_LOOP_15_modExp_1_while_C_3,
      COMP_LOOP_15_modExp_1_while_C_4, COMP_LOOP_15_modExp_1_while_C_5, COMP_LOOP_15_modExp_1_while_C_6,
      COMP_LOOP_15_modExp_1_while_C_7, COMP_LOOP_15_modExp_1_while_C_8, COMP_LOOP_15_modExp_1_while_C_9,
      COMP_LOOP_15_modExp_1_while_C_10, COMP_LOOP_15_modExp_1_while_C_11, COMP_LOOP_15_modExp_1_while_C_12,
      COMP_LOOP_15_modExp_1_while_C_13, COMP_LOOP_15_modExp_1_while_C_14, COMP_LOOP_15_modExp_1_while_C_15,
      COMP_LOOP_15_modExp_1_while_C_16, COMP_LOOP_15_modExp_1_while_C_17, COMP_LOOP_15_modExp_1_while_C_18,
      COMP_LOOP_15_modExp_1_while_C_19, COMP_LOOP_15_modExp_1_while_C_20, COMP_LOOP_15_modExp_1_while_C_21,
      COMP_LOOP_15_modExp_1_while_C_22, COMP_LOOP_15_modExp_1_while_C_23, COMP_LOOP_15_modExp_1_while_C_24,
      COMP_LOOP_15_modExp_1_while_C_25, COMP_LOOP_15_modExp_1_while_C_26, COMP_LOOP_15_modExp_1_while_C_27,
      COMP_LOOP_15_modExp_1_while_C_28, COMP_LOOP_15_modExp_1_while_C_29, COMP_LOOP_15_modExp_1_while_C_30,
      COMP_LOOP_15_modExp_1_while_C_31, COMP_LOOP_15_modExp_1_while_C_32, COMP_LOOP_15_modExp_1_while_C_33,
      COMP_LOOP_15_modExp_1_while_C_34, COMP_LOOP_15_modExp_1_while_C_35, COMP_LOOP_15_modExp_1_while_C_36,
      COMP_LOOP_15_modExp_1_while_C_37, COMP_LOOP_15_modExp_1_while_C_38, COMP_LOOP_C_898,
      COMP_LOOP_C_899, COMP_LOOP_C_900, COMP_LOOP_C_901, COMP_LOOP_C_902, COMP_LOOP_C_903,
      COMP_LOOP_C_904, COMP_LOOP_C_905, COMP_LOOP_C_906, COMP_LOOP_C_907, COMP_LOOP_C_908,
      COMP_LOOP_C_909, COMP_LOOP_C_910, COMP_LOOP_C_911, COMP_LOOP_C_912, COMP_LOOP_C_913,
      COMP_LOOP_C_914, COMP_LOOP_C_915, COMP_LOOP_C_916, COMP_LOOP_C_917, COMP_LOOP_C_918,
      COMP_LOOP_C_919, COMP_LOOP_C_920, COMP_LOOP_C_921, COMP_LOOP_C_922, COMP_LOOP_C_923,
      COMP_LOOP_C_924, COMP_LOOP_C_925, COMP_LOOP_C_926, COMP_LOOP_C_927, COMP_LOOP_C_928,
      COMP_LOOP_C_929, COMP_LOOP_C_930, COMP_LOOP_C_931, COMP_LOOP_C_932, COMP_LOOP_C_933,
      COMP_LOOP_C_934, COMP_LOOP_C_935, COMP_LOOP_C_936, COMP_LOOP_C_937, COMP_LOOP_C_938,
      COMP_LOOP_C_939, COMP_LOOP_C_940, COMP_LOOP_C_941, COMP_LOOP_C_942, COMP_LOOP_C_943,
      COMP_LOOP_C_944, COMP_LOOP_C_945, COMP_LOOP_C_946, COMP_LOOP_C_947, COMP_LOOP_C_948,
      COMP_LOOP_C_949, COMP_LOOP_C_950, COMP_LOOP_C_951, COMP_LOOP_C_952, COMP_LOOP_C_953,
      COMP_LOOP_C_954, COMP_LOOP_C_955, COMP_LOOP_C_956, COMP_LOOP_C_957, COMP_LOOP_C_958,
      COMP_LOOP_C_959, COMP_LOOP_C_960, COMP_LOOP_C_961, COMP_LOOP_16_modExp_1_while_C_0,
      COMP_LOOP_16_modExp_1_while_C_1, COMP_LOOP_16_modExp_1_while_C_2, COMP_LOOP_16_modExp_1_while_C_3,
      COMP_LOOP_16_modExp_1_while_C_4, COMP_LOOP_16_modExp_1_while_C_5, COMP_LOOP_16_modExp_1_while_C_6,
      COMP_LOOP_16_modExp_1_while_C_7, COMP_LOOP_16_modExp_1_while_C_8, COMP_LOOP_16_modExp_1_while_C_9,
      COMP_LOOP_16_modExp_1_while_C_10, COMP_LOOP_16_modExp_1_while_C_11, COMP_LOOP_16_modExp_1_while_C_12,
      COMP_LOOP_16_modExp_1_while_C_13, COMP_LOOP_16_modExp_1_while_C_14, COMP_LOOP_16_modExp_1_while_C_15,
      COMP_LOOP_16_modExp_1_while_C_16, COMP_LOOP_16_modExp_1_while_C_17, COMP_LOOP_16_modExp_1_while_C_18,
      COMP_LOOP_16_modExp_1_while_C_19, COMP_LOOP_16_modExp_1_while_C_20, COMP_LOOP_16_modExp_1_while_C_21,
      COMP_LOOP_16_modExp_1_while_C_22, COMP_LOOP_16_modExp_1_while_C_23, COMP_LOOP_16_modExp_1_while_C_24,
      COMP_LOOP_16_modExp_1_while_C_25, COMP_LOOP_16_modExp_1_while_C_26, COMP_LOOP_16_modExp_1_while_C_27,
      COMP_LOOP_16_modExp_1_while_C_28, COMP_LOOP_16_modExp_1_while_C_29, COMP_LOOP_16_modExp_1_while_C_30,
      COMP_LOOP_16_modExp_1_while_C_31, COMP_LOOP_16_modExp_1_while_C_32, COMP_LOOP_16_modExp_1_while_C_33,
      COMP_LOOP_16_modExp_1_while_C_34, COMP_LOOP_16_modExp_1_while_C_35, COMP_LOOP_16_modExp_1_while_C_36,
      COMP_LOOP_16_modExp_1_while_C_37, COMP_LOOP_16_modExp_1_while_C_38, COMP_LOOP_C_962,
      COMP_LOOP_C_963, COMP_LOOP_C_964, COMP_LOOP_C_965, COMP_LOOP_C_966, COMP_LOOP_C_967,
      COMP_LOOP_C_968, COMP_LOOP_C_969, COMP_LOOP_C_970, COMP_LOOP_C_971, COMP_LOOP_C_972,
      COMP_LOOP_C_973, COMP_LOOP_C_974, COMP_LOOP_C_975, COMP_LOOP_C_976, COMP_LOOP_C_977,
      COMP_LOOP_C_978, COMP_LOOP_C_979, COMP_LOOP_C_980, COMP_LOOP_C_981, COMP_LOOP_C_982,
      COMP_LOOP_C_983, COMP_LOOP_C_984, COMP_LOOP_C_985, COMP_LOOP_C_986, COMP_LOOP_C_987,
      COMP_LOOP_C_988, COMP_LOOP_C_989, COMP_LOOP_C_990, COMP_LOOP_C_991, COMP_LOOP_C_992,
      COMP_LOOP_C_993, COMP_LOOP_C_994, COMP_LOOP_C_995, COMP_LOOP_C_996, COMP_LOOP_C_997,
      COMP_LOOP_C_998, COMP_LOOP_C_999, COMP_LOOP_C_1000, COMP_LOOP_C_1001, COMP_LOOP_C_1002,
      COMP_LOOP_C_1003, COMP_LOOP_C_1004, COMP_LOOP_C_1005, COMP_LOOP_C_1006, COMP_LOOP_C_1007,
      COMP_LOOP_C_1008, COMP_LOOP_C_1009, COMP_LOOP_C_1010, COMP_LOOP_C_1011, COMP_LOOP_C_1012,
      COMP_LOOP_C_1013, COMP_LOOP_C_1014, COMP_LOOP_C_1015, COMP_LOOP_C_1016, COMP_LOOP_C_1017,
      COMP_LOOP_C_1018, COMP_LOOP_C_1019, COMP_LOOP_C_1020, COMP_LOOP_C_1021, COMP_LOOP_C_1022,
      COMP_LOOP_C_1023, COMP_LOOP_C_1024, VEC_LOOP_C_0, STAGE_LOOP_C_9, main_C_1);

  SIGNAL state_var : inPlaceNTT_DIT_core_core_fsm_1_ST;
  SIGNAL state_var_NS : inPlaceNTT_DIT_core_core_fsm_1_ST;

BEGIN
  inPlaceNTT_DIT_core_core_fsm_1 : PROCESS (STAGE_LOOP_C_8_tr0, modExp_while_C_38_tr0,
      COMP_LOOP_C_1_tr0, COMP_LOOP_1_modExp_1_while_C_38_tr0, COMP_LOOP_C_64_tr0,
      COMP_LOOP_2_modExp_1_while_C_38_tr0, COMP_LOOP_C_128_tr0, COMP_LOOP_3_modExp_1_while_C_38_tr0,
      COMP_LOOP_C_192_tr0, COMP_LOOP_4_modExp_1_while_C_38_tr0, COMP_LOOP_C_256_tr0,
      COMP_LOOP_5_modExp_1_while_C_38_tr0, COMP_LOOP_C_320_tr0, COMP_LOOP_6_modExp_1_while_C_38_tr0,
      COMP_LOOP_C_384_tr0, COMP_LOOP_7_modExp_1_while_C_38_tr0, COMP_LOOP_C_448_tr0,
      COMP_LOOP_8_modExp_1_while_C_38_tr0, COMP_LOOP_C_512_tr0, COMP_LOOP_9_modExp_1_while_C_38_tr0,
      COMP_LOOP_C_576_tr0, COMP_LOOP_10_modExp_1_while_C_38_tr0, COMP_LOOP_C_640_tr0,
      COMP_LOOP_11_modExp_1_while_C_38_tr0, COMP_LOOP_C_704_tr0, COMP_LOOP_12_modExp_1_while_C_38_tr0,
      COMP_LOOP_C_768_tr0, COMP_LOOP_13_modExp_1_while_C_38_tr0, COMP_LOOP_C_832_tr0,
      COMP_LOOP_14_modExp_1_while_C_38_tr0, COMP_LOOP_C_896_tr0, COMP_LOOP_15_modExp_1_while_C_38_tr0,
      COMP_LOOP_C_960_tr0, COMP_LOOP_16_modExp_1_while_C_38_tr0, COMP_LOOP_C_1024_tr0,
      VEC_LOOP_C_0_tr0, STAGE_LOOP_C_9_tr0, state_var)
  BEGIN
    CASE state_var IS
      WHEN STAGE_LOOP_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000001");
        state_var_NS <= STAGE_LOOP_C_1;
      WHEN STAGE_LOOP_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000010");
        state_var_NS <= STAGE_LOOP_C_2;
      WHEN STAGE_LOOP_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000011");
        state_var_NS <= STAGE_LOOP_C_3;
      WHEN STAGE_LOOP_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000100");
        state_var_NS <= STAGE_LOOP_C_4;
      WHEN STAGE_LOOP_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000101");
        state_var_NS <= STAGE_LOOP_C_5;
      WHEN STAGE_LOOP_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000110");
        state_var_NS <= STAGE_LOOP_C_6;
      WHEN STAGE_LOOP_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000111");
        state_var_NS <= STAGE_LOOP_C_7;
      WHEN STAGE_LOOP_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000001000");
        state_var_NS <= STAGE_LOOP_C_8;
      WHEN STAGE_LOOP_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000001001");
        IF ( STAGE_LOOP_C_8_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_0;
        ELSE
          state_var_NS <= modExp_while_C_0;
        END IF;
      WHEN modExp_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000001010");
        state_var_NS <= modExp_while_C_1;
      WHEN modExp_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000001011");
        state_var_NS <= modExp_while_C_2;
      WHEN modExp_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000001100");
        state_var_NS <= modExp_while_C_3;
      WHEN modExp_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000001101");
        state_var_NS <= modExp_while_C_4;
      WHEN modExp_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000001110");
        state_var_NS <= modExp_while_C_5;
      WHEN modExp_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000001111");
        state_var_NS <= modExp_while_C_6;
      WHEN modExp_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000010000");
        state_var_NS <= modExp_while_C_7;
      WHEN modExp_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000010001");
        state_var_NS <= modExp_while_C_8;
      WHEN modExp_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000010010");
        state_var_NS <= modExp_while_C_9;
      WHEN modExp_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000010011");
        state_var_NS <= modExp_while_C_10;
      WHEN modExp_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000010100");
        state_var_NS <= modExp_while_C_11;
      WHEN modExp_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000010101");
        state_var_NS <= modExp_while_C_12;
      WHEN modExp_while_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000010110");
        state_var_NS <= modExp_while_C_13;
      WHEN modExp_while_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000010111");
        state_var_NS <= modExp_while_C_14;
      WHEN modExp_while_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000011000");
        state_var_NS <= modExp_while_C_15;
      WHEN modExp_while_C_15 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000011001");
        state_var_NS <= modExp_while_C_16;
      WHEN modExp_while_C_16 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000011010");
        state_var_NS <= modExp_while_C_17;
      WHEN modExp_while_C_17 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000011011");
        state_var_NS <= modExp_while_C_18;
      WHEN modExp_while_C_18 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000011100");
        state_var_NS <= modExp_while_C_19;
      WHEN modExp_while_C_19 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000011101");
        state_var_NS <= modExp_while_C_20;
      WHEN modExp_while_C_20 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000011110");
        state_var_NS <= modExp_while_C_21;
      WHEN modExp_while_C_21 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000011111");
        state_var_NS <= modExp_while_C_22;
      WHEN modExp_while_C_22 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000100000");
        state_var_NS <= modExp_while_C_23;
      WHEN modExp_while_C_23 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000100001");
        state_var_NS <= modExp_while_C_24;
      WHEN modExp_while_C_24 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000100010");
        state_var_NS <= modExp_while_C_25;
      WHEN modExp_while_C_25 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000100011");
        state_var_NS <= modExp_while_C_26;
      WHEN modExp_while_C_26 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000100100");
        state_var_NS <= modExp_while_C_27;
      WHEN modExp_while_C_27 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000100101");
        state_var_NS <= modExp_while_C_28;
      WHEN modExp_while_C_28 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000100110");
        state_var_NS <= modExp_while_C_29;
      WHEN modExp_while_C_29 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000100111");
        state_var_NS <= modExp_while_C_30;
      WHEN modExp_while_C_30 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000101000");
        state_var_NS <= modExp_while_C_31;
      WHEN modExp_while_C_31 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000101001");
        state_var_NS <= modExp_while_C_32;
      WHEN modExp_while_C_32 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000101010");
        state_var_NS <= modExp_while_C_33;
      WHEN modExp_while_C_33 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000101011");
        state_var_NS <= modExp_while_C_34;
      WHEN modExp_while_C_34 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000101100");
        state_var_NS <= modExp_while_C_35;
      WHEN modExp_while_C_35 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000101101");
        state_var_NS <= modExp_while_C_36;
      WHEN modExp_while_C_36 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000101110");
        state_var_NS <= modExp_while_C_37;
      WHEN modExp_while_C_37 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000101111");
        state_var_NS <= modExp_while_C_38;
      WHEN modExp_while_C_38 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000110000");
        IF ( modExp_while_C_38_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_0;
        ELSE
          state_var_NS <= modExp_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000110001");
        state_var_NS <= COMP_LOOP_C_1;
      WHEN COMP_LOOP_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000110010");
        IF ( COMP_LOOP_C_1_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_2;
        ELSE
          state_var_NS <= COMP_LOOP_1_modExp_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_1_modExp_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000110011");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_1;
      WHEN COMP_LOOP_1_modExp_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000110100");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_2;
      WHEN COMP_LOOP_1_modExp_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000110101");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_3;
      WHEN COMP_LOOP_1_modExp_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000110110");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_4;
      WHEN COMP_LOOP_1_modExp_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000110111");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_5;
      WHEN COMP_LOOP_1_modExp_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000111000");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_6;
      WHEN COMP_LOOP_1_modExp_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000111001");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_7;
      WHEN COMP_LOOP_1_modExp_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000111010");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_8;
      WHEN COMP_LOOP_1_modExp_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000111011");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_9;
      WHEN COMP_LOOP_1_modExp_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000111100");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_10;
      WHEN COMP_LOOP_1_modExp_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000111101");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_11;
      WHEN COMP_LOOP_1_modExp_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000111110");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_12;
      WHEN COMP_LOOP_1_modExp_1_while_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000111111");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_13;
      WHEN COMP_LOOP_1_modExp_1_while_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001000000");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_14;
      WHEN COMP_LOOP_1_modExp_1_while_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001000001");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_15;
      WHEN COMP_LOOP_1_modExp_1_while_C_15 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001000010");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_16;
      WHEN COMP_LOOP_1_modExp_1_while_C_16 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001000011");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_17;
      WHEN COMP_LOOP_1_modExp_1_while_C_17 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001000100");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_18;
      WHEN COMP_LOOP_1_modExp_1_while_C_18 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001000101");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_19;
      WHEN COMP_LOOP_1_modExp_1_while_C_19 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001000110");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_20;
      WHEN COMP_LOOP_1_modExp_1_while_C_20 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001000111");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_21;
      WHEN COMP_LOOP_1_modExp_1_while_C_21 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001001000");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_22;
      WHEN COMP_LOOP_1_modExp_1_while_C_22 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001001001");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_23;
      WHEN COMP_LOOP_1_modExp_1_while_C_23 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001001010");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_24;
      WHEN COMP_LOOP_1_modExp_1_while_C_24 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001001011");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_25;
      WHEN COMP_LOOP_1_modExp_1_while_C_25 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001001100");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_26;
      WHEN COMP_LOOP_1_modExp_1_while_C_26 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001001101");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_27;
      WHEN COMP_LOOP_1_modExp_1_while_C_27 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001001110");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_28;
      WHEN COMP_LOOP_1_modExp_1_while_C_28 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001001111");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_29;
      WHEN COMP_LOOP_1_modExp_1_while_C_29 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001010000");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_30;
      WHEN COMP_LOOP_1_modExp_1_while_C_30 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001010001");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_31;
      WHEN COMP_LOOP_1_modExp_1_while_C_31 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001010010");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_32;
      WHEN COMP_LOOP_1_modExp_1_while_C_32 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001010011");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_33;
      WHEN COMP_LOOP_1_modExp_1_while_C_33 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001010100");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_34;
      WHEN COMP_LOOP_1_modExp_1_while_C_34 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001010101");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_35;
      WHEN COMP_LOOP_1_modExp_1_while_C_35 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001010110");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_36;
      WHEN COMP_LOOP_1_modExp_1_while_C_36 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001010111");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_37;
      WHEN COMP_LOOP_1_modExp_1_while_C_37 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001011000");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_38;
      WHEN COMP_LOOP_1_modExp_1_while_C_38 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001011001");
        IF ( COMP_LOOP_1_modExp_1_while_C_38_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_2;
        ELSE
          state_var_NS <= COMP_LOOP_1_modExp_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001011010");
        state_var_NS <= COMP_LOOP_C_3;
      WHEN COMP_LOOP_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001011011");
        state_var_NS <= COMP_LOOP_C_4;
      WHEN COMP_LOOP_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001011100");
        state_var_NS <= COMP_LOOP_C_5;
      WHEN COMP_LOOP_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001011101");
        state_var_NS <= COMP_LOOP_C_6;
      WHEN COMP_LOOP_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001011110");
        state_var_NS <= COMP_LOOP_C_7;
      WHEN COMP_LOOP_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001011111");
        state_var_NS <= COMP_LOOP_C_8;
      WHEN COMP_LOOP_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001100000");
        state_var_NS <= COMP_LOOP_C_9;
      WHEN COMP_LOOP_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001100001");
        state_var_NS <= COMP_LOOP_C_10;
      WHEN COMP_LOOP_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001100010");
        state_var_NS <= COMP_LOOP_C_11;
      WHEN COMP_LOOP_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001100011");
        state_var_NS <= COMP_LOOP_C_12;
      WHEN COMP_LOOP_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001100100");
        state_var_NS <= COMP_LOOP_C_13;
      WHEN COMP_LOOP_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001100101");
        state_var_NS <= COMP_LOOP_C_14;
      WHEN COMP_LOOP_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001100110");
        state_var_NS <= COMP_LOOP_C_15;
      WHEN COMP_LOOP_C_15 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001100111");
        state_var_NS <= COMP_LOOP_C_16;
      WHEN COMP_LOOP_C_16 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001101000");
        state_var_NS <= COMP_LOOP_C_17;
      WHEN COMP_LOOP_C_17 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001101001");
        state_var_NS <= COMP_LOOP_C_18;
      WHEN COMP_LOOP_C_18 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001101010");
        state_var_NS <= COMP_LOOP_C_19;
      WHEN COMP_LOOP_C_19 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001101011");
        state_var_NS <= COMP_LOOP_C_20;
      WHEN COMP_LOOP_C_20 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001101100");
        state_var_NS <= COMP_LOOP_C_21;
      WHEN COMP_LOOP_C_21 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001101101");
        state_var_NS <= COMP_LOOP_C_22;
      WHEN COMP_LOOP_C_22 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001101110");
        state_var_NS <= COMP_LOOP_C_23;
      WHEN COMP_LOOP_C_23 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001101111");
        state_var_NS <= COMP_LOOP_C_24;
      WHEN COMP_LOOP_C_24 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001110000");
        state_var_NS <= COMP_LOOP_C_25;
      WHEN COMP_LOOP_C_25 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001110001");
        state_var_NS <= COMP_LOOP_C_26;
      WHEN COMP_LOOP_C_26 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001110010");
        state_var_NS <= COMP_LOOP_C_27;
      WHEN COMP_LOOP_C_27 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001110011");
        state_var_NS <= COMP_LOOP_C_28;
      WHEN COMP_LOOP_C_28 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001110100");
        state_var_NS <= COMP_LOOP_C_29;
      WHEN COMP_LOOP_C_29 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001110101");
        state_var_NS <= COMP_LOOP_C_30;
      WHEN COMP_LOOP_C_30 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001110110");
        state_var_NS <= COMP_LOOP_C_31;
      WHEN COMP_LOOP_C_31 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001110111");
        state_var_NS <= COMP_LOOP_C_32;
      WHEN COMP_LOOP_C_32 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001111000");
        state_var_NS <= COMP_LOOP_C_33;
      WHEN COMP_LOOP_C_33 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001111001");
        state_var_NS <= COMP_LOOP_C_34;
      WHEN COMP_LOOP_C_34 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001111010");
        state_var_NS <= COMP_LOOP_C_35;
      WHEN COMP_LOOP_C_35 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001111011");
        state_var_NS <= COMP_LOOP_C_36;
      WHEN COMP_LOOP_C_36 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001111100");
        state_var_NS <= COMP_LOOP_C_37;
      WHEN COMP_LOOP_C_37 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001111101");
        state_var_NS <= COMP_LOOP_C_38;
      WHEN COMP_LOOP_C_38 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001111110");
        state_var_NS <= COMP_LOOP_C_39;
      WHEN COMP_LOOP_C_39 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001111111");
        state_var_NS <= COMP_LOOP_C_40;
      WHEN COMP_LOOP_C_40 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010000000");
        state_var_NS <= COMP_LOOP_C_41;
      WHEN COMP_LOOP_C_41 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010000001");
        state_var_NS <= COMP_LOOP_C_42;
      WHEN COMP_LOOP_C_42 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010000010");
        state_var_NS <= COMP_LOOP_C_43;
      WHEN COMP_LOOP_C_43 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010000011");
        state_var_NS <= COMP_LOOP_C_44;
      WHEN COMP_LOOP_C_44 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010000100");
        state_var_NS <= COMP_LOOP_C_45;
      WHEN COMP_LOOP_C_45 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010000101");
        state_var_NS <= COMP_LOOP_C_46;
      WHEN COMP_LOOP_C_46 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010000110");
        state_var_NS <= COMP_LOOP_C_47;
      WHEN COMP_LOOP_C_47 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010000111");
        state_var_NS <= COMP_LOOP_C_48;
      WHEN COMP_LOOP_C_48 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010001000");
        state_var_NS <= COMP_LOOP_C_49;
      WHEN COMP_LOOP_C_49 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010001001");
        state_var_NS <= COMP_LOOP_C_50;
      WHEN COMP_LOOP_C_50 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010001010");
        state_var_NS <= COMP_LOOP_C_51;
      WHEN COMP_LOOP_C_51 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010001011");
        state_var_NS <= COMP_LOOP_C_52;
      WHEN COMP_LOOP_C_52 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010001100");
        state_var_NS <= COMP_LOOP_C_53;
      WHEN COMP_LOOP_C_53 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010001101");
        state_var_NS <= COMP_LOOP_C_54;
      WHEN COMP_LOOP_C_54 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010001110");
        state_var_NS <= COMP_LOOP_C_55;
      WHEN COMP_LOOP_C_55 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010001111");
        state_var_NS <= COMP_LOOP_C_56;
      WHEN COMP_LOOP_C_56 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010010000");
        state_var_NS <= COMP_LOOP_C_57;
      WHEN COMP_LOOP_C_57 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010010001");
        state_var_NS <= COMP_LOOP_C_58;
      WHEN COMP_LOOP_C_58 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010010010");
        state_var_NS <= COMP_LOOP_C_59;
      WHEN COMP_LOOP_C_59 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010010011");
        state_var_NS <= COMP_LOOP_C_60;
      WHEN COMP_LOOP_C_60 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010010100");
        state_var_NS <= COMP_LOOP_C_61;
      WHEN COMP_LOOP_C_61 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010010101");
        state_var_NS <= COMP_LOOP_C_62;
      WHEN COMP_LOOP_C_62 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010010110");
        state_var_NS <= COMP_LOOP_C_63;
      WHEN COMP_LOOP_C_63 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010010111");
        state_var_NS <= COMP_LOOP_C_64;
      WHEN COMP_LOOP_C_64 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010011000");
        IF ( COMP_LOOP_C_64_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_65;
        END IF;
      WHEN COMP_LOOP_C_65 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010011001");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_0;
      WHEN COMP_LOOP_2_modExp_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010011010");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_1;
      WHEN COMP_LOOP_2_modExp_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010011011");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_2;
      WHEN COMP_LOOP_2_modExp_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010011100");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_3;
      WHEN COMP_LOOP_2_modExp_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010011101");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_4;
      WHEN COMP_LOOP_2_modExp_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010011110");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_5;
      WHEN COMP_LOOP_2_modExp_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010011111");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_6;
      WHEN COMP_LOOP_2_modExp_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010100000");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_7;
      WHEN COMP_LOOP_2_modExp_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010100001");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_8;
      WHEN COMP_LOOP_2_modExp_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010100010");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_9;
      WHEN COMP_LOOP_2_modExp_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010100011");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_10;
      WHEN COMP_LOOP_2_modExp_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010100100");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_11;
      WHEN COMP_LOOP_2_modExp_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010100101");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_12;
      WHEN COMP_LOOP_2_modExp_1_while_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010100110");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_13;
      WHEN COMP_LOOP_2_modExp_1_while_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010100111");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_14;
      WHEN COMP_LOOP_2_modExp_1_while_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010101000");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_15;
      WHEN COMP_LOOP_2_modExp_1_while_C_15 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010101001");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_16;
      WHEN COMP_LOOP_2_modExp_1_while_C_16 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010101010");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_17;
      WHEN COMP_LOOP_2_modExp_1_while_C_17 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010101011");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_18;
      WHEN COMP_LOOP_2_modExp_1_while_C_18 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010101100");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_19;
      WHEN COMP_LOOP_2_modExp_1_while_C_19 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010101101");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_20;
      WHEN COMP_LOOP_2_modExp_1_while_C_20 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010101110");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_21;
      WHEN COMP_LOOP_2_modExp_1_while_C_21 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010101111");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_22;
      WHEN COMP_LOOP_2_modExp_1_while_C_22 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010110000");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_23;
      WHEN COMP_LOOP_2_modExp_1_while_C_23 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010110001");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_24;
      WHEN COMP_LOOP_2_modExp_1_while_C_24 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010110010");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_25;
      WHEN COMP_LOOP_2_modExp_1_while_C_25 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010110011");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_26;
      WHEN COMP_LOOP_2_modExp_1_while_C_26 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010110100");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_27;
      WHEN COMP_LOOP_2_modExp_1_while_C_27 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010110101");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_28;
      WHEN COMP_LOOP_2_modExp_1_while_C_28 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010110110");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_29;
      WHEN COMP_LOOP_2_modExp_1_while_C_29 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010110111");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_30;
      WHEN COMP_LOOP_2_modExp_1_while_C_30 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010111000");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_31;
      WHEN COMP_LOOP_2_modExp_1_while_C_31 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010111001");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_32;
      WHEN COMP_LOOP_2_modExp_1_while_C_32 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010111010");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_33;
      WHEN COMP_LOOP_2_modExp_1_while_C_33 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010111011");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_34;
      WHEN COMP_LOOP_2_modExp_1_while_C_34 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010111100");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_35;
      WHEN COMP_LOOP_2_modExp_1_while_C_35 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010111101");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_36;
      WHEN COMP_LOOP_2_modExp_1_while_C_36 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010111110");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_37;
      WHEN COMP_LOOP_2_modExp_1_while_C_37 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010111111");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_38;
      WHEN COMP_LOOP_2_modExp_1_while_C_38 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011000000");
        IF ( COMP_LOOP_2_modExp_1_while_C_38_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_66;
        ELSE
          state_var_NS <= COMP_LOOP_2_modExp_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_66 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011000001");
        state_var_NS <= COMP_LOOP_C_67;
      WHEN COMP_LOOP_C_67 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011000010");
        state_var_NS <= COMP_LOOP_C_68;
      WHEN COMP_LOOP_C_68 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011000011");
        state_var_NS <= COMP_LOOP_C_69;
      WHEN COMP_LOOP_C_69 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011000100");
        state_var_NS <= COMP_LOOP_C_70;
      WHEN COMP_LOOP_C_70 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011000101");
        state_var_NS <= COMP_LOOP_C_71;
      WHEN COMP_LOOP_C_71 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011000110");
        state_var_NS <= COMP_LOOP_C_72;
      WHEN COMP_LOOP_C_72 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011000111");
        state_var_NS <= COMP_LOOP_C_73;
      WHEN COMP_LOOP_C_73 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011001000");
        state_var_NS <= COMP_LOOP_C_74;
      WHEN COMP_LOOP_C_74 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011001001");
        state_var_NS <= COMP_LOOP_C_75;
      WHEN COMP_LOOP_C_75 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011001010");
        state_var_NS <= COMP_LOOP_C_76;
      WHEN COMP_LOOP_C_76 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011001011");
        state_var_NS <= COMP_LOOP_C_77;
      WHEN COMP_LOOP_C_77 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011001100");
        state_var_NS <= COMP_LOOP_C_78;
      WHEN COMP_LOOP_C_78 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011001101");
        state_var_NS <= COMP_LOOP_C_79;
      WHEN COMP_LOOP_C_79 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011001110");
        state_var_NS <= COMP_LOOP_C_80;
      WHEN COMP_LOOP_C_80 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011001111");
        state_var_NS <= COMP_LOOP_C_81;
      WHEN COMP_LOOP_C_81 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011010000");
        state_var_NS <= COMP_LOOP_C_82;
      WHEN COMP_LOOP_C_82 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011010001");
        state_var_NS <= COMP_LOOP_C_83;
      WHEN COMP_LOOP_C_83 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011010010");
        state_var_NS <= COMP_LOOP_C_84;
      WHEN COMP_LOOP_C_84 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011010011");
        state_var_NS <= COMP_LOOP_C_85;
      WHEN COMP_LOOP_C_85 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011010100");
        state_var_NS <= COMP_LOOP_C_86;
      WHEN COMP_LOOP_C_86 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011010101");
        state_var_NS <= COMP_LOOP_C_87;
      WHEN COMP_LOOP_C_87 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011010110");
        state_var_NS <= COMP_LOOP_C_88;
      WHEN COMP_LOOP_C_88 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011010111");
        state_var_NS <= COMP_LOOP_C_89;
      WHEN COMP_LOOP_C_89 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011011000");
        state_var_NS <= COMP_LOOP_C_90;
      WHEN COMP_LOOP_C_90 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011011001");
        state_var_NS <= COMP_LOOP_C_91;
      WHEN COMP_LOOP_C_91 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011011010");
        state_var_NS <= COMP_LOOP_C_92;
      WHEN COMP_LOOP_C_92 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011011011");
        state_var_NS <= COMP_LOOP_C_93;
      WHEN COMP_LOOP_C_93 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011011100");
        state_var_NS <= COMP_LOOP_C_94;
      WHEN COMP_LOOP_C_94 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011011101");
        state_var_NS <= COMP_LOOP_C_95;
      WHEN COMP_LOOP_C_95 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011011110");
        state_var_NS <= COMP_LOOP_C_96;
      WHEN COMP_LOOP_C_96 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011011111");
        state_var_NS <= COMP_LOOP_C_97;
      WHEN COMP_LOOP_C_97 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011100000");
        state_var_NS <= COMP_LOOP_C_98;
      WHEN COMP_LOOP_C_98 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011100001");
        state_var_NS <= COMP_LOOP_C_99;
      WHEN COMP_LOOP_C_99 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011100010");
        state_var_NS <= COMP_LOOP_C_100;
      WHEN COMP_LOOP_C_100 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011100011");
        state_var_NS <= COMP_LOOP_C_101;
      WHEN COMP_LOOP_C_101 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011100100");
        state_var_NS <= COMP_LOOP_C_102;
      WHEN COMP_LOOP_C_102 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011100101");
        state_var_NS <= COMP_LOOP_C_103;
      WHEN COMP_LOOP_C_103 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011100110");
        state_var_NS <= COMP_LOOP_C_104;
      WHEN COMP_LOOP_C_104 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011100111");
        state_var_NS <= COMP_LOOP_C_105;
      WHEN COMP_LOOP_C_105 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011101000");
        state_var_NS <= COMP_LOOP_C_106;
      WHEN COMP_LOOP_C_106 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011101001");
        state_var_NS <= COMP_LOOP_C_107;
      WHEN COMP_LOOP_C_107 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011101010");
        state_var_NS <= COMP_LOOP_C_108;
      WHEN COMP_LOOP_C_108 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011101011");
        state_var_NS <= COMP_LOOP_C_109;
      WHEN COMP_LOOP_C_109 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011101100");
        state_var_NS <= COMP_LOOP_C_110;
      WHEN COMP_LOOP_C_110 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011101101");
        state_var_NS <= COMP_LOOP_C_111;
      WHEN COMP_LOOP_C_111 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011101110");
        state_var_NS <= COMP_LOOP_C_112;
      WHEN COMP_LOOP_C_112 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011101111");
        state_var_NS <= COMP_LOOP_C_113;
      WHEN COMP_LOOP_C_113 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011110000");
        state_var_NS <= COMP_LOOP_C_114;
      WHEN COMP_LOOP_C_114 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011110001");
        state_var_NS <= COMP_LOOP_C_115;
      WHEN COMP_LOOP_C_115 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011110010");
        state_var_NS <= COMP_LOOP_C_116;
      WHEN COMP_LOOP_C_116 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011110011");
        state_var_NS <= COMP_LOOP_C_117;
      WHEN COMP_LOOP_C_117 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011110100");
        state_var_NS <= COMP_LOOP_C_118;
      WHEN COMP_LOOP_C_118 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011110101");
        state_var_NS <= COMP_LOOP_C_119;
      WHEN COMP_LOOP_C_119 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011110110");
        state_var_NS <= COMP_LOOP_C_120;
      WHEN COMP_LOOP_C_120 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011110111");
        state_var_NS <= COMP_LOOP_C_121;
      WHEN COMP_LOOP_C_121 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011111000");
        state_var_NS <= COMP_LOOP_C_122;
      WHEN COMP_LOOP_C_122 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011111001");
        state_var_NS <= COMP_LOOP_C_123;
      WHEN COMP_LOOP_C_123 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011111010");
        state_var_NS <= COMP_LOOP_C_124;
      WHEN COMP_LOOP_C_124 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011111011");
        state_var_NS <= COMP_LOOP_C_125;
      WHEN COMP_LOOP_C_125 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011111100");
        state_var_NS <= COMP_LOOP_C_126;
      WHEN COMP_LOOP_C_126 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011111101");
        state_var_NS <= COMP_LOOP_C_127;
      WHEN COMP_LOOP_C_127 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011111110");
        state_var_NS <= COMP_LOOP_C_128;
      WHEN COMP_LOOP_C_128 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011111111");
        IF ( COMP_LOOP_C_128_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_129;
        END IF;
      WHEN COMP_LOOP_C_129 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100000000");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_0;
      WHEN COMP_LOOP_3_modExp_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100000001");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_1;
      WHEN COMP_LOOP_3_modExp_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100000010");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_2;
      WHEN COMP_LOOP_3_modExp_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100000011");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_3;
      WHEN COMP_LOOP_3_modExp_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100000100");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_4;
      WHEN COMP_LOOP_3_modExp_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100000101");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_5;
      WHEN COMP_LOOP_3_modExp_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100000110");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_6;
      WHEN COMP_LOOP_3_modExp_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100000111");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_7;
      WHEN COMP_LOOP_3_modExp_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100001000");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_8;
      WHEN COMP_LOOP_3_modExp_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100001001");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_9;
      WHEN COMP_LOOP_3_modExp_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100001010");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_10;
      WHEN COMP_LOOP_3_modExp_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100001011");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_11;
      WHEN COMP_LOOP_3_modExp_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100001100");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_12;
      WHEN COMP_LOOP_3_modExp_1_while_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100001101");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_13;
      WHEN COMP_LOOP_3_modExp_1_while_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100001110");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_14;
      WHEN COMP_LOOP_3_modExp_1_while_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100001111");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_15;
      WHEN COMP_LOOP_3_modExp_1_while_C_15 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100010000");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_16;
      WHEN COMP_LOOP_3_modExp_1_while_C_16 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100010001");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_17;
      WHEN COMP_LOOP_3_modExp_1_while_C_17 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100010010");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_18;
      WHEN COMP_LOOP_3_modExp_1_while_C_18 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100010011");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_19;
      WHEN COMP_LOOP_3_modExp_1_while_C_19 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100010100");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_20;
      WHEN COMP_LOOP_3_modExp_1_while_C_20 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100010101");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_21;
      WHEN COMP_LOOP_3_modExp_1_while_C_21 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100010110");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_22;
      WHEN COMP_LOOP_3_modExp_1_while_C_22 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100010111");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_23;
      WHEN COMP_LOOP_3_modExp_1_while_C_23 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100011000");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_24;
      WHEN COMP_LOOP_3_modExp_1_while_C_24 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100011001");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_25;
      WHEN COMP_LOOP_3_modExp_1_while_C_25 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100011010");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_26;
      WHEN COMP_LOOP_3_modExp_1_while_C_26 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100011011");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_27;
      WHEN COMP_LOOP_3_modExp_1_while_C_27 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100011100");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_28;
      WHEN COMP_LOOP_3_modExp_1_while_C_28 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100011101");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_29;
      WHEN COMP_LOOP_3_modExp_1_while_C_29 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100011110");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_30;
      WHEN COMP_LOOP_3_modExp_1_while_C_30 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100011111");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_31;
      WHEN COMP_LOOP_3_modExp_1_while_C_31 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100100000");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_32;
      WHEN COMP_LOOP_3_modExp_1_while_C_32 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100100001");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_33;
      WHEN COMP_LOOP_3_modExp_1_while_C_33 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100100010");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_34;
      WHEN COMP_LOOP_3_modExp_1_while_C_34 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100100011");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_35;
      WHEN COMP_LOOP_3_modExp_1_while_C_35 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100100100");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_36;
      WHEN COMP_LOOP_3_modExp_1_while_C_36 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100100101");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_37;
      WHEN COMP_LOOP_3_modExp_1_while_C_37 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100100110");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_38;
      WHEN COMP_LOOP_3_modExp_1_while_C_38 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100100111");
        IF ( COMP_LOOP_3_modExp_1_while_C_38_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_130;
        ELSE
          state_var_NS <= COMP_LOOP_3_modExp_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_130 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100101000");
        state_var_NS <= COMP_LOOP_C_131;
      WHEN COMP_LOOP_C_131 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100101001");
        state_var_NS <= COMP_LOOP_C_132;
      WHEN COMP_LOOP_C_132 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100101010");
        state_var_NS <= COMP_LOOP_C_133;
      WHEN COMP_LOOP_C_133 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100101011");
        state_var_NS <= COMP_LOOP_C_134;
      WHEN COMP_LOOP_C_134 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100101100");
        state_var_NS <= COMP_LOOP_C_135;
      WHEN COMP_LOOP_C_135 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100101101");
        state_var_NS <= COMP_LOOP_C_136;
      WHEN COMP_LOOP_C_136 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100101110");
        state_var_NS <= COMP_LOOP_C_137;
      WHEN COMP_LOOP_C_137 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100101111");
        state_var_NS <= COMP_LOOP_C_138;
      WHEN COMP_LOOP_C_138 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100110000");
        state_var_NS <= COMP_LOOP_C_139;
      WHEN COMP_LOOP_C_139 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100110001");
        state_var_NS <= COMP_LOOP_C_140;
      WHEN COMP_LOOP_C_140 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100110010");
        state_var_NS <= COMP_LOOP_C_141;
      WHEN COMP_LOOP_C_141 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100110011");
        state_var_NS <= COMP_LOOP_C_142;
      WHEN COMP_LOOP_C_142 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100110100");
        state_var_NS <= COMP_LOOP_C_143;
      WHEN COMP_LOOP_C_143 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100110101");
        state_var_NS <= COMP_LOOP_C_144;
      WHEN COMP_LOOP_C_144 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100110110");
        state_var_NS <= COMP_LOOP_C_145;
      WHEN COMP_LOOP_C_145 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100110111");
        state_var_NS <= COMP_LOOP_C_146;
      WHEN COMP_LOOP_C_146 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100111000");
        state_var_NS <= COMP_LOOP_C_147;
      WHEN COMP_LOOP_C_147 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100111001");
        state_var_NS <= COMP_LOOP_C_148;
      WHEN COMP_LOOP_C_148 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100111010");
        state_var_NS <= COMP_LOOP_C_149;
      WHEN COMP_LOOP_C_149 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100111011");
        state_var_NS <= COMP_LOOP_C_150;
      WHEN COMP_LOOP_C_150 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100111100");
        state_var_NS <= COMP_LOOP_C_151;
      WHEN COMP_LOOP_C_151 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100111101");
        state_var_NS <= COMP_LOOP_C_152;
      WHEN COMP_LOOP_C_152 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100111110");
        state_var_NS <= COMP_LOOP_C_153;
      WHEN COMP_LOOP_C_153 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100111111");
        state_var_NS <= COMP_LOOP_C_154;
      WHEN COMP_LOOP_C_154 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101000000");
        state_var_NS <= COMP_LOOP_C_155;
      WHEN COMP_LOOP_C_155 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101000001");
        state_var_NS <= COMP_LOOP_C_156;
      WHEN COMP_LOOP_C_156 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101000010");
        state_var_NS <= COMP_LOOP_C_157;
      WHEN COMP_LOOP_C_157 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101000011");
        state_var_NS <= COMP_LOOP_C_158;
      WHEN COMP_LOOP_C_158 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101000100");
        state_var_NS <= COMP_LOOP_C_159;
      WHEN COMP_LOOP_C_159 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101000101");
        state_var_NS <= COMP_LOOP_C_160;
      WHEN COMP_LOOP_C_160 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101000110");
        state_var_NS <= COMP_LOOP_C_161;
      WHEN COMP_LOOP_C_161 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101000111");
        state_var_NS <= COMP_LOOP_C_162;
      WHEN COMP_LOOP_C_162 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101001000");
        state_var_NS <= COMP_LOOP_C_163;
      WHEN COMP_LOOP_C_163 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101001001");
        state_var_NS <= COMP_LOOP_C_164;
      WHEN COMP_LOOP_C_164 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101001010");
        state_var_NS <= COMP_LOOP_C_165;
      WHEN COMP_LOOP_C_165 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101001011");
        state_var_NS <= COMP_LOOP_C_166;
      WHEN COMP_LOOP_C_166 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101001100");
        state_var_NS <= COMP_LOOP_C_167;
      WHEN COMP_LOOP_C_167 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101001101");
        state_var_NS <= COMP_LOOP_C_168;
      WHEN COMP_LOOP_C_168 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101001110");
        state_var_NS <= COMP_LOOP_C_169;
      WHEN COMP_LOOP_C_169 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101001111");
        state_var_NS <= COMP_LOOP_C_170;
      WHEN COMP_LOOP_C_170 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101010000");
        state_var_NS <= COMP_LOOP_C_171;
      WHEN COMP_LOOP_C_171 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101010001");
        state_var_NS <= COMP_LOOP_C_172;
      WHEN COMP_LOOP_C_172 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101010010");
        state_var_NS <= COMP_LOOP_C_173;
      WHEN COMP_LOOP_C_173 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101010011");
        state_var_NS <= COMP_LOOP_C_174;
      WHEN COMP_LOOP_C_174 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101010100");
        state_var_NS <= COMP_LOOP_C_175;
      WHEN COMP_LOOP_C_175 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101010101");
        state_var_NS <= COMP_LOOP_C_176;
      WHEN COMP_LOOP_C_176 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101010110");
        state_var_NS <= COMP_LOOP_C_177;
      WHEN COMP_LOOP_C_177 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101010111");
        state_var_NS <= COMP_LOOP_C_178;
      WHEN COMP_LOOP_C_178 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101011000");
        state_var_NS <= COMP_LOOP_C_179;
      WHEN COMP_LOOP_C_179 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101011001");
        state_var_NS <= COMP_LOOP_C_180;
      WHEN COMP_LOOP_C_180 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101011010");
        state_var_NS <= COMP_LOOP_C_181;
      WHEN COMP_LOOP_C_181 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101011011");
        state_var_NS <= COMP_LOOP_C_182;
      WHEN COMP_LOOP_C_182 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101011100");
        state_var_NS <= COMP_LOOP_C_183;
      WHEN COMP_LOOP_C_183 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101011101");
        state_var_NS <= COMP_LOOP_C_184;
      WHEN COMP_LOOP_C_184 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101011110");
        state_var_NS <= COMP_LOOP_C_185;
      WHEN COMP_LOOP_C_185 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101011111");
        state_var_NS <= COMP_LOOP_C_186;
      WHEN COMP_LOOP_C_186 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101100000");
        state_var_NS <= COMP_LOOP_C_187;
      WHEN COMP_LOOP_C_187 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101100001");
        state_var_NS <= COMP_LOOP_C_188;
      WHEN COMP_LOOP_C_188 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101100010");
        state_var_NS <= COMP_LOOP_C_189;
      WHEN COMP_LOOP_C_189 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101100011");
        state_var_NS <= COMP_LOOP_C_190;
      WHEN COMP_LOOP_C_190 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101100100");
        state_var_NS <= COMP_LOOP_C_191;
      WHEN COMP_LOOP_C_191 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101100101");
        state_var_NS <= COMP_LOOP_C_192;
      WHEN COMP_LOOP_C_192 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101100110");
        IF ( COMP_LOOP_C_192_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_193;
        END IF;
      WHEN COMP_LOOP_C_193 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101100111");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_0;
      WHEN COMP_LOOP_4_modExp_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101101000");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_1;
      WHEN COMP_LOOP_4_modExp_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101101001");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_2;
      WHEN COMP_LOOP_4_modExp_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101101010");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_3;
      WHEN COMP_LOOP_4_modExp_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101101011");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_4;
      WHEN COMP_LOOP_4_modExp_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101101100");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_5;
      WHEN COMP_LOOP_4_modExp_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101101101");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_6;
      WHEN COMP_LOOP_4_modExp_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101101110");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_7;
      WHEN COMP_LOOP_4_modExp_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101101111");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_8;
      WHEN COMP_LOOP_4_modExp_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101110000");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_9;
      WHEN COMP_LOOP_4_modExp_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101110001");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_10;
      WHEN COMP_LOOP_4_modExp_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101110010");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_11;
      WHEN COMP_LOOP_4_modExp_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101110011");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_12;
      WHEN COMP_LOOP_4_modExp_1_while_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101110100");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_13;
      WHEN COMP_LOOP_4_modExp_1_while_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101110101");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_14;
      WHEN COMP_LOOP_4_modExp_1_while_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101110110");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_15;
      WHEN COMP_LOOP_4_modExp_1_while_C_15 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101110111");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_16;
      WHEN COMP_LOOP_4_modExp_1_while_C_16 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101111000");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_17;
      WHEN COMP_LOOP_4_modExp_1_while_C_17 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101111001");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_18;
      WHEN COMP_LOOP_4_modExp_1_while_C_18 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101111010");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_19;
      WHEN COMP_LOOP_4_modExp_1_while_C_19 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101111011");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_20;
      WHEN COMP_LOOP_4_modExp_1_while_C_20 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101111100");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_21;
      WHEN COMP_LOOP_4_modExp_1_while_C_21 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101111101");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_22;
      WHEN COMP_LOOP_4_modExp_1_while_C_22 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101111110");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_23;
      WHEN COMP_LOOP_4_modExp_1_while_C_23 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101111111");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_24;
      WHEN COMP_LOOP_4_modExp_1_while_C_24 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110000000");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_25;
      WHEN COMP_LOOP_4_modExp_1_while_C_25 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110000001");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_26;
      WHEN COMP_LOOP_4_modExp_1_while_C_26 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110000010");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_27;
      WHEN COMP_LOOP_4_modExp_1_while_C_27 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110000011");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_28;
      WHEN COMP_LOOP_4_modExp_1_while_C_28 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110000100");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_29;
      WHEN COMP_LOOP_4_modExp_1_while_C_29 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110000101");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_30;
      WHEN COMP_LOOP_4_modExp_1_while_C_30 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110000110");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_31;
      WHEN COMP_LOOP_4_modExp_1_while_C_31 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110000111");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_32;
      WHEN COMP_LOOP_4_modExp_1_while_C_32 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110001000");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_33;
      WHEN COMP_LOOP_4_modExp_1_while_C_33 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110001001");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_34;
      WHEN COMP_LOOP_4_modExp_1_while_C_34 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110001010");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_35;
      WHEN COMP_LOOP_4_modExp_1_while_C_35 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110001011");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_36;
      WHEN COMP_LOOP_4_modExp_1_while_C_36 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110001100");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_37;
      WHEN COMP_LOOP_4_modExp_1_while_C_37 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110001101");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_38;
      WHEN COMP_LOOP_4_modExp_1_while_C_38 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110001110");
        IF ( COMP_LOOP_4_modExp_1_while_C_38_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_194;
        ELSE
          state_var_NS <= COMP_LOOP_4_modExp_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_194 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110001111");
        state_var_NS <= COMP_LOOP_C_195;
      WHEN COMP_LOOP_C_195 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110010000");
        state_var_NS <= COMP_LOOP_C_196;
      WHEN COMP_LOOP_C_196 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110010001");
        state_var_NS <= COMP_LOOP_C_197;
      WHEN COMP_LOOP_C_197 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110010010");
        state_var_NS <= COMP_LOOP_C_198;
      WHEN COMP_LOOP_C_198 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110010011");
        state_var_NS <= COMP_LOOP_C_199;
      WHEN COMP_LOOP_C_199 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110010100");
        state_var_NS <= COMP_LOOP_C_200;
      WHEN COMP_LOOP_C_200 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110010101");
        state_var_NS <= COMP_LOOP_C_201;
      WHEN COMP_LOOP_C_201 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110010110");
        state_var_NS <= COMP_LOOP_C_202;
      WHEN COMP_LOOP_C_202 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110010111");
        state_var_NS <= COMP_LOOP_C_203;
      WHEN COMP_LOOP_C_203 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110011000");
        state_var_NS <= COMP_LOOP_C_204;
      WHEN COMP_LOOP_C_204 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110011001");
        state_var_NS <= COMP_LOOP_C_205;
      WHEN COMP_LOOP_C_205 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110011010");
        state_var_NS <= COMP_LOOP_C_206;
      WHEN COMP_LOOP_C_206 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110011011");
        state_var_NS <= COMP_LOOP_C_207;
      WHEN COMP_LOOP_C_207 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110011100");
        state_var_NS <= COMP_LOOP_C_208;
      WHEN COMP_LOOP_C_208 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110011101");
        state_var_NS <= COMP_LOOP_C_209;
      WHEN COMP_LOOP_C_209 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110011110");
        state_var_NS <= COMP_LOOP_C_210;
      WHEN COMP_LOOP_C_210 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110011111");
        state_var_NS <= COMP_LOOP_C_211;
      WHEN COMP_LOOP_C_211 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110100000");
        state_var_NS <= COMP_LOOP_C_212;
      WHEN COMP_LOOP_C_212 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110100001");
        state_var_NS <= COMP_LOOP_C_213;
      WHEN COMP_LOOP_C_213 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110100010");
        state_var_NS <= COMP_LOOP_C_214;
      WHEN COMP_LOOP_C_214 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110100011");
        state_var_NS <= COMP_LOOP_C_215;
      WHEN COMP_LOOP_C_215 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110100100");
        state_var_NS <= COMP_LOOP_C_216;
      WHEN COMP_LOOP_C_216 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110100101");
        state_var_NS <= COMP_LOOP_C_217;
      WHEN COMP_LOOP_C_217 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110100110");
        state_var_NS <= COMP_LOOP_C_218;
      WHEN COMP_LOOP_C_218 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110100111");
        state_var_NS <= COMP_LOOP_C_219;
      WHEN COMP_LOOP_C_219 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110101000");
        state_var_NS <= COMP_LOOP_C_220;
      WHEN COMP_LOOP_C_220 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110101001");
        state_var_NS <= COMP_LOOP_C_221;
      WHEN COMP_LOOP_C_221 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110101010");
        state_var_NS <= COMP_LOOP_C_222;
      WHEN COMP_LOOP_C_222 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110101011");
        state_var_NS <= COMP_LOOP_C_223;
      WHEN COMP_LOOP_C_223 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110101100");
        state_var_NS <= COMP_LOOP_C_224;
      WHEN COMP_LOOP_C_224 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110101101");
        state_var_NS <= COMP_LOOP_C_225;
      WHEN COMP_LOOP_C_225 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110101110");
        state_var_NS <= COMP_LOOP_C_226;
      WHEN COMP_LOOP_C_226 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110101111");
        state_var_NS <= COMP_LOOP_C_227;
      WHEN COMP_LOOP_C_227 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110110000");
        state_var_NS <= COMP_LOOP_C_228;
      WHEN COMP_LOOP_C_228 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110110001");
        state_var_NS <= COMP_LOOP_C_229;
      WHEN COMP_LOOP_C_229 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110110010");
        state_var_NS <= COMP_LOOP_C_230;
      WHEN COMP_LOOP_C_230 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110110011");
        state_var_NS <= COMP_LOOP_C_231;
      WHEN COMP_LOOP_C_231 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110110100");
        state_var_NS <= COMP_LOOP_C_232;
      WHEN COMP_LOOP_C_232 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110110101");
        state_var_NS <= COMP_LOOP_C_233;
      WHEN COMP_LOOP_C_233 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110110110");
        state_var_NS <= COMP_LOOP_C_234;
      WHEN COMP_LOOP_C_234 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110110111");
        state_var_NS <= COMP_LOOP_C_235;
      WHEN COMP_LOOP_C_235 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110111000");
        state_var_NS <= COMP_LOOP_C_236;
      WHEN COMP_LOOP_C_236 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110111001");
        state_var_NS <= COMP_LOOP_C_237;
      WHEN COMP_LOOP_C_237 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110111010");
        state_var_NS <= COMP_LOOP_C_238;
      WHEN COMP_LOOP_C_238 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110111011");
        state_var_NS <= COMP_LOOP_C_239;
      WHEN COMP_LOOP_C_239 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110111100");
        state_var_NS <= COMP_LOOP_C_240;
      WHEN COMP_LOOP_C_240 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110111101");
        state_var_NS <= COMP_LOOP_C_241;
      WHEN COMP_LOOP_C_241 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110111110");
        state_var_NS <= COMP_LOOP_C_242;
      WHEN COMP_LOOP_C_242 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110111111");
        state_var_NS <= COMP_LOOP_C_243;
      WHEN COMP_LOOP_C_243 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111000000");
        state_var_NS <= COMP_LOOP_C_244;
      WHEN COMP_LOOP_C_244 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111000001");
        state_var_NS <= COMP_LOOP_C_245;
      WHEN COMP_LOOP_C_245 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111000010");
        state_var_NS <= COMP_LOOP_C_246;
      WHEN COMP_LOOP_C_246 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111000011");
        state_var_NS <= COMP_LOOP_C_247;
      WHEN COMP_LOOP_C_247 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111000100");
        state_var_NS <= COMP_LOOP_C_248;
      WHEN COMP_LOOP_C_248 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111000101");
        state_var_NS <= COMP_LOOP_C_249;
      WHEN COMP_LOOP_C_249 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111000110");
        state_var_NS <= COMP_LOOP_C_250;
      WHEN COMP_LOOP_C_250 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111000111");
        state_var_NS <= COMP_LOOP_C_251;
      WHEN COMP_LOOP_C_251 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111001000");
        state_var_NS <= COMP_LOOP_C_252;
      WHEN COMP_LOOP_C_252 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111001001");
        state_var_NS <= COMP_LOOP_C_253;
      WHEN COMP_LOOP_C_253 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111001010");
        state_var_NS <= COMP_LOOP_C_254;
      WHEN COMP_LOOP_C_254 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111001011");
        state_var_NS <= COMP_LOOP_C_255;
      WHEN COMP_LOOP_C_255 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111001100");
        state_var_NS <= COMP_LOOP_C_256;
      WHEN COMP_LOOP_C_256 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111001101");
        IF ( COMP_LOOP_C_256_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_257;
        END IF;
      WHEN COMP_LOOP_C_257 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111001110");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_0;
      WHEN COMP_LOOP_5_modExp_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111001111");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_1;
      WHEN COMP_LOOP_5_modExp_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111010000");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_2;
      WHEN COMP_LOOP_5_modExp_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111010001");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_3;
      WHEN COMP_LOOP_5_modExp_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111010010");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_4;
      WHEN COMP_LOOP_5_modExp_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111010011");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_5;
      WHEN COMP_LOOP_5_modExp_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111010100");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_6;
      WHEN COMP_LOOP_5_modExp_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111010101");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_7;
      WHEN COMP_LOOP_5_modExp_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111010110");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_8;
      WHEN COMP_LOOP_5_modExp_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111010111");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_9;
      WHEN COMP_LOOP_5_modExp_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111011000");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_10;
      WHEN COMP_LOOP_5_modExp_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111011001");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_11;
      WHEN COMP_LOOP_5_modExp_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111011010");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_12;
      WHEN COMP_LOOP_5_modExp_1_while_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111011011");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_13;
      WHEN COMP_LOOP_5_modExp_1_while_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111011100");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_14;
      WHEN COMP_LOOP_5_modExp_1_while_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111011101");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_15;
      WHEN COMP_LOOP_5_modExp_1_while_C_15 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111011110");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_16;
      WHEN COMP_LOOP_5_modExp_1_while_C_16 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111011111");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_17;
      WHEN COMP_LOOP_5_modExp_1_while_C_17 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111100000");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_18;
      WHEN COMP_LOOP_5_modExp_1_while_C_18 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111100001");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_19;
      WHEN COMP_LOOP_5_modExp_1_while_C_19 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111100010");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_20;
      WHEN COMP_LOOP_5_modExp_1_while_C_20 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111100011");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_21;
      WHEN COMP_LOOP_5_modExp_1_while_C_21 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111100100");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_22;
      WHEN COMP_LOOP_5_modExp_1_while_C_22 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111100101");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_23;
      WHEN COMP_LOOP_5_modExp_1_while_C_23 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111100110");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_24;
      WHEN COMP_LOOP_5_modExp_1_while_C_24 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111100111");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_25;
      WHEN COMP_LOOP_5_modExp_1_while_C_25 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111101000");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_26;
      WHEN COMP_LOOP_5_modExp_1_while_C_26 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111101001");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_27;
      WHEN COMP_LOOP_5_modExp_1_while_C_27 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111101010");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_28;
      WHEN COMP_LOOP_5_modExp_1_while_C_28 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111101011");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_29;
      WHEN COMP_LOOP_5_modExp_1_while_C_29 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111101100");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_30;
      WHEN COMP_LOOP_5_modExp_1_while_C_30 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111101101");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_31;
      WHEN COMP_LOOP_5_modExp_1_while_C_31 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111101110");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_32;
      WHEN COMP_LOOP_5_modExp_1_while_C_32 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111101111");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_33;
      WHEN COMP_LOOP_5_modExp_1_while_C_33 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111110000");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_34;
      WHEN COMP_LOOP_5_modExp_1_while_C_34 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111110001");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_35;
      WHEN COMP_LOOP_5_modExp_1_while_C_35 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111110010");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_36;
      WHEN COMP_LOOP_5_modExp_1_while_C_36 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111110011");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_37;
      WHEN COMP_LOOP_5_modExp_1_while_C_37 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111110100");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_38;
      WHEN COMP_LOOP_5_modExp_1_while_C_38 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111110101");
        IF ( COMP_LOOP_5_modExp_1_while_C_38_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_258;
        ELSE
          state_var_NS <= COMP_LOOP_5_modExp_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_258 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111110110");
        state_var_NS <= COMP_LOOP_C_259;
      WHEN COMP_LOOP_C_259 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111110111");
        state_var_NS <= COMP_LOOP_C_260;
      WHEN COMP_LOOP_C_260 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111111000");
        state_var_NS <= COMP_LOOP_C_261;
      WHEN COMP_LOOP_C_261 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111111001");
        state_var_NS <= COMP_LOOP_C_262;
      WHEN COMP_LOOP_C_262 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111111010");
        state_var_NS <= COMP_LOOP_C_263;
      WHEN COMP_LOOP_C_263 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111111011");
        state_var_NS <= COMP_LOOP_C_264;
      WHEN COMP_LOOP_C_264 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111111100");
        state_var_NS <= COMP_LOOP_C_265;
      WHEN COMP_LOOP_C_265 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111111101");
        state_var_NS <= COMP_LOOP_C_266;
      WHEN COMP_LOOP_C_266 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111111110");
        state_var_NS <= COMP_LOOP_C_267;
      WHEN COMP_LOOP_C_267 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111111111");
        state_var_NS <= COMP_LOOP_C_268;
      WHEN COMP_LOOP_C_268 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000000000");
        state_var_NS <= COMP_LOOP_C_269;
      WHEN COMP_LOOP_C_269 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000000001");
        state_var_NS <= COMP_LOOP_C_270;
      WHEN COMP_LOOP_C_270 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000000010");
        state_var_NS <= COMP_LOOP_C_271;
      WHEN COMP_LOOP_C_271 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000000011");
        state_var_NS <= COMP_LOOP_C_272;
      WHEN COMP_LOOP_C_272 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000000100");
        state_var_NS <= COMP_LOOP_C_273;
      WHEN COMP_LOOP_C_273 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000000101");
        state_var_NS <= COMP_LOOP_C_274;
      WHEN COMP_LOOP_C_274 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000000110");
        state_var_NS <= COMP_LOOP_C_275;
      WHEN COMP_LOOP_C_275 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000000111");
        state_var_NS <= COMP_LOOP_C_276;
      WHEN COMP_LOOP_C_276 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000001000");
        state_var_NS <= COMP_LOOP_C_277;
      WHEN COMP_LOOP_C_277 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000001001");
        state_var_NS <= COMP_LOOP_C_278;
      WHEN COMP_LOOP_C_278 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000001010");
        state_var_NS <= COMP_LOOP_C_279;
      WHEN COMP_LOOP_C_279 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000001011");
        state_var_NS <= COMP_LOOP_C_280;
      WHEN COMP_LOOP_C_280 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000001100");
        state_var_NS <= COMP_LOOP_C_281;
      WHEN COMP_LOOP_C_281 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000001101");
        state_var_NS <= COMP_LOOP_C_282;
      WHEN COMP_LOOP_C_282 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000001110");
        state_var_NS <= COMP_LOOP_C_283;
      WHEN COMP_LOOP_C_283 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000001111");
        state_var_NS <= COMP_LOOP_C_284;
      WHEN COMP_LOOP_C_284 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000010000");
        state_var_NS <= COMP_LOOP_C_285;
      WHEN COMP_LOOP_C_285 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000010001");
        state_var_NS <= COMP_LOOP_C_286;
      WHEN COMP_LOOP_C_286 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000010010");
        state_var_NS <= COMP_LOOP_C_287;
      WHEN COMP_LOOP_C_287 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000010011");
        state_var_NS <= COMP_LOOP_C_288;
      WHEN COMP_LOOP_C_288 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000010100");
        state_var_NS <= COMP_LOOP_C_289;
      WHEN COMP_LOOP_C_289 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000010101");
        state_var_NS <= COMP_LOOP_C_290;
      WHEN COMP_LOOP_C_290 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000010110");
        state_var_NS <= COMP_LOOP_C_291;
      WHEN COMP_LOOP_C_291 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000010111");
        state_var_NS <= COMP_LOOP_C_292;
      WHEN COMP_LOOP_C_292 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000011000");
        state_var_NS <= COMP_LOOP_C_293;
      WHEN COMP_LOOP_C_293 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000011001");
        state_var_NS <= COMP_LOOP_C_294;
      WHEN COMP_LOOP_C_294 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000011010");
        state_var_NS <= COMP_LOOP_C_295;
      WHEN COMP_LOOP_C_295 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000011011");
        state_var_NS <= COMP_LOOP_C_296;
      WHEN COMP_LOOP_C_296 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000011100");
        state_var_NS <= COMP_LOOP_C_297;
      WHEN COMP_LOOP_C_297 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000011101");
        state_var_NS <= COMP_LOOP_C_298;
      WHEN COMP_LOOP_C_298 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000011110");
        state_var_NS <= COMP_LOOP_C_299;
      WHEN COMP_LOOP_C_299 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000011111");
        state_var_NS <= COMP_LOOP_C_300;
      WHEN COMP_LOOP_C_300 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000100000");
        state_var_NS <= COMP_LOOP_C_301;
      WHEN COMP_LOOP_C_301 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000100001");
        state_var_NS <= COMP_LOOP_C_302;
      WHEN COMP_LOOP_C_302 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000100010");
        state_var_NS <= COMP_LOOP_C_303;
      WHEN COMP_LOOP_C_303 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000100011");
        state_var_NS <= COMP_LOOP_C_304;
      WHEN COMP_LOOP_C_304 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000100100");
        state_var_NS <= COMP_LOOP_C_305;
      WHEN COMP_LOOP_C_305 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000100101");
        state_var_NS <= COMP_LOOP_C_306;
      WHEN COMP_LOOP_C_306 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000100110");
        state_var_NS <= COMP_LOOP_C_307;
      WHEN COMP_LOOP_C_307 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000100111");
        state_var_NS <= COMP_LOOP_C_308;
      WHEN COMP_LOOP_C_308 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000101000");
        state_var_NS <= COMP_LOOP_C_309;
      WHEN COMP_LOOP_C_309 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000101001");
        state_var_NS <= COMP_LOOP_C_310;
      WHEN COMP_LOOP_C_310 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000101010");
        state_var_NS <= COMP_LOOP_C_311;
      WHEN COMP_LOOP_C_311 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000101011");
        state_var_NS <= COMP_LOOP_C_312;
      WHEN COMP_LOOP_C_312 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000101100");
        state_var_NS <= COMP_LOOP_C_313;
      WHEN COMP_LOOP_C_313 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000101101");
        state_var_NS <= COMP_LOOP_C_314;
      WHEN COMP_LOOP_C_314 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000101110");
        state_var_NS <= COMP_LOOP_C_315;
      WHEN COMP_LOOP_C_315 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000101111");
        state_var_NS <= COMP_LOOP_C_316;
      WHEN COMP_LOOP_C_316 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000110000");
        state_var_NS <= COMP_LOOP_C_317;
      WHEN COMP_LOOP_C_317 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000110001");
        state_var_NS <= COMP_LOOP_C_318;
      WHEN COMP_LOOP_C_318 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000110010");
        state_var_NS <= COMP_LOOP_C_319;
      WHEN COMP_LOOP_C_319 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000110011");
        state_var_NS <= COMP_LOOP_C_320;
      WHEN COMP_LOOP_C_320 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000110100");
        IF ( COMP_LOOP_C_320_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_321;
        END IF;
      WHEN COMP_LOOP_C_321 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000110101");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_0;
      WHEN COMP_LOOP_6_modExp_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000110110");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_1;
      WHEN COMP_LOOP_6_modExp_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000110111");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_2;
      WHEN COMP_LOOP_6_modExp_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000111000");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_3;
      WHEN COMP_LOOP_6_modExp_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000111001");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_4;
      WHEN COMP_LOOP_6_modExp_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000111010");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_5;
      WHEN COMP_LOOP_6_modExp_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000111011");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_6;
      WHEN COMP_LOOP_6_modExp_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000111100");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_7;
      WHEN COMP_LOOP_6_modExp_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000111101");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_8;
      WHEN COMP_LOOP_6_modExp_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000111110");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_9;
      WHEN COMP_LOOP_6_modExp_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000111111");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_10;
      WHEN COMP_LOOP_6_modExp_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001000000");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_11;
      WHEN COMP_LOOP_6_modExp_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001000001");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_12;
      WHEN COMP_LOOP_6_modExp_1_while_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001000010");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_13;
      WHEN COMP_LOOP_6_modExp_1_while_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001000011");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_14;
      WHEN COMP_LOOP_6_modExp_1_while_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001000100");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_15;
      WHEN COMP_LOOP_6_modExp_1_while_C_15 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001000101");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_16;
      WHEN COMP_LOOP_6_modExp_1_while_C_16 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001000110");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_17;
      WHEN COMP_LOOP_6_modExp_1_while_C_17 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001000111");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_18;
      WHEN COMP_LOOP_6_modExp_1_while_C_18 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001001000");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_19;
      WHEN COMP_LOOP_6_modExp_1_while_C_19 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001001001");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_20;
      WHEN COMP_LOOP_6_modExp_1_while_C_20 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001001010");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_21;
      WHEN COMP_LOOP_6_modExp_1_while_C_21 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001001011");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_22;
      WHEN COMP_LOOP_6_modExp_1_while_C_22 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001001100");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_23;
      WHEN COMP_LOOP_6_modExp_1_while_C_23 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001001101");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_24;
      WHEN COMP_LOOP_6_modExp_1_while_C_24 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001001110");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_25;
      WHEN COMP_LOOP_6_modExp_1_while_C_25 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001001111");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_26;
      WHEN COMP_LOOP_6_modExp_1_while_C_26 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001010000");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_27;
      WHEN COMP_LOOP_6_modExp_1_while_C_27 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001010001");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_28;
      WHEN COMP_LOOP_6_modExp_1_while_C_28 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001010010");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_29;
      WHEN COMP_LOOP_6_modExp_1_while_C_29 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001010011");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_30;
      WHEN COMP_LOOP_6_modExp_1_while_C_30 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001010100");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_31;
      WHEN COMP_LOOP_6_modExp_1_while_C_31 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001010101");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_32;
      WHEN COMP_LOOP_6_modExp_1_while_C_32 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001010110");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_33;
      WHEN COMP_LOOP_6_modExp_1_while_C_33 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001010111");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_34;
      WHEN COMP_LOOP_6_modExp_1_while_C_34 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001011000");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_35;
      WHEN COMP_LOOP_6_modExp_1_while_C_35 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001011001");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_36;
      WHEN COMP_LOOP_6_modExp_1_while_C_36 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001011010");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_37;
      WHEN COMP_LOOP_6_modExp_1_while_C_37 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001011011");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_38;
      WHEN COMP_LOOP_6_modExp_1_while_C_38 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001011100");
        IF ( COMP_LOOP_6_modExp_1_while_C_38_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_322;
        ELSE
          state_var_NS <= COMP_LOOP_6_modExp_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_322 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001011101");
        state_var_NS <= COMP_LOOP_C_323;
      WHEN COMP_LOOP_C_323 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001011110");
        state_var_NS <= COMP_LOOP_C_324;
      WHEN COMP_LOOP_C_324 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001011111");
        state_var_NS <= COMP_LOOP_C_325;
      WHEN COMP_LOOP_C_325 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001100000");
        state_var_NS <= COMP_LOOP_C_326;
      WHEN COMP_LOOP_C_326 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001100001");
        state_var_NS <= COMP_LOOP_C_327;
      WHEN COMP_LOOP_C_327 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001100010");
        state_var_NS <= COMP_LOOP_C_328;
      WHEN COMP_LOOP_C_328 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001100011");
        state_var_NS <= COMP_LOOP_C_329;
      WHEN COMP_LOOP_C_329 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001100100");
        state_var_NS <= COMP_LOOP_C_330;
      WHEN COMP_LOOP_C_330 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001100101");
        state_var_NS <= COMP_LOOP_C_331;
      WHEN COMP_LOOP_C_331 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001100110");
        state_var_NS <= COMP_LOOP_C_332;
      WHEN COMP_LOOP_C_332 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001100111");
        state_var_NS <= COMP_LOOP_C_333;
      WHEN COMP_LOOP_C_333 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001101000");
        state_var_NS <= COMP_LOOP_C_334;
      WHEN COMP_LOOP_C_334 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001101001");
        state_var_NS <= COMP_LOOP_C_335;
      WHEN COMP_LOOP_C_335 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001101010");
        state_var_NS <= COMP_LOOP_C_336;
      WHEN COMP_LOOP_C_336 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001101011");
        state_var_NS <= COMP_LOOP_C_337;
      WHEN COMP_LOOP_C_337 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001101100");
        state_var_NS <= COMP_LOOP_C_338;
      WHEN COMP_LOOP_C_338 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001101101");
        state_var_NS <= COMP_LOOP_C_339;
      WHEN COMP_LOOP_C_339 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001101110");
        state_var_NS <= COMP_LOOP_C_340;
      WHEN COMP_LOOP_C_340 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001101111");
        state_var_NS <= COMP_LOOP_C_341;
      WHEN COMP_LOOP_C_341 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001110000");
        state_var_NS <= COMP_LOOP_C_342;
      WHEN COMP_LOOP_C_342 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001110001");
        state_var_NS <= COMP_LOOP_C_343;
      WHEN COMP_LOOP_C_343 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001110010");
        state_var_NS <= COMP_LOOP_C_344;
      WHEN COMP_LOOP_C_344 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001110011");
        state_var_NS <= COMP_LOOP_C_345;
      WHEN COMP_LOOP_C_345 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001110100");
        state_var_NS <= COMP_LOOP_C_346;
      WHEN COMP_LOOP_C_346 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001110101");
        state_var_NS <= COMP_LOOP_C_347;
      WHEN COMP_LOOP_C_347 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001110110");
        state_var_NS <= COMP_LOOP_C_348;
      WHEN COMP_LOOP_C_348 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001110111");
        state_var_NS <= COMP_LOOP_C_349;
      WHEN COMP_LOOP_C_349 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001111000");
        state_var_NS <= COMP_LOOP_C_350;
      WHEN COMP_LOOP_C_350 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001111001");
        state_var_NS <= COMP_LOOP_C_351;
      WHEN COMP_LOOP_C_351 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001111010");
        state_var_NS <= COMP_LOOP_C_352;
      WHEN COMP_LOOP_C_352 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001111011");
        state_var_NS <= COMP_LOOP_C_353;
      WHEN COMP_LOOP_C_353 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001111100");
        state_var_NS <= COMP_LOOP_C_354;
      WHEN COMP_LOOP_C_354 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001111101");
        state_var_NS <= COMP_LOOP_C_355;
      WHEN COMP_LOOP_C_355 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001111110");
        state_var_NS <= COMP_LOOP_C_356;
      WHEN COMP_LOOP_C_356 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001111111");
        state_var_NS <= COMP_LOOP_C_357;
      WHEN COMP_LOOP_C_357 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010000000");
        state_var_NS <= COMP_LOOP_C_358;
      WHEN COMP_LOOP_C_358 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010000001");
        state_var_NS <= COMP_LOOP_C_359;
      WHEN COMP_LOOP_C_359 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010000010");
        state_var_NS <= COMP_LOOP_C_360;
      WHEN COMP_LOOP_C_360 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010000011");
        state_var_NS <= COMP_LOOP_C_361;
      WHEN COMP_LOOP_C_361 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010000100");
        state_var_NS <= COMP_LOOP_C_362;
      WHEN COMP_LOOP_C_362 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010000101");
        state_var_NS <= COMP_LOOP_C_363;
      WHEN COMP_LOOP_C_363 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010000110");
        state_var_NS <= COMP_LOOP_C_364;
      WHEN COMP_LOOP_C_364 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010000111");
        state_var_NS <= COMP_LOOP_C_365;
      WHEN COMP_LOOP_C_365 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010001000");
        state_var_NS <= COMP_LOOP_C_366;
      WHEN COMP_LOOP_C_366 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010001001");
        state_var_NS <= COMP_LOOP_C_367;
      WHEN COMP_LOOP_C_367 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010001010");
        state_var_NS <= COMP_LOOP_C_368;
      WHEN COMP_LOOP_C_368 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010001011");
        state_var_NS <= COMP_LOOP_C_369;
      WHEN COMP_LOOP_C_369 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010001100");
        state_var_NS <= COMP_LOOP_C_370;
      WHEN COMP_LOOP_C_370 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010001101");
        state_var_NS <= COMP_LOOP_C_371;
      WHEN COMP_LOOP_C_371 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010001110");
        state_var_NS <= COMP_LOOP_C_372;
      WHEN COMP_LOOP_C_372 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010001111");
        state_var_NS <= COMP_LOOP_C_373;
      WHEN COMP_LOOP_C_373 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010010000");
        state_var_NS <= COMP_LOOP_C_374;
      WHEN COMP_LOOP_C_374 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010010001");
        state_var_NS <= COMP_LOOP_C_375;
      WHEN COMP_LOOP_C_375 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010010010");
        state_var_NS <= COMP_LOOP_C_376;
      WHEN COMP_LOOP_C_376 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010010011");
        state_var_NS <= COMP_LOOP_C_377;
      WHEN COMP_LOOP_C_377 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010010100");
        state_var_NS <= COMP_LOOP_C_378;
      WHEN COMP_LOOP_C_378 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010010101");
        state_var_NS <= COMP_LOOP_C_379;
      WHEN COMP_LOOP_C_379 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010010110");
        state_var_NS <= COMP_LOOP_C_380;
      WHEN COMP_LOOP_C_380 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010010111");
        state_var_NS <= COMP_LOOP_C_381;
      WHEN COMP_LOOP_C_381 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010011000");
        state_var_NS <= COMP_LOOP_C_382;
      WHEN COMP_LOOP_C_382 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010011001");
        state_var_NS <= COMP_LOOP_C_383;
      WHEN COMP_LOOP_C_383 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010011010");
        state_var_NS <= COMP_LOOP_C_384;
      WHEN COMP_LOOP_C_384 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010011011");
        IF ( COMP_LOOP_C_384_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_385;
        END IF;
      WHEN COMP_LOOP_C_385 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010011100");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_0;
      WHEN COMP_LOOP_7_modExp_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010011101");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_1;
      WHEN COMP_LOOP_7_modExp_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010011110");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_2;
      WHEN COMP_LOOP_7_modExp_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010011111");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_3;
      WHEN COMP_LOOP_7_modExp_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010100000");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_4;
      WHEN COMP_LOOP_7_modExp_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010100001");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_5;
      WHEN COMP_LOOP_7_modExp_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010100010");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_6;
      WHEN COMP_LOOP_7_modExp_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010100011");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_7;
      WHEN COMP_LOOP_7_modExp_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010100100");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_8;
      WHEN COMP_LOOP_7_modExp_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010100101");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_9;
      WHEN COMP_LOOP_7_modExp_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010100110");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_10;
      WHEN COMP_LOOP_7_modExp_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010100111");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_11;
      WHEN COMP_LOOP_7_modExp_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010101000");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_12;
      WHEN COMP_LOOP_7_modExp_1_while_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010101001");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_13;
      WHEN COMP_LOOP_7_modExp_1_while_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010101010");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_14;
      WHEN COMP_LOOP_7_modExp_1_while_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010101011");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_15;
      WHEN COMP_LOOP_7_modExp_1_while_C_15 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010101100");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_16;
      WHEN COMP_LOOP_7_modExp_1_while_C_16 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010101101");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_17;
      WHEN COMP_LOOP_7_modExp_1_while_C_17 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010101110");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_18;
      WHEN COMP_LOOP_7_modExp_1_while_C_18 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010101111");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_19;
      WHEN COMP_LOOP_7_modExp_1_while_C_19 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010110000");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_20;
      WHEN COMP_LOOP_7_modExp_1_while_C_20 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010110001");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_21;
      WHEN COMP_LOOP_7_modExp_1_while_C_21 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010110010");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_22;
      WHEN COMP_LOOP_7_modExp_1_while_C_22 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010110011");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_23;
      WHEN COMP_LOOP_7_modExp_1_while_C_23 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010110100");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_24;
      WHEN COMP_LOOP_7_modExp_1_while_C_24 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010110101");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_25;
      WHEN COMP_LOOP_7_modExp_1_while_C_25 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010110110");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_26;
      WHEN COMP_LOOP_7_modExp_1_while_C_26 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010110111");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_27;
      WHEN COMP_LOOP_7_modExp_1_while_C_27 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010111000");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_28;
      WHEN COMP_LOOP_7_modExp_1_while_C_28 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010111001");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_29;
      WHEN COMP_LOOP_7_modExp_1_while_C_29 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010111010");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_30;
      WHEN COMP_LOOP_7_modExp_1_while_C_30 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010111011");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_31;
      WHEN COMP_LOOP_7_modExp_1_while_C_31 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010111100");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_32;
      WHEN COMP_LOOP_7_modExp_1_while_C_32 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010111101");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_33;
      WHEN COMP_LOOP_7_modExp_1_while_C_33 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010111110");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_34;
      WHEN COMP_LOOP_7_modExp_1_while_C_34 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010111111");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_35;
      WHEN COMP_LOOP_7_modExp_1_while_C_35 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011000000");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_36;
      WHEN COMP_LOOP_7_modExp_1_while_C_36 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011000001");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_37;
      WHEN COMP_LOOP_7_modExp_1_while_C_37 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011000010");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_38;
      WHEN COMP_LOOP_7_modExp_1_while_C_38 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011000011");
        IF ( COMP_LOOP_7_modExp_1_while_C_38_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_386;
        ELSE
          state_var_NS <= COMP_LOOP_7_modExp_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_386 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011000100");
        state_var_NS <= COMP_LOOP_C_387;
      WHEN COMP_LOOP_C_387 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011000101");
        state_var_NS <= COMP_LOOP_C_388;
      WHEN COMP_LOOP_C_388 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011000110");
        state_var_NS <= COMP_LOOP_C_389;
      WHEN COMP_LOOP_C_389 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011000111");
        state_var_NS <= COMP_LOOP_C_390;
      WHEN COMP_LOOP_C_390 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011001000");
        state_var_NS <= COMP_LOOP_C_391;
      WHEN COMP_LOOP_C_391 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011001001");
        state_var_NS <= COMP_LOOP_C_392;
      WHEN COMP_LOOP_C_392 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011001010");
        state_var_NS <= COMP_LOOP_C_393;
      WHEN COMP_LOOP_C_393 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011001011");
        state_var_NS <= COMP_LOOP_C_394;
      WHEN COMP_LOOP_C_394 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011001100");
        state_var_NS <= COMP_LOOP_C_395;
      WHEN COMP_LOOP_C_395 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011001101");
        state_var_NS <= COMP_LOOP_C_396;
      WHEN COMP_LOOP_C_396 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011001110");
        state_var_NS <= COMP_LOOP_C_397;
      WHEN COMP_LOOP_C_397 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011001111");
        state_var_NS <= COMP_LOOP_C_398;
      WHEN COMP_LOOP_C_398 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011010000");
        state_var_NS <= COMP_LOOP_C_399;
      WHEN COMP_LOOP_C_399 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011010001");
        state_var_NS <= COMP_LOOP_C_400;
      WHEN COMP_LOOP_C_400 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011010010");
        state_var_NS <= COMP_LOOP_C_401;
      WHEN COMP_LOOP_C_401 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011010011");
        state_var_NS <= COMP_LOOP_C_402;
      WHEN COMP_LOOP_C_402 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011010100");
        state_var_NS <= COMP_LOOP_C_403;
      WHEN COMP_LOOP_C_403 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011010101");
        state_var_NS <= COMP_LOOP_C_404;
      WHEN COMP_LOOP_C_404 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011010110");
        state_var_NS <= COMP_LOOP_C_405;
      WHEN COMP_LOOP_C_405 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011010111");
        state_var_NS <= COMP_LOOP_C_406;
      WHEN COMP_LOOP_C_406 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011011000");
        state_var_NS <= COMP_LOOP_C_407;
      WHEN COMP_LOOP_C_407 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011011001");
        state_var_NS <= COMP_LOOP_C_408;
      WHEN COMP_LOOP_C_408 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011011010");
        state_var_NS <= COMP_LOOP_C_409;
      WHEN COMP_LOOP_C_409 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011011011");
        state_var_NS <= COMP_LOOP_C_410;
      WHEN COMP_LOOP_C_410 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011011100");
        state_var_NS <= COMP_LOOP_C_411;
      WHEN COMP_LOOP_C_411 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011011101");
        state_var_NS <= COMP_LOOP_C_412;
      WHEN COMP_LOOP_C_412 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011011110");
        state_var_NS <= COMP_LOOP_C_413;
      WHEN COMP_LOOP_C_413 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011011111");
        state_var_NS <= COMP_LOOP_C_414;
      WHEN COMP_LOOP_C_414 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011100000");
        state_var_NS <= COMP_LOOP_C_415;
      WHEN COMP_LOOP_C_415 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011100001");
        state_var_NS <= COMP_LOOP_C_416;
      WHEN COMP_LOOP_C_416 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011100010");
        state_var_NS <= COMP_LOOP_C_417;
      WHEN COMP_LOOP_C_417 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011100011");
        state_var_NS <= COMP_LOOP_C_418;
      WHEN COMP_LOOP_C_418 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011100100");
        state_var_NS <= COMP_LOOP_C_419;
      WHEN COMP_LOOP_C_419 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011100101");
        state_var_NS <= COMP_LOOP_C_420;
      WHEN COMP_LOOP_C_420 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011100110");
        state_var_NS <= COMP_LOOP_C_421;
      WHEN COMP_LOOP_C_421 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011100111");
        state_var_NS <= COMP_LOOP_C_422;
      WHEN COMP_LOOP_C_422 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011101000");
        state_var_NS <= COMP_LOOP_C_423;
      WHEN COMP_LOOP_C_423 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011101001");
        state_var_NS <= COMP_LOOP_C_424;
      WHEN COMP_LOOP_C_424 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011101010");
        state_var_NS <= COMP_LOOP_C_425;
      WHEN COMP_LOOP_C_425 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011101011");
        state_var_NS <= COMP_LOOP_C_426;
      WHEN COMP_LOOP_C_426 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011101100");
        state_var_NS <= COMP_LOOP_C_427;
      WHEN COMP_LOOP_C_427 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011101101");
        state_var_NS <= COMP_LOOP_C_428;
      WHEN COMP_LOOP_C_428 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011101110");
        state_var_NS <= COMP_LOOP_C_429;
      WHEN COMP_LOOP_C_429 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011101111");
        state_var_NS <= COMP_LOOP_C_430;
      WHEN COMP_LOOP_C_430 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011110000");
        state_var_NS <= COMP_LOOP_C_431;
      WHEN COMP_LOOP_C_431 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011110001");
        state_var_NS <= COMP_LOOP_C_432;
      WHEN COMP_LOOP_C_432 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011110010");
        state_var_NS <= COMP_LOOP_C_433;
      WHEN COMP_LOOP_C_433 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011110011");
        state_var_NS <= COMP_LOOP_C_434;
      WHEN COMP_LOOP_C_434 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011110100");
        state_var_NS <= COMP_LOOP_C_435;
      WHEN COMP_LOOP_C_435 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011110101");
        state_var_NS <= COMP_LOOP_C_436;
      WHEN COMP_LOOP_C_436 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011110110");
        state_var_NS <= COMP_LOOP_C_437;
      WHEN COMP_LOOP_C_437 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011110111");
        state_var_NS <= COMP_LOOP_C_438;
      WHEN COMP_LOOP_C_438 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011111000");
        state_var_NS <= COMP_LOOP_C_439;
      WHEN COMP_LOOP_C_439 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011111001");
        state_var_NS <= COMP_LOOP_C_440;
      WHEN COMP_LOOP_C_440 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011111010");
        state_var_NS <= COMP_LOOP_C_441;
      WHEN COMP_LOOP_C_441 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011111011");
        state_var_NS <= COMP_LOOP_C_442;
      WHEN COMP_LOOP_C_442 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011111100");
        state_var_NS <= COMP_LOOP_C_443;
      WHEN COMP_LOOP_C_443 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011111101");
        state_var_NS <= COMP_LOOP_C_444;
      WHEN COMP_LOOP_C_444 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011111110");
        state_var_NS <= COMP_LOOP_C_445;
      WHEN COMP_LOOP_C_445 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011111111");
        state_var_NS <= COMP_LOOP_C_446;
      WHEN COMP_LOOP_C_446 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100000000");
        state_var_NS <= COMP_LOOP_C_447;
      WHEN COMP_LOOP_C_447 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100000001");
        state_var_NS <= COMP_LOOP_C_448;
      WHEN COMP_LOOP_C_448 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100000010");
        IF ( COMP_LOOP_C_448_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_449;
        END IF;
      WHEN COMP_LOOP_C_449 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100000011");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_0;
      WHEN COMP_LOOP_8_modExp_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100000100");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_1;
      WHEN COMP_LOOP_8_modExp_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100000101");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_2;
      WHEN COMP_LOOP_8_modExp_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100000110");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_3;
      WHEN COMP_LOOP_8_modExp_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100000111");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_4;
      WHEN COMP_LOOP_8_modExp_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100001000");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_5;
      WHEN COMP_LOOP_8_modExp_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100001001");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_6;
      WHEN COMP_LOOP_8_modExp_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100001010");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_7;
      WHEN COMP_LOOP_8_modExp_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100001011");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_8;
      WHEN COMP_LOOP_8_modExp_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100001100");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_9;
      WHEN COMP_LOOP_8_modExp_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100001101");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_10;
      WHEN COMP_LOOP_8_modExp_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100001110");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_11;
      WHEN COMP_LOOP_8_modExp_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100001111");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_12;
      WHEN COMP_LOOP_8_modExp_1_while_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100010000");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_13;
      WHEN COMP_LOOP_8_modExp_1_while_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100010001");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_14;
      WHEN COMP_LOOP_8_modExp_1_while_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100010010");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_15;
      WHEN COMP_LOOP_8_modExp_1_while_C_15 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100010011");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_16;
      WHEN COMP_LOOP_8_modExp_1_while_C_16 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100010100");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_17;
      WHEN COMP_LOOP_8_modExp_1_while_C_17 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100010101");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_18;
      WHEN COMP_LOOP_8_modExp_1_while_C_18 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100010110");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_19;
      WHEN COMP_LOOP_8_modExp_1_while_C_19 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100010111");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_20;
      WHEN COMP_LOOP_8_modExp_1_while_C_20 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100011000");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_21;
      WHEN COMP_LOOP_8_modExp_1_while_C_21 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100011001");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_22;
      WHEN COMP_LOOP_8_modExp_1_while_C_22 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100011010");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_23;
      WHEN COMP_LOOP_8_modExp_1_while_C_23 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100011011");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_24;
      WHEN COMP_LOOP_8_modExp_1_while_C_24 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100011100");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_25;
      WHEN COMP_LOOP_8_modExp_1_while_C_25 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100011101");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_26;
      WHEN COMP_LOOP_8_modExp_1_while_C_26 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100011110");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_27;
      WHEN COMP_LOOP_8_modExp_1_while_C_27 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100011111");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_28;
      WHEN COMP_LOOP_8_modExp_1_while_C_28 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100100000");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_29;
      WHEN COMP_LOOP_8_modExp_1_while_C_29 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100100001");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_30;
      WHEN COMP_LOOP_8_modExp_1_while_C_30 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100100010");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_31;
      WHEN COMP_LOOP_8_modExp_1_while_C_31 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100100011");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_32;
      WHEN COMP_LOOP_8_modExp_1_while_C_32 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100100100");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_33;
      WHEN COMP_LOOP_8_modExp_1_while_C_33 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100100101");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_34;
      WHEN COMP_LOOP_8_modExp_1_while_C_34 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100100110");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_35;
      WHEN COMP_LOOP_8_modExp_1_while_C_35 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100100111");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_36;
      WHEN COMP_LOOP_8_modExp_1_while_C_36 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100101000");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_37;
      WHEN COMP_LOOP_8_modExp_1_while_C_37 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100101001");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_38;
      WHEN COMP_LOOP_8_modExp_1_while_C_38 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100101010");
        IF ( COMP_LOOP_8_modExp_1_while_C_38_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_450;
        ELSE
          state_var_NS <= COMP_LOOP_8_modExp_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_450 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100101011");
        state_var_NS <= COMP_LOOP_C_451;
      WHEN COMP_LOOP_C_451 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100101100");
        state_var_NS <= COMP_LOOP_C_452;
      WHEN COMP_LOOP_C_452 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100101101");
        state_var_NS <= COMP_LOOP_C_453;
      WHEN COMP_LOOP_C_453 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100101110");
        state_var_NS <= COMP_LOOP_C_454;
      WHEN COMP_LOOP_C_454 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100101111");
        state_var_NS <= COMP_LOOP_C_455;
      WHEN COMP_LOOP_C_455 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100110000");
        state_var_NS <= COMP_LOOP_C_456;
      WHEN COMP_LOOP_C_456 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100110001");
        state_var_NS <= COMP_LOOP_C_457;
      WHEN COMP_LOOP_C_457 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100110010");
        state_var_NS <= COMP_LOOP_C_458;
      WHEN COMP_LOOP_C_458 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100110011");
        state_var_NS <= COMP_LOOP_C_459;
      WHEN COMP_LOOP_C_459 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100110100");
        state_var_NS <= COMP_LOOP_C_460;
      WHEN COMP_LOOP_C_460 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100110101");
        state_var_NS <= COMP_LOOP_C_461;
      WHEN COMP_LOOP_C_461 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100110110");
        state_var_NS <= COMP_LOOP_C_462;
      WHEN COMP_LOOP_C_462 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100110111");
        state_var_NS <= COMP_LOOP_C_463;
      WHEN COMP_LOOP_C_463 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100111000");
        state_var_NS <= COMP_LOOP_C_464;
      WHEN COMP_LOOP_C_464 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100111001");
        state_var_NS <= COMP_LOOP_C_465;
      WHEN COMP_LOOP_C_465 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100111010");
        state_var_NS <= COMP_LOOP_C_466;
      WHEN COMP_LOOP_C_466 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100111011");
        state_var_NS <= COMP_LOOP_C_467;
      WHEN COMP_LOOP_C_467 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100111100");
        state_var_NS <= COMP_LOOP_C_468;
      WHEN COMP_LOOP_C_468 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100111101");
        state_var_NS <= COMP_LOOP_C_469;
      WHEN COMP_LOOP_C_469 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100111110");
        state_var_NS <= COMP_LOOP_C_470;
      WHEN COMP_LOOP_C_470 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100111111");
        state_var_NS <= COMP_LOOP_C_471;
      WHEN COMP_LOOP_C_471 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101000000");
        state_var_NS <= COMP_LOOP_C_472;
      WHEN COMP_LOOP_C_472 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101000001");
        state_var_NS <= COMP_LOOP_C_473;
      WHEN COMP_LOOP_C_473 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101000010");
        state_var_NS <= COMP_LOOP_C_474;
      WHEN COMP_LOOP_C_474 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101000011");
        state_var_NS <= COMP_LOOP_C_475;
      WHEN COMP_LOOP_C_475 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101000100");
        state_var_NS <= COMP_LOOP_C_476;
      WHEN COMP_LOOP_C_476 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101000101");
        state_var_NS <= COMP_LOOP_C_477;
      WHEN COMP_LOOP_C_477 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101000110");
        state_var_NS <= COMP_LOOP_C_478;
      WHEN COMP_LOOP_C_478 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101000111");
        state_var_NS <= COMP_LOOP_C_479;
      WHEN COMP_LOOP_C_479 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101001000");
        state_var_NS <= COMP_LOOP_C_480;
      WHEN COMP_LOOP_C_480 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101001001");
        state_var_NS <= COMP_LOOP_C_481;
      WHEN COMP_LOOP_C_481 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101001010");
        state_var_NS <= COMP_LOOP_C_482;
      WHEN COMP_LOOP_C_482 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101001011");
        state_var_NS <= COMP_LOOP_C_483;
      WHEN COMP_LOOP_C_483 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101001100");
        state_var_NS <= COMP_LOOP_C_484;
      WHEN COMP_LOOP_C_484 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101001101");
        state_var_NS <= COMP_LOOP_C_485;
      WHEN COMP_LOOP_C_485 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101001110");
        state_var_NS <= COMP_LOOP_C_486;
      WHEN COMP_LOOP_C_486 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101001111");
        state_var_NS <= COMP_LOOP_C_487;
      WHEN COMP_LOOP_C_487 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101010000");
        state_var_NS <= COMP_LOOP_C_488;
      WHEN COMP_LOOP_C_488 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101010001");
        state_var_NS <= COMP_LOOP_C_489;
      WHEN COMP_LOOP_C_489 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101010010");
        state_var_NS <= COMP_LOOP_C_490;
      WHEN COMP_LOOP_C_490 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101010011");
        state_var_NS <= COMP_LOOP_C_491;
      WHEN COMP_LOOP_C_491 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101010100");
        state_var_NS <= COMP_LOOP_C_492;
      WHEN COMP_LOOP_C_492 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101010101");
        state_var_NS <= COMP_LOOP_C_493;
      WHEN COMP_LOOP_C_493 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101010110");
        state_var_NS <= COMP_LOOP_C_494;
      WHEN COMP_LOOP_C_494 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101010111");
        state_var_NS <= COMP_LOOP_C_495;
      WHEN COMP_LOOP_C_495 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101011000");
        state_var_NS <= COMP_LOOP_C_496;
      WHEN COMP_LOOP_C_496 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101011001");
        state_var_NS <= COMP_LOOP_C_497;
      WHEN COMP_LOOP_C_497 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101011010");
        state_var_NS <= COMP_LOOP_C_498;
      WHEN COMP_LOOP_C_498 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101011011");
        state_var_NS <= COMP_LOOP_C_499;
      WHEN COMP_LOOP_C_499 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101011100");
        state_var_NS <= COMP_LOOP_C_500;
      WHEN COMP_LOOP_C_500 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101011101");
        state_var_NS <= COMP_LOOP_C_501;
      WHEN COMP_LOOP_C_501 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101011110");
        state_var_NS <= COMP_LOOP_C_502;
      WHEN COMP_LOOP_C_502 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101011111");
        state_var_NS <= COMP_LOOP_C_503;
      WHEN COMP_LOOP_C_503 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101100000");
        state_var_NS <= COMP_LOOP_C_504;
      WHEN COMP_LOOP_C_504 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101100001");
        state_var_NS <= COMP_LOOP_C_505;
      WHEN COMP_LOOP_C_505 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101100010");
        state_var_NS <= COMP_LOOP_C_506;
      WHEN COMP_LOOP_C_506 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101100011");
        state_var_NS <= COMP_LOOP_C_507;
      WHEN COMP_LOOP_C_507 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101100100");
        state_var_NS <= COMP_LOOP_C_508;
      WHEN COMP_LOOP_C_508 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101100101");
        state_var_NS <= COMP_LOOP_C_509;
      WHEN COMP_LOOP_C_509 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101100110");
        state_var_NS <= COMP_LOOP_C_510;
      WHEN COMP_LOOP_C_510 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101100111");
        state_var_NS <= COMP_LOOP_C_511;
      WHEN COMP_LOOP_C_511 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101101000");
        state_var_NS <= COMP_LOOP_C_512;
      WHEN COMP_LOOP_C_512 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101101001");
        IF ( COMP_LOOP_C_512_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_513;
        END IF;
      WHEN COMP_LOOP_C_513 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101101010");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_0;
      WHEN COMP_LOOP_9_modExp_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101101011");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_1;
      WHEN COMP_LOOP_9_modExp_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101101100");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_2;
      WHEN COMP_LOOP_9_modExp_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101101101");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_3;
      WHEN COMP_LOOP_9_modExp_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101101110");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_4;
      WHEN COMP_LOOP_9_modExp_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101101111");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_5;
      WHEN COMP_LOOP_9_modExp_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101110000");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_6;
      WHEN COMP_LOOP_9_modExp_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101110001");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_7;
      WHEN COMP_LOOP_9_modExp_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101110010");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_8;
      WHEN COMP_LOOP_9_modExp_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101110011");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_9;
      WHEN COMP_LOOP_9_modExp_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101110100");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_10;
      WHEN COMP_LOOP_9_modExp_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101110101");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_11;
      WHEN COMP_LOOP_9_modExp_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101110110");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_12;
      WHEN COMP_LOOP_9_modExp_1_while_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101110111");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_13;
      WHEN COMP_LOOP_9_modExp_1_while_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101111000");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_14;
      WHEN COMP_LOOP_9_modExp_1_while_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101111001");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_15;
      WHEN COMP_LOOP_9_modExp_1_while_C_15 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101111010");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_16;
      WHEN COMP_LOOP_9_modExp_1_while_C_16 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101111011");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_17;
      WHEN COMP_LOOP_9_modExp_1_while_C_17 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101111100");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_18;
      WHEN COMP_LOOP_9_modExp_1_while_C_18 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101111101");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_19;
      WHEN COMP_LOOP_9_modExp_1_while_C_19 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101111110");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_20;
      WHEN COMP_LOOP_9_modExp_1_while_C_20 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101111111");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_21;
      WHEN COMP_LOOP_9_modExp_1_while_C_21 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110000000");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_22;
      WHEN COMP_LOOP_9_modExp_1_while_C_22 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110000001");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_23;
      WHEN COMP_LOOP_9_modExp_1_while_C_23 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110000010");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_24;
      WHEN COMP_LOOP_9_modExp_1_while_C_24 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110000011");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_25;
      WHEN COMP_LOOP_9_modExp_1_while_C_25 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110000100");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_26;
      WHEN COMP_LOOP_9_modExp_1_while_C_26 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110000101");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_27;
      WHEN COMP_LOOP_9_modExp_1_while_C_27 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110000110");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_28;
      WHEN COMP_LOOP_9_modExp_1_while_C_28 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110000111");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_29;
      WHEN COMP_LOOP_9_modExp_1_while_C_29 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110001000");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_30;
      WHEN COMP_LOOP_9_modExp_1_while_C_30 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110001001");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_31;
      WHEN COMP_LOOP_9_modExp_1_while_C_31 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110001010");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_32;
      WHEN COMP_LOOP_9_modExp_1_while_C_32 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110001011");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_33;
      WHEN COMP_LOOP_9_modExp_1_while_C_33 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110001100");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_34;
      WHEN COMP_LOOP_9_modExp_1_while_C_34 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110001101");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_35;
      WHEN COMP_LOOP_9_modExp_1_while_C_35 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110001110");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_36;
      WHEN COMP_LOOP_9_modExp_1_while_C_36 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110001111");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_37;
      WHEN COMP_LOOP_9_modExp_1_while_C_37 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110010000");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_38;
      WHEN COMP_LOOP_9_modExp_1_while_C_38 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110010001");
        IF ( COMP_LOOP_9_modExp_1_while_C_38_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_514;
        ELSE
          state_var_NS <= COMP_LOOP_9_modExp_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_514 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110010010");
        state_var_NS <= COMP_LOOP_C_515;
      WHEN COMP_LOOP_C_515 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110010011");
        state_var_NS <= COMP_LOOP_C_516;
      WHEN COMP_LOOP_C_516 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110010100");
        state_var_NS <= COMP_LOOP_C_517;
      WHEN COMP_LOOP_C_517 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110010101");
        state_var_NS <= COMP_LOOP_C_518;
      WHEN COMP_LOOP_C_518 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110010110");
        state_var_NS <= COMP_LOOP_C_519;
      WHEN COMP_LOOP_C_519 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110010111");
        state_var_NS <= COMP_LOOP_C_520;
      WHEN COMP_LOOP_C_520 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110011000");
        state_var_NS <= COMP_LOOP_C_521;
      WHEN COMP_LOOP_C_521 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110011001");
        state_var_NS <= COMP_LOOP_C_522;
      WHEN COMP_LOOP_C_522 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110011010");
        state_var_NS <= COMP_LOOP_C_523;
      WHEN COMP_LOOP_C_523 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110011011");
        state_var_NS <= COMP_LOOP_C_524;
      WHEN COMP_LOOP_C_524 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110011100");
        state_var_NS <= COMP_LOOP_C_525;
      WHEN COMP_LOOP_C_525 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110011101");
        state_var_NS <= COMP_LOOP_C_526;
      WHEN COMP_LOOP_C_526 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110011110");
        state_var_NS <= COMP_LOOP_C_527;
      WHEN COMP_LOOP_C_527 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110011111");
        state_var_NS <= COMP_LOOP_C_528;
      WHEN COMP_LOOP_C_528 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110100000");
        state_var_NS <= COMP_LOOP_C_529;
      WHEN COMP_LOOP_C_529 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110100001");
        state_var_NS <= COMP_LOOP_C_530;
      WHEN COMP_LOOP_C_530 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110100010");
        state_var_NS <= COMP_LOOP_C_531;
      WHEN COMP_LOOP_C_531 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110100011");
        state_var_NS <= COMP_LOOP_C_532;
      WHEN COMP_LOOP_C_532 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110100100");
        state_var_NS <= COMP_LOOP_C_533;
      WHEN COMP_LOOP_C_533 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110100101");
        state_var_NS <= COMP_LOOP_C_534;
      WHEN COMP_LOOP_C_534 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110100110");
        state_var_NS <= COMP_LOOP_C_535;
      WHEN COMP_LOOP_C_535 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110100111");
        state_var_NS <= COMP_LOOP_C_536;
      WHEN COMP_LOOP_C_536 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110101000");
        state_var_NS <= COMP_LOOP_C_537;
      WHEN COMP_LOOP_C_537 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110101001");
        state_var_NS <= COMP_LOOP_C_538;
      WHEN COMP_LOOP_C_538 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110101010");
        state_var_NS <= COMP_LOOP_C_539;
      WHEN COMP_LOOP_C_539 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110101011");
        state_var_NS <= COMP_LOOP_C_540;
      WHEN COMP_LOOP_C_540 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110101100");
        state_var_NS <= COMP_LOOP_C_541;
      WHEN COMP_LOOP_C_541 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110101101");
        state_var_NS <= COMP_LOOP_C_542;
      WHEN COMP_LOOP_C_542 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110101110");
        state_var_NS <= COMP_LOOP_C_543;
      WHEN COMP_LOOP_C_543 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110101111");
        state_var_NS <= COMP_LOOP_C_544;
      WHEN COMP_LOOP_C_544 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110110000");
        state_var_NS <= COMP_LOOP_C_545;
      WHEN COMP_LOOP_C_545 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110110001");
        state_var_NS <= COMP_LOOP_C_546;
      WHEN COMP_LOOP_C_546 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110110010");
        state_var_NS <= COMP_LOOP_C_547;
      WHEN COMP_LOOP_C_547 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110110011");
        state_var_NS <= COMP_LOOP_C_548;
      WHEN COMP_LOOP_C_548 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110110100");
        state_var_NS <= COMP_LOOP_C_549;
      WHEN COMP_LOOP_C_549 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110110101");
        state_var_NS <= COMP_LOOP_C_550;
      WHEN COMP_LOOP_C_550 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110110110");
        state_var_NS <= COMP_LOOP_C_551;
      WHEN COMP_LOOP_C_551 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110110111");
        state_var_NS <= COMP_LOOP_C_552;
      WHEN COMP_LOOP_C_552 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110111000");
        state_var_NS <= COMP_LOOP_C_553;
      WHEN COMP_LOOP_C_553 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110111001");
        state_var_NS <= COMP_LOOP_C_554;
      WHEN COMP_LOOP_C_554 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110111010");
        state_var_NS <= COMP_LOOP_C_555;
      WHEN COMP_LOOP_C_555 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110111011");
        state_var_NS <= COMP_LOOP_C_556;
      WHEN COMP_LOOP_C_556 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110111100");
        state_var_NS <= COMP_LOOP_C_557;
      WHEN COMP_LOOP_C_557 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110111101");
        state_var_NS <= COMP_LOOP_C_558;
      WHEN COMP_LOOP_C_558 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110111110");
        state_var_NS <= COMP_LOOP_C_559;
      WHEN COMP_LOOP_C_559 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110111111");
        state_var_NS <= COMP_LOOP_C_560;
      WHEN COMP_LOOP_C_560 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111000000");
        state_var_NS <= COMP_LOOP_C_561;
      WHEN COMP_LOOP_C_561 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111000001");
        state_var_NS <= COMP_LOOP_C_562;
      WHEN COMP_LOOP_C_562 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111000010");
        state_var_NS <= COMP_LOOP_C_563;
      WHEN COMP_LOOP_C_563 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111000011");
        state_var_NS <= COMP_LOOP_C_564;
      WHEN COMP_LOOP_C_564 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111000100");
        state_var_NS <= COMP_LOOP_C_565;
      WHEN COMP_LOOP_C_565 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111000101");
        state_var_NS <= COMP_LOOP_C_566;
      WHEN COMP_LOOP_C_566 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111000110");
        state_var_NS <= COMP_LOOP_C_567;
      WHEN COMP_LOOP_C_567 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111000111");
        state_var_NS <= COMP_LOOP_C_568;
      WHEN COMP_LOOP_C_568 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111001000");
        state_var_NS <= COMP_LOOP_C_569;
      WHEN COMP_LOOP_C_569 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111001001");
        state_var_NS <= COMP_LOOP_C_570;
      WHEN COMP_LOOP_C_570 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111001010");
        state_var_NS <= COMP_LOOP_C_571;
      WHEN COMP_LOOP_C_571 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111001011");
        state_var_NS <= COMP_LOOP_C_572;
      WHEN COMP_LOOP_C_572 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111001100");
        state_var_NS <= COMP_LOOP_C_573;
      WHEN COMP_LOOP_C_573 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111001101");
        state_var_NS <= COMP_LOOP_C_574;
      WHEN COMP_LOOP_C_574 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111001110");
        state_var_NS <= COMP_LOOP_C_575;
      WHEN COMP_LOOP_C_575 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111001111");
        state_var_NS <= COMP_LOOP_C_576;
      WHEN COMP_LOOP_C_576 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111010000");
        IF ( COMP_LOOP_C_576_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_577;
        END IF;
      WHEN COMP_LOOP_C_577 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111010001");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_0;
      WHEN COMP_LOOP_10_modExp_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111010010");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_1;
      WHEN COMP_LOOP_10_modExp_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111010011");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_2;
      WHEN COMP_LOOP_10_modExp_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111010100");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_3;
      WHEN COMP_LOOP_10_modExp_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111010101");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_4;
      WHEN COMP_LOOP_10_modExp_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111010110");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_5;
      WHEN COMP_LOOP_10_modExp_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111010111");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_6;
      WHEN COMP_LOOP_10_modExp_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111011000");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_7;
      WHEN COMP_LOOP_10_modExp_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111011001");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_8;
      WHEN COMP_LOOP_10_modExp_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111011010");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_9;
      WHEN COMP_LOOP_10_modExp_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111011011");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_10;
      WHEN COMP_LOOP_10_modExp_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111011100");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_11;
      WHEN COMP_LOOP_10_modExp_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111011101");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_12;
      WHEN COMP_LOOP_10_modExp_1_while_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111011110");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_13;
      WHEN COMP_LOOP_10_modExp_1_while_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111011111");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_14;
      WHEN COMP_LOOP_10_modExp_1_while_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111100000");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_15;
      WHEN COMP_LOOP_10_modExp_1_while_C_15 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111100001");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_16;
      WHEN COMP_LOOP_10_modExp_1_while_C_16 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111100010");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_17;
      WHEN COMP_LOOP_10_modExp_1_while_C_17 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111100011");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_18;
      WHEN COMP_LOOP_10_modExp_1_while_C_18 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111100100");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_19;
      WHEN COMP_LOOP_10_modExp_1_while_C_19 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111100101");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_20;
      WHEN COMP_LOOP_10_modExp_1_while_C_20 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111100110");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_21;
      WHEN COMP_LOOP_10_modExp_1_while_C_21 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111100111");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_22;
      WHEN COMP_LOOP_10_modExp_1_while_C_22 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111101000");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_23;
      WHEN COMP_LOOP_10_modExp_1_while_C_23 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111101001");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_24;
      WHEN COMP_LOOP_10_modExp_1_while_C_24 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111101010");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_25;
      WHEN COMP_LOOP_10_modExp_1_while_C_25 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111101011");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_26;
      WHEN COMP_LOOP_10_modExp_1_while_C_26 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111101100");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_27;
      WHEN COMP_LOOP_10_modExp_1_while_C_27 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111101101");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_28;
      WHEN COMP_LOOP_10_modExp_1_while_C_28 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111101110");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_29;
      WHEN COMP_LOOP_10_modExp_1_while_C_29 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111101111");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_30;
      WHEN COMP_LOOP_10_modExp_1_while_C_30 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111110000");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_31;
      WHEN COMP_LOOP_10_modExp_1_while_C_31 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111110001");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_32;
      WHEN COMP_LOOP_10_modExp_1_while_C_32 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111110010");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_33;
      WHEN COMP_LOOP_10_modExp_1_while_C_33 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111110011");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_34;
      WHEN COMP_LOOP_10_modExp_1_while_C_34 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111110100");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_35;
      WHEN COMP_LOOP_10_modExp_1_while_C_35 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111110101");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_36;
      WHEN COMP_LOOP_10_modExp_1_while_C_36 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111110110");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_37;
      WHEN COMP_LOOP_10_modExp_1_while_C_37 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111110111");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_38;
      WHEN COMP_LOOP_10_modExp_1_while_C_38 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111111000");
        IF ( COMP_LOOP_10_modExp_1_while_C_38_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_578;
        ELSE
          state_var_NS <= COMP_LOOP_10_modExp_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_578 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111111001");
        state_var_NS <= COMP_LOOP_C_579;
      WHEN COMP_LOOP_C_579 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111111010");
        state_var_NS <= COMP_LOOP_C_580;
      WHEN COMP_LOOP_C_580 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111111011");
        state_var_NS <= COMP_LOOP_C_581;
      WHEN COMP_LOOP_C_581 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111111100");
        state_var_NS <= COMP_LOOP_C_582;
      WHEN COMP_LOOP_C_582 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111111101");
        state_var_NS <= COMP_LOOP_C_583;
      WHEN COMP_LOOP_C_583 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111111110");
        state_var_NS <= COMP_LOOP_C_584;
      WHEN COMP_LOOP_C_584 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111111111");
        state_var_NS <= COMP_LOOP_C_585;
      WHEN COMP_LOOP_C_585 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000000000");
        state_var_NS <= COMP_LOOP_C_586;
      WHEN COMP_LOOP_C_586 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000000001");
        state_var_NS <= COMP_LOOP_C_587;
      WHEN COMP_LOOP_C_587 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000000010");
        state_var_NS <= COMP_LOOP_C_588;
      WHEN COMP_LOOP_C_588 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000000011");
        state_var_NS <= COMP_LOOP_C_589;
      WHEN COMP_LOOP_C_589 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000000100");
        state_var_NS <= COMP_LOOP_C_590;
      WHEN COMP_LOOP_C_590 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000000101");
        state_var_NS <= COMP_LOOP_C_591;
      WHEN COMP_LOOP_C_591 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000000110");
        state_var_NS <= COMP_LOOP_C_592;
      WHEN COMP_LOOP_C_592 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000000111");
        state_var_NS <= COMP_LOOP_C_593;
      WHEN COMP_LOOP_C_593 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000001000");
        state_var_NS <= COMP_LOOP_C_594;
      WHEN COMP_LOOP_C_594 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000001001");
        state_var_NS <= COMP_LOOP_C_595;
      WHEN COMP_LOOP_C_595 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000001010");
        state_var_NS <= COMP_LOOP_C_596;
      WHEN COMP_LOOP_C_596 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000001011");
        state_var_NS <= COMP_LOOP_C_597;
      WHEN COMP_LOOP_C_597 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000001100");
        state_var_NS <= COMP_LOOP_C_598;
      WHEN COMP_LOOP_C_598 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000001101");
        state_var_NS <= COMP_LOOP_C_599;
      WHEN COMP_LOOP_C_599 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000001110");
        state_var_NS <= COMP_LOOP_C_600;
      WHEN COMP_LOOP_C_600 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000001111");
        state_var_NS <= COMP_LOOP_C_601;
      WHEN COMP_LOOP_C_601 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000010000");
        state_var_NS <= COMP_LOOP_C_602;
      WHEN COMP_LOOP_C_602 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000010001");
        state_var_NS <= COMP_LOOP_C_603;
      WHEN COMP_LOOP_C_603 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000010010");
        state_var_NS <= COMP_LOOP_C_604;
      WHEN COMP_LOOP_C_604 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000010011");
        state_var_NS <= COMP_LOOP_C_605;
      WHEN COMP_LOOP_C_605 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000010100");
        state_var_NS <= COMP_LOOP_C_606;
      WHEN COMP_LOOP_C_606 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000010101");
        state_var_NS <= COMP_LOOP_C_607;
      WHEN COMP_LOOP_C_607 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000010110");
        state_var_NS <= COMP_LOOP_C_608;
      WHEN COMP_LOOP_C_608 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000010111");
        state_var_NS <= COMP_LOOP_C_609;
      WHEN COMP_LOOP_C_609 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000011000");
        state_var_NS <= COMP_LOOP_C_610;
      WHEN COMP_LOOP_C_610 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000011001");
        state_var_NS <= COMP_LOOP_C_611;
      WHEN COMP_LOOP_C_611 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000011010");
        state_var_NS <= COMP_LOOP_C_612;
      WHEN COMP_LOOP_C_612 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000011011");
        state_var_NS <= COMP_LOOP_C_613;
      WHEN COMP_LOOP_C_613 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000011100");
        state_var_NS <= COMP_LOOP_C_614;
      WHEN COMP_LOOP_C_614 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000011101");
        state_var_NS <= COMP_LOOP_C_615;
      WHEN COMP_LOOP_C_615 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000011110");
        state_var_NS <= COMP_LOOP_C_616;
      WHEN COMP_LOOP_C_616 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000011111");
        state_var_NS <= COMP_LOOP_C_617;
      WHEN COMP_LOOP_C_617 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000100000");
        state_var_NS <= COMP_LOOP_C_618;
      WHEN COMP_LOOP_C_618 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000100001");
        state_var_NS <= COMP_LOOP_C_619;
      WHEN COMP_LOOP_C_619 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000100010");
        state_var_NS <= COMP_LOOP_C_620;
      WHEN COMP_LOOP_C_620 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000100011");
        state_var_NS <= COMP_LOOP_C_621;
      WHEN COMP_LOOP_C_621 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000100100");
        state_var_NS <= COMP_LOOP_C_622;
      WHEN COMP_LOOP_C_622 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000100101");
        state_var_NS <= COMP_LOOP_C_623;
      WHEN COMP_LOOP_C_623 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000100110");
        state_var_NS <= COMP_LOOP_C_624;
      WHEN COMP_LOOP_C_624 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000100111");
        state_var_NS <= COMP_LOOP_C_625;
      WHEN COMP_LOOP_C_625 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000101000");
        state_var_NS <= COMP_LOOP_C_626;
      WHEN COMP_LOOP_C_626 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000101001");
        state_var_NS <= COMP_LOOP_C_627;
      WHEN COMP_LOOP_C_627 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000101010");
        state_var_NS <= COMP_LOOP_C_628;
      WHEN COMP_LOOP_C_628 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000101011");
        state_var_NS <= COMP_LOOP_C_629;
      WHEN COMP_LOOP_C_629 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000101100");
        state_var_NS <= COMP_LOOP_C_630;
      WHEN COMP_LOOP_C_630 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000101101");
        state_var_NS <= COMP_LOOP_C_631;
      WHEN COMP_LOOP_C_631 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000101110");
        state_var_NS <= COMP_LOOP_C_632;
      WHEN COMP_LOOP_C_632 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000101111");
        state_var_NS <= COMP_LOOP_C_633;
      WHEN COMP_LOOP_C_633 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000110000");
        state_var_NS <= COMP_LOOP_C_634;
      WHEN COMP_LOOP_C_634 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000110001");
        state_var_NS <= COMP_LOOP_C_635;
      WHEN COMP_LOOP_C_635 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000110010");
        state_var_NS <= COMP_LOOP_C_636;
      WHEN COMP_LOOP_C_636 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000110011");
        state_var_NS <= COMP_LOOP_C_637;
      WHEN COMP_LOOP_C_637 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000110100");
        state_var_NS <= COMP_LOOP_C_638;
      WHEN COMP_LOOP_C_638 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000110101");
        state_var_NS <= COMP_LOOP_C_639;
      WHEN COMP_LOOP_C_639 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000110110");
        state_var_NS <= COMP_LOOP_C_640;
      WHEN COMP_LOOP_C_640 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000110111");
        IF ( COMP_LOOP_C_640_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_641;
        END IF;
      WHEN COMP_LOOP_C_641 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000111000");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_0;
      WHEN COMP_LOOP_11_modExp_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000111001");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_1;
      WHEN COMP_LOOP_11_modExp_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000111010");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_2;
      WHEN COMP_LOOP_11_modExp_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000111011");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_3;
      WHEN COMP_LOOP_11_modExp_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000111100");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_4;
      WHEN COMP_LOOP_11_modExp_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000111101");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_5;
      WHEN COMP_LOOP_11_modExp_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000111110");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_6;
      WHEN COMP_LOOP_11_modExp_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000111111");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_7;
      WHEN COMP_LOOP_11_modExp_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001000000");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_8;
      WHEN COMP_LOOP_11_modExp_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001000001");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_9;
      WHEN COMP_LOOP_11_modExp_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001000010");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_10;
      WHEN COMP_LOOP_11_modExp_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001000011");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_11;
      WHEN COMP_LOOP_11_modExp_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001000100");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_12;
      WHEN COMP_LOOP_11_modExp_1_while_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001000101");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_13;
      WHEN COMP_LOOP_11_modExp_1_while_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001000110");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_14;
      WHEN COMP_LOOP_11_modExp_1_while_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001000111");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_15;
      WHEN COMP_LOOP_11_modExp_1_while_C_15 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001001000");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_16;
      WHEN COMP_LOOP_11_modExp_1_while_C_16 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001001001");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_17;
      WHEN COMP_LOOP_11_modExp_1_while_C_17 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001001010");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_18;
      WHEN COMP_LOOP_11_modExp_1_while_C_18 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001001011");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_19;
      WHEN COMP_LOOP_11_modExp_1_while_C_19 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001001100");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_20;
      WHEN COMP_LOOP_11_modExp_1_while_C_20 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001001101");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_21;
      WHEN COMP_LOOP_11_modExp_1_while_C_21 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001001110");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_22;
      WHEN COMP_LOOP_11_modExp_1_while_C_22 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001001111");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_23;
      WHEN COMP_LOOP_11_modExp_1_while_C_23 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001010000");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_24;
      WHEN COMP_LOOP_11_modExp_1_while_C_24 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001010001");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_25;
      WHEN COMP_LOOP_11_modExp_1_while_C_25 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001010010");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_26;
      WHEN COMP_LOOP_11_modExp_1_while_C_26 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001010011");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_27;
      WHEN COMP_LOOP_11_modExp_1_while_C_27 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001010100");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_28;
      WHEN COMP_LOOP_11_modExp_1_while_C_28 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001010101");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_29;
      WHEN COMP_LOOP_11_modExp_1_while_C_29 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001010110");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_30;
      WHEN COMP_LOOP_11_modExp_1_while_C_30 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001010111");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_31;
      WHEN COMP_LOOP_11_modExp_1_while_C_31 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001011000");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_32;
      WHEN COMP_LOOP_11_modExp_1_while_C_32 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001011001");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_33;
      WHEN COMP_LOOP_11_modExp_1_while_C_33 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001011010");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_34;
      WHEN COMP_LOOP_11_modExp_1_while_C_34 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001011011");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_35;
      WHEN COMP_LOOP_11_modExp_1_while_C_35 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001011100");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_36;
      WHEN COMP_LOOP_11_modExp_1_while_C_36 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001011101");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_37;
      WHEN COMP_LOOP_11_modExp_1_while_C_37 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001011110");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_38;
      WHEN COMP_LOOP_11_modExp_1_while_C_38 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001011111");
        IF ( COMP_LOOP_11_modExp_1_while_C_38_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_642;
        ELSE
          state_var_NS <= COMP_LOOP_11_modExp_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_642 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001100000");
        state_var_NS <= COMP_LOOP_C_643;
      WHEN COMP_LOOP_C_643 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001100001");
        state_var_NS <= COMP_LOOP_C_644;
      WHEN COMP_LOOP_C_644 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001100010");
        state_var_NS <= COMP_LOOP_C_645;
      WHEN COMP_LOOP_C_645 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001100011");
        state_var_NS <= COMP_LOOP_C_646;
      WHEN COMP_LOOP_C_646 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001100100");
        state_var_NS <= COMP_LOOP_C_647;
      WHEN COMP_LOOP_C_647 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001100101");
        state_var_NS <= COMP_LOOP_C_648;
      WHEN COMP_LOOP_C_648 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001100110");
        state_var_NS <= COMP_LOOP_C_649;
      WHEN COMP_LOOP_C_649 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001100111");
        state_var_NS <= COMP_LOOP_C_650;
      WHEN COMP_LOOP_C_650 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001101000");
        state_var_NS <= COMP_LOOP_C_651;
      WHEN COMP_LOOP_C_651 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001101001");
        state_var_NS <= COMP_LOOP_C_652;
      WHEN COMP_LOOP_C_652 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001101010");
        state_var_NS <= COMP_LOOP_C_653;
      WHEN COMP_LOOP_C_653 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001101011");
        state_var_NS <= COMP_LOOP_C_654;
      WHEN COMP_LOOP_C_654 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001101100");
        state_var_NS <= COMP_LOOP_C_655;
      WHEN COMP_LOOP_C_655 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001101101");
        state_var_NS <= COMP_LOOP_C_656;
      WHEN COMP_LOOP_C_656 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001101110");
        state_var_NS <= COMP_LOOP_C_657;
      WHEN COMP_LOOP_C_657 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001101111");
        state_var_NS <= COMP_LOOP_C_658;
      WHEN COMP_LOOP_C_658 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001110000");
        state_var_NS <= COMP_LOOP_C_659;
      WHEN COMP_LOOP_C_659 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001110001");
        state_var_NS <= COMP_LOOP_C_660;
      WHEN COMP_LOOP_C_660 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001110010");
        state_var_NS <= COMP_LOOP_C_661;
      WHEN COMP_LOOP_C_661 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001110011");
        state_var_NS <= COMP_LOOP_C_662;
      WHEN COMP_LOOP_C_662 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001110100");
        state_var_NS <= COMP_LOOP_C_663;
      WHEN COMP_LOOP_C_663 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001110101");
        state_var_NS <= COMP_LOOP_C_664;
      WHEN COMP_LOOP_C_664 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001110110");
        state_var_NS <= COMP_LOOP_C_665;
      WHEN COMP_LOOP_C_665 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001110111");
        state_var_NS <= COMP_LOOP_C_666;
      WHEN COMP_LOOP_C_666 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001111000");
        state_var_NS <= COMP_LOOP_C_667;
      WHEN COMP_LOOP_C_667 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001111001");
        state_var_NS <= COMP_LOOP_C_668;
      WHEN COMP_LOOP_C_668 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001111010");
        state_var_NS <= COMP_LOOP_C_669;
      WHEN COMP_LOOP_C_669 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001111011");
        state_var_NS <= COMP_LOOP_C_670;
      WHEN COMP_LOOP_C_670 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001111100");
        state_var_NS <= COMP_LOOP_C_671;
      WHEN COMP_LOOP_C_671 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001111101");
        state_var_NS <= COMP_LOOP_C_672;
      WHEN COMP_LOOP_C_672 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001111110");
        state_var_NS <= COMP_LOOP_C_673;
      WHEN COMP_LOOP_C_673 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001111111");
        state_var_NS <= COMP_LOOP_C_674;
      WHEN COMP_LOOP_C_674 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010000000");
        state_var_NS <= COMP_LOOP_C_675;
      WHEN COMP_LOOP_C_675 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010000001");
        state_var_NS <= COMP_LOOP_C_676;
      WHEN COMP_LOOP_C_676 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010000010");
        state_var_NS <= COMP_LOOP_C_677;
      WHEN COMP_LOOP_C_677 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010000011");
        state_var_NS <= COMP_LOOP_C_678;
      WHEN COMP_LOOP_C_678 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010000100");
        state_var_NS <= COMP_LOOP_C_679;
      WHEN COMP_LOOP_C_679 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010000101");
        state_var_NS <= COMP_LOOP_C_680;
      WHEN COMP_LOOP_C_680 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010000110");
        state_var_NS <= COMP_LOOP_C_681;
      WHEN COMP_LOOP_C_681 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010000111");
        state_var_NS <= COMP_LOOP_C_682;
      WHEN COMP_LOOP_C_682 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010001000");
        state_var_NS <= COMP_LOOP_C_683;
      WHEN COMP_LOOP_C_683 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010001001");
        state_var_NS <= COMP_LOOP_C_684;
      WHEN COMP_LOOP_C_684 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010001010");
        state_var_NS <= COMP_LOOP_C_685;
      WHEN COMP_LOOP_C_685 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010001011");
        state_var_NS <= COMP_LOOP_C_686;
      WHEN COMP_LOOP_C_686 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010001100");
        state_var_NS <= COMP_LOOP_C_687;
      WHEN COMP_LOOP_C_687 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010001101");
        state_var_NS <= COMP_LOOP_C_688;
      WHEN COMP_LOOP_C_688 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010001110");
        state_var_NS <= COMP_LOOP_C_689;
      WHEN COMP_LOOP_C_689 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010001111");
        state_var_NS <= COMP_LOOP_C_690;
      WHEN COMP_LOOP_C_690 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010010000");
        state_var_NS <= COMP_LOOP_C_691;
      WHEN COMP_LOOP_C_691 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010010001");
        state_var_NS <= COMP_LOOP_C_692;
      WHEN COMP_LOOP_C_692 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010010010");
        state_var_NS <= COMP_LOOP_C_693;
      WHEN COMP_LOOP_C_693 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010010011");
        state_var_NS <= COMP_LOOP_C_694;
      WHEN COMP_LOOP_C_694 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010010100");
        state_var_NS <= COMP_LOOP_C_695;
      WHEN COMP_LOOP_C_695 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010010101");
        state_var_NS <= COMP_LOOP_C_696;
      WHEN COMP_LOOP_C_696 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010010110");
        state_var_NS <= COMP_LOOP_C_697;
      WHEN COMP_LOOP_C_697 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010010111");
        state_var_NS <= COMP_LOOP_C_698;
      WHEN COMP_LOOP_C_698 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010011000");
        state_var_NS <= COMP_LOOP_C_699;
      WHEN COMP_LOOP_C_699 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010011001");
        state_var_NS <= COMP_LOOP_C_700;
      WHEN COMP_LOOP_C_700 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010011010");
        state_var_NS <= COMP_LOOP_C_701;
      WHEN COMP_LOOP_C_701 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010011011");
        state_var_NS <= COMP_LOOP_C_702;
      WHEN COMP_LOOP_C_702 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010011100");
        state_var_NS <= COMP_LOOP_C_703;
      WHEN COMP_LOOP_C_703 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010011101");
        state_var_NS <= COMP_LOOP_C_704;
      WHEN COMP_LOOP_C_704 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010011110");
        IF ( COMP_LOOP_C_704_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_705;
        END IF;
      WHEN COMP_LOOP_C_705 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010011111");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_0;
      WHEN COMP_LOOP_12_modExp_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010100000");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_1;
      WHEN COMP_LOOP_12_modExp_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010100001");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_2;
      WHEN COMP_LOOP_12_modExp_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010100010");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_3;
      WHEN COMP_LOOP_12_modExp_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010100011");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_4;
      WHEN COMP_LOOP_12_modExp_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010100100");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_5;
      WHEN COMP_LOOP_12_modExp_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010100101");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_6;
      WHEN COMP_LOOP_12_modExp_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010100110");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_7;
      WHEN COMP_LOOP_12_modExp_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010100111");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_8;
      WHEN COMP_LOOP_12_modExp_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010101000");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_9;
      WHEN COMP_LOOP_12_modExp_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010101001");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_10;
      WHEN COMP_LOOP_12_modExp_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010101010");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_11;
      WHEN COMP_LOOP_12_modExp_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010101011");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_12;
      WHEN COMP_LOOP_12_modExp_1_while_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010101100");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_13;
      WHEN COMP_LOOP_12_modExp_1_while_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010101101");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_14;
      WHEN COMP_LOOP_12_modExp_1_while_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010101110");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_15;
      WHEN COMP_LOOP_12_modExp_1_while_C_15 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010101111");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_16;
      WHEN COMP_LOOP_12_modExp_1_while_C_16 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010110000");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_17;
      WHEN COMP_LOOP_12_modExp_1_while_C_17 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010110001");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_18;
      WHEN COMP_LOOP_12_modExp_1_while_C_18 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010110010");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_19;
      WHEN COMP_LOOP_12_modExp_1_while_C_19 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010110011");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_20;
      WHEN COMP_LOOP_12_modExp_1_while_C_20 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010110100");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_21;
      WHEN COMP_LOOP_12_modExp_1_while_C_21 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010110101");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_22;
      WHEN COMP_LOOP_12_modExp_1_while_C_22 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010110110");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_23;
      WHEN COMP_LOOP_12_modExp_1_while_C_23 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010110111");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_24;
      WHEN COMP_LOOP_12_modExp_1_while_C_24 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010111000");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_25;
      WHEN COMP_LOOP_12_modExp_1_while_C_25 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010111001");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_26;
      WHEN COMP_LOOP_12_modExp_1_while_C_26 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010111010");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_27;
      WHEN COMP_LOOP_12_modExp_1_while_C_27 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010111011");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_28;
      WHEN COMP_LOOP_12_modExp_1_while_C_28 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010111100");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_29;
      WHEN COMP_LOOP_12_modExp_1_while_C_29 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010111101");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_30;
      WHEN COMP_LOOP_12_modExp_1_while_C_30 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010111110");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_31;
      WHEN COMP_LOOP_12_modExp_1_while_C_31 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010111111");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_32;
      WHEN COMP_LOOP_12_modExp_1_while_C_32 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011000000");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_33;
      WHEN COMP_LOOP_12_modExp_1_while_C_33 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011000001");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_34;
      WHEN COMP_LOOP_12_modExp_1_while_C_34 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011000010");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_35;
      WHEN COMP_LOOP_12_modExp_1_while_C_35 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011000011");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_36;
      WHEN COMP_LOOP_12_modExp_1_while_C_36 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011000100");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_37;
      WHEN COMP_LOOP_12_modExp_1_while_C_37 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011000101");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_38;
      WHEN COMP_LOOP_12_modExp_1_while_C_38 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011000110");
        IF ( COMP_LOOP_12_modExp_1_while_C_38_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_706;
        ELSE
          state_var_NS <= COMP_LOOP_12_modExp_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_706 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011000111");
        state_var_NS <= COMP_LOOP_C_707;
      WHEN COMP_LOOP_C_707 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011001000");
        state_var_NS <= COMP_LOOP_C_708;
      WHEN COMP_LOOP_C_708 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011001001");
        state_var_NS <= COMP_LOOP_C_709;
      WHEN COMP_LOOP_C_709 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011001010");
        state_var_NS <= COMP_LOOP_C_710;
      WHEN COMP_LOOP_C_710 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011001011");
        state_var_NS <= COMP_LOOP_C_711;
      WHEN COMP_LOOP_C_711 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011001100");
        state_var_NS <= COMP_LOOP_C_712;
      WHEN COMP_LOOP_C_712 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011001101");
        state_var_NS <= COMP_LOOP_C_713;
      WHEN COMP_LOOP_C_713 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011001110");
        state_var_NS <= COMP_LOOP_C_714;
      WHEN COMP_LOOP_C_714 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011001111");
        state_var_NS <= COMP_LOOP_C_715;
      WHEN COMP_LOOP_C_715 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011010000");
        state_var_NS <= COMP_LOOP_C_716;
      WHEN COMP_LOOP_C_716 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011010001");
        state_var_NS <= COMP_LOOP_C_717;
      WHEN COMP_LOOP_C_717 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011010010");
        state_var_NS <= COMP_LOOP_C_718;
      WHEN COMP_LOOP_C_718 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011010011");
        state_var_NS <= COMP_LOOP_C_719;
      WHEN COMP_LOOP_C_719 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011010100");
        state_var_NS <= COMP_LOOP_C_720;
      WHEN COMP_LOOP_C_720 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011010101");
        state_var_NS <= COMP_LOOP_C_721;
      WHEN COMP_LOOP_C_721 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011010110");
        state_var_NS <= COMP_LOOP_C_722;
      WHEN COMP_LOOP_C_722 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011010111");
        state_var_NS <= COMP_LOOP_C_723;
      WHEN COMP_LOOP_C_723 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011011000");
        state_var_NS <= COMP_LOOP_C_724;
      WHEN COMP_LOOP_C_724 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011011001");
        state_var_NS <= COMP_LOOP_C_725;
      WHEN COMP_LOOP_C_725 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011011010");
        state_var_NS <= COMP_LOOP_C_726;
      WHEN COMP_LOOP_C_726 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011011011");
        state_var_NS <= COMP_LOOP_C_727;
      WHEN COMP_LOOP_C_727 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011011100");
        state_var_NS <= COMP_LOOP_C_728;
      WHEN COMP_LOOP_C_728 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011011101");
        state_var_NS <= COMP_LOOP_C_729;
      WHEN COMP_LOOP_C_729 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011011110");
        state_var_NS <= COMP_LOOP_C_730;
      WHEN COMP_LOOP_C_730 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011011111");
        state_var_NS <= COMP_LOOP_C_731;
      WHEN COMP_LOOP_C_731 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011100000");
        state_var_NS <= COMP_LOOP_C_732;
      WHEN COMP_LOOP_C_732 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011100001");
        state_var_NS <= COMP_LOOP_C_733;
      WHEN COMP_LOOP_C_733 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011100010");
        state_var_NS <= COMP_LOOP_C_734;
      WHEN COMP_LOOP_C_734 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011100011");
        state_var_NS <= COMP_LOOP_C_735;
      WHEN COMP_LOOP_C_735 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011100100");
        state_var_NS <= COMP_LOOP_C_736;
      WHEN COMP_LOOP_C_736 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011100101");
        state_var_NS <= COMP_LOOP_C_737;
      WHEN COMP_LOOP_C_737 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011100110");
        state_var_NS <= COMP_LOOP_C_738;
      WHEN COMP_LOOP_C_738 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011100111");
        state_var_NS <= COMP_LOOP_C_739;
      WHEN COMP_LOOP_C_739 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011101000");
        state_var_NS <= COMP_LOOP_C_740;
      WHEN COMP_LOOP_C_740 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011101001");
        state_var_NS <= COMP_LOOP_C_741;
      WHEN COMP_LOOP_C_741 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011101010");
        state_var_NS <= COMP_LOOP_C_742;
      WHEN COMP_LOOP_C_742 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011101011");
        state_var_NS <= COMP_LOOP_C_743;
      WHEN COMP_LOOP_C_743 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011101100");
        state_var_NS <= COMP_LOOP_C_744;
      WHEN COMP_LOOP_C_744 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011101101");
        state_var_NS <= COMP_LOOP_C_745;
      WHEN COMP_LOOP_C_745 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011101110");
        state_var_NS <= COMP_LOOP_C_746;
      WHEN COMP_LOOP_C_746 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011101111");
        state_var_NS <= COMP_LOOP_C_747;
      WHEN COMP_LOOP_C_747 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011110000");
        state_var_NS <= COMP_LOOP_C_748;
      WHEN COMP_LOOP_C_748 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011110001");
        state_var_NS <= COMP_LOOP_C_749;
      WHEN COMP_LOOP_C_749 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011110010");
        state_var_NS <= COMP_LOOP_C_750;
      WHEN COMP_LOOP_C_750 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011110011");
        state_var_NS <= COMP_LOOP_C_751;
      WHEN COMP_LOOP_C_751 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011110100");
        state_var_NS <= COMP_LOOP_C_752;
      WHEN COMP_LOOP_C_752 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011110101");
        state_var_NS <= COMP_LOOP_C_753;
      WHEN COMP_LOOP_C_753 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011110110");
        state_var_NS <= COMP_LOOP_C_754;
      WHEN COMP_LOOP_C_754 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011110111");
        state_var_NS <= COMP_LOOP_C_755;
      WHEN COMP_LOOP_C_755 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011111000");
        state_var_NS <= COMP_LOOP_C_756;
      WHEN COMP_LOOP_C_756 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011111001");
        state_var_NS <= COMP_LOOP_C_757;
      WHEN COMP_LOOP_C_757 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011111010");
        state_var_NS <= COMP_LOOP_C_758;
      WHEN COMP_LOOP_C_758 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011111011");
        state_var_NS <= COMP_LOOP_C_759;
      WHEN COMP_LOOP_C_759 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011111100");
        state_var_NS <= COMP_LOOP_C_760;
      WHEN COMP_LOOP_C_760 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011111101");
        state_var_NS <= COMP_LOOP_C_761;
      WHEN COMP_LOOP_C_761 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011111110");
        state_var_NS <= COMP_LOOP_C_762;
      WHEN COMP_LOOP_C_762 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011111111");
        state_var_NS <= COMP_LOOP_C_763;
      WHEN COMP_LOOP_C_763 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100000000");
        state_var_NS <= COMP_LOOP_C_764;
      WHEN COMP_LOOP_C_764 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100000001");
        state_var_NS <= COMP_LOOP_C_765;
      WHEN COMP_LOOP_C_765 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100000010");
        state_var_NS <= COMP_LOOP_C_766;
      WHEN COMP_LOOP_C_766 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100000011");
        state_var_NS <= COMP_LOOP_C_767;
      WHEN COMP_LOOP_C_767 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100000100");
        state_var_NS <= COMP_LOOP_C_768;
      WHEN COMP_LOOP_C_768 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100000101");
        IF ( COMP_LOOP_C_768_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_769;
        END IF;
      WHEN COMP_LOOP_C_769 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100000110");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_0;
      WHEN COMP_LOOP_13_modExp_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100000111");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_1;
      WHEN COMP_LOOP_13_modExp_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100001000");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_2;
      WHEN COMP_LOOP_13_modExp_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100001001");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_3;
      WHEN COMP_LOOP_13_modExp_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100001010");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_4;
      WHEN COMP_LOOP_13_modExp_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100001011");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_5;
      WHEN COMP_LOOP_13_modExp_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100001100");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_6;
      WHEN COMP_LOOP_13_modExp_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100001101");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_7;
      WHEN COMP_LOOP_13_modExp_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100001110");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_8;
      WHEN COMP_LOOP_13_modExp_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100001111");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_9;
      WHEN COMP_LOOP_13_modExp_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100010000");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_10;
      WHEN COMP_LOOP_13_modExp_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100010001");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_11;
      WHEN COMP_LOOP_13_modExp_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100010010");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_12;
      WHEN COMP_LOOP_13_modExp_1_while_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100010011");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_13;
      WHEN COMP_LOOP_13_modExp_1_while_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100010100");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_14;
      WHEN COMP_LOOP_13_modExp_1_while_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100010101");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_15;
      WHEN COMP_LOOP_13_modExp_1_while_C_15 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100010110");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_16;
      WHEN COMP_LOOP_13_modExp_1_while_C_16 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100010111");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_17;
      WHEN COMP_LOOP_13_modExp_1_while_C_17 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100011000");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_18;
      WHEN COMP_LOOP_13_modExp_1_while_C_18 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100011001");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_19;
      WHEN COMP_LOOP_13_modExp_1_while_C_19 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100011010");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_20;
      WHEN COMP_LOOP_13_modExp_1_while_C_20 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100011011");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_21;
      WHEN COMP_LOOP_13_modExp_1_while_C_21 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100011100");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_22;
      WHEN COMP_LOOP_13_modExp_1_while_C_22 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100011101");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_23;
      WHEN COMP_LOOP_13_modExp_1_while_C_23 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100011110");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_24;
      WHEN COMP_LOOP_13_modExp_1_while_C_24 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100011111");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_25;
      WHEN COMP_LOOP_13_modExp_1_while_C_25 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100100000");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_26;
      WHEN COMP_LOOP_13_modExp_1_while_C_26 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100100001");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_27;
      WHEN COMP_LOOP_13_modExp_1_while_C_27 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100100010");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_28;
      WHEN COMP_LOOP_13_modExp_1_while_C_28 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100100011");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_29;
      WHEN COMP_LOOP_13_modExp_1_while_C_29 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100100100");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_30;
      WHEN COMP_LOOP_13_modExp_1_while_C_30 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100100101");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_31;
      WHEN COMP_LOOP_13_modExp_1_while_C_31 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100100110");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_32;
      WHEN COMP_LOOP_13_modExp_1_while_C_32 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100100111");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_33;
      WHEN COMP_LOOP_13_modExp_1_while_C_33 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100101000");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_34;
      WHEN COMP_LOOP_13_modExp_1_while_C_34 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100101001");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_35;
      WHEN COMP_LOOP_13_modExp_1_while_C_35 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100101010");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_36;
      WHEN COMP_LOOP_13_modExp_1_while_C_36 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100101011");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_37;
      WHEN COMP_LOOP_13_modExp_1_while_C_37 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100101100");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_38;
      WHEN COMP_LOOP_13_modExp_1_while_C_38 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100101101");
        IF ( COMP_LOOP_13_modExp_1_while_C_38_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_770;
        ELSE
          state_var_NS <= COMP_LOOP_13_modExp_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_770 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100101110");
        state_var_NS <= COMP_LOOP_C_771;
      WHEN COMP_LOOP_C_771 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100101111");
        state_var_NS <= COMP_LOOP_C_772;
      WHEN COMP_LOOP_C_772 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100110000");
        state_var_NS <= COMP_LOOP_C_773;
      WHEN COMP_LOOP_C_773 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100110001");
        state_var_NS <= COMP_LOOP_C_774;
      WHEN COMP_LOOP_C_774 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100110010");
        state_var_NS <= COMP_LOOP_C_775;
      WHEN COMP_LOOP_C_775 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100110011");
        state_var_NS <= COMP_LOOP_C_776;
      WHEN COMP_LOOP_C_776 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100110100");
        state_var_NS <= COMP_LOOP_C_777;
      WHEN COMP_LOOP_C_777 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100110101");
        state_var_NS <= COMP_LOOP_C_778;
      WHEN COMP_LOOP_C_778 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100110110");
        state_var_NS <= COMP_LOOP_C_779;
      WHEN COMP_LOOP_C_779 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100110111");
        state_var_NS <= COMP_LOOP_C_780;
      WHEN COMP_LOOP_C_780 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100111000");
        state_var_NS <= COMP_LOOP_C_781;
      WHEN COMP_LOOP_C_781 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100111001");
        state_var_NS <= COMP_LOOP_C_782;
      WHEN COMP_LOOP_C_782 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100111010");
        state_var_NS <= COMP_LOOP_C_783;
      WHEN COMP_LOOP_C_783 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100111011");
        state_var_NS <= COMP_LOOP_C_784;
      WHEN COMP_LOOP_C_784 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100111100");
        state_var_NS <= COMP_LOOP_C_785;
      WHEN COMP_LOOP_C_785 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100111101");
        state_var_NS <= COMP_LOOP_C_786;
      WHEN COMP_LOOP_C_786 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100111110");
        state_var_NS <= COMP_LOOP_C_787;
      WHEN COMP_LOOP_C_787 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100111111");
        state_var_NS <= COMP_LOOP_C_788;
      WHEN COMP_LOOP_C_788 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101000000");
        state_var_NS <= COMP_LOOP_C_789;
      WHEN COMP_LOOP_C_789 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101000001");
        state_var_NS <= COMP_LOOP_C_790;
      WHEN COMP_LOOP_C_790 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101000010");
        state_var_NS <= COMP_LOOP_C_791;
      WHEN COMP_LOOP_C_791 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101000011");
        state_var_NS <= COMP_LOOP_C_792;
      WHEN COMP_LOOP_C_792 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101000100");
        state_var_NS <= COMP_LOOP_C_793;
      WHEN COMP_LOOP_C_793 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101000101");
        state_var_NS <= COMP_LOOP_C_794;
      WHEN COMP_LOOP_C_794 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101000110");
        state_var_NS <= COMP_LOOP_C_795;
      WHEN COMP_LOOP_C_795 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101000111");
        state_var_NS <= COMP_LOOP_C_796;
      WHEN COMP_LOOP_C_796 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101001000");
        state_var_NS <= COMP_LOOP_C_797;
      WHEN COMP_LOOP_C_797 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101001001");
        state_var_NS <= COMP_LOOP_C_798;
      WHEN COMP_LOOP_C_798 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101001010");
        state_var_NS <= COMP_LOOP_C_799;
      WHEN COMP_LOOP_C_799 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101001011");
        state_var_NS <= COMP_LOOP_C_800;
      WHEN COMP_LOOP_C_800 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101001100");
        state_var_NS <= COMP_LOOP_C_801;
      WHEN COMP_LOOP_C_801 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101001101");
        state_var_NS <= COMP_LOOP_C_802;
      WHEN COMP_LOOP_C_802 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101001110");
        state_var_NS <= COMP_LOOP_C_803;
      WHEN COMP_LOOP_C_803 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101001111");
        state_var_NS <= COMP_LOOP_C_804;
      WHEN COMP_LOOP_C_804 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101010000");
        state_var_NS <= COMP_LOOP_C_805;
      WHEN COMP_LOOP_C_805 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101010001");
        state_var_NS <= COMP_LOOP_C_806;
      WHEN COMP_LOOP_C_806 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101010010");
        state_var_NS <= COMP_LOOP_C_807;
      WHEN COMP_LOOP_C_807 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101010011");
        state_var_NS <= COMP_LOOP_C_808;
      WHEN COMP_LOOP_C_808 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101010100");
        state_var_NS <= COMP_LOOP_C_809;
      WHEN COMP_LOOP_C_809 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101010101");
        state_var_NS <= COMP_LOOP_C_810;
      WHEN COMP_LOOP_C_810 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101010110");
        state_var_NS <= COMP_LOOP_C_811;
      WHEN COMP_LOOP_C_811 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101010111");
        state_var_NS <= COMP_LOOP_C_812;
      WHEN COMP_LOOP_C_812 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101011000");
        state_var_NS <= COMP_LOOP_C_813;
      WHEN COMP_LOOP_C_813 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101011001");
        state_var_NS <= COMP_LOOP_C_814;
      WHEN COMP_LOOP_C_814 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101011010");
        state_var_NS <= COMP_LOOP_C_815;
      WHEN COMP_LOOP_C_815 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101011011");
        state_var_NS <= COMP_LOOP_C_816;
      WHEN COMP_LOOP_C_816 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101011100");
        state_var_NS <= COMP_LOOP_C_817;
      WHEN COMP_LOOP_C_817 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101011101");
        state_var_NS <= COMP_LOOP_C_818;
      WHEN COMP_LOOP_C_818 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101011110");
        state_var_NS <= COMP_LOOP_C_819;
      WHEN COMP_LOOP_C_819 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101011111");
        state_var_NS <= COMP_LOOP_C_820;
      WHEN COMP_LOOP_C_820 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101100000");
        state_var_NS <= COMP_LOOP_C_821;
      WHEN COMP_LOOP_C_821 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101100001");
        state_var_NS <= COMP_LOOP_C_822;
      WHEN COMP_LOOP_C_822 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101100010");
        state_var_NS <= COMP_LOOP_C_823;
      WHEN COMP_LOOP_C_823 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101100011");
        state_var_NS <= COMP_LOOP_C_824;
      WHEN COMP_LOOP_C_824 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101100100");
        state_var_NS <= COMP_LOOP_C_825;
      WHEN COMP_LOOP_C_825 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101100101");
        state_var_NS <= COMP_LOOP_C_826;
      WHEN COMP_LOOP_C_826 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101100110");
        state_var_NS <= COMP_LOOP_C_827;
      WHEN COMP_LOOP_C_827 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101100111");
        state_var_NS <= COMP_LOOP_C_828;
      WHEN COMP_LOOP_C_828 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101101000");
        state_var_NS <= COMP_LOOP_C_829;
      WHEN COMP_LOOP_C_829 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101101001");
        state_var_NS <= COMP_LOOP_C_830;
      WHEN COMP_LOOP_C_830 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101101010");
        state_var_NS <= COMP_LOOP_C_831;
      WHEN COMP_LOOP_C_831 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101101011");
        state_var_NS <= COMP_LOOP_C_832;
      WHEN COMP_LOOP_C_832 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101101100");
        IF ( COMP_LOOP_C_832_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_833;
        END IF;
      WHEN COMP_LOOP_C_833 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101101101");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_0;
      WHEN COMP_LOOP_14_modExp_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101101110");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_1;
      WHEN COMP_LOOP_14_modExp_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101101111");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_2;
      WHEN COMP_LOOP_14_modExp_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101110000");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_3;
      WHEN COMP_LOOP_14_modExp_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101110001");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_4;
      WHEN COMP_LOOP_14_modExp_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101110010");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_5;
      WHEN COMP_LOOP_14_modExp_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101110011");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_6;
      WHEN COMP_LOOP_14_modExp_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101110100");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_7;
      WHEN COMP_LOOP_14_modExp_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101110101");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_8;
      WHEN COMP_LOOP_14_modExp_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101110110");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_9;
      WHEN COMP_LOOP_14_modExp_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101110111");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_10;
      WHEN COMP_LOOP_14_modExp_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101111000");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_11;
      WHEN COMP_LOOP_14_modExp_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101111001");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_12;
      WHEN COMP_LOOP_14_modExp_1_while_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101111010");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_13;
      WHEN COMP_LOOP_14_modExp_1_while_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101111011");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_14;
      WHEN COMP_LOOP_14_modExp_1_while_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101111100");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_15;
      WHEN COMP_LOOP_14_modExp_1_while_C_15 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101111101");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_16;
      WHEN COMP_LOOP_14_modExp_1_while_C_16 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101111110");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_17;
      WHEN COMP_LOOP_14_modExp_1_while_C_17 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101111111");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_18;
      WHEN COMP_LOOP_14_modExp_1_while_C_18 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110000000");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_19;
      WHEN COMP_LOOP_14_modExp_1_while_C_19 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110000001");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_20;
      WHEN COMP_LOOP_14_modExp_1_while_C_20 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110000010");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_21;
      WHEN COMP_LOOP_14_modExp_1_while_C_21 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110000011");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_22;
      WHEN COMP_LOOP_14_modExp_1_while_C_22 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110000100");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_23;
      WHEN COMP_LOOP_14_modExp_1_while_C_23 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110000101");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_24;
      WHEN COMP_LOOP_14_modExp_1_while_C_24 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110000110");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_25;
      WHEN COMP_LOOP_14_modExp_1_while_C_25 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110000111");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_26;
      WHEN COMP_LOOP_14_modExp_1_while_C_26 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110001000");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_27;
      WHEN COMP_LOOP_14_modExp_1_while_C_27 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110001001");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_28;
      WHEN COMP_LOOP_14_modExp_1_while_C_28 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110001010");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_29;
      WHEN COMP_LOOP_14_modExp_1_while_C_29 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110001011");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_30;
      WHEN COMP_LOOP_14_modExp_1_while_C_30 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110001100");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_31;
      WHEN COMP_LOOP_14_modExp_1_while_C_31 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110001101");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_32;
      WHEN COMP_LOOP_14_modExp_1_while_C_32 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110001110");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_33;
      WHEN COMP_LOOP_14_modExp_1_while_C_33 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110001111");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_34;
      WHEN COMP_LOOP_14_modExp_1_while_C_34 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110010000");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_35;
      WHEN COMP_LOOP_14_modExp_1_while_C_35 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110010001");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_36;
      WHEN COMP_LOOP_14_modExp_1_while_C_36 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110010010");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_37;
      WHEN COMP_LOOP_14_modExp_1_while_C_37 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110010011");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_38;
      WHEN COMP_LOOP_14_modExp_1_while_C_38 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110010100");
        IF ( COMP_LOOP_14_modExp_1_while_C_38_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_834;
        ELSE
          state_var_NS <= COMP_LOOP_14_modExp_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_834 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110010101");
        state_var_NS <= COMP_LOOP_C_835;
      WHEN COMP_LOOP_C_835 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110010110");
        state_var_NS <= COMP_LOOP_C_836;
      WHEN COMP_LOOP_C_836 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110010111");
        state_var_NS <= COMP_LOOP_C_837;
      WHEN COMP_LOOP_C_837 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110011000");
        state_var_NS <= COMP_LOOP_C_838;
      WHEN COMP_LOOP_C_838 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110011001");
        state_var_NS <= COMP_LOOP_C_839;
      WHEN COMP_LOOP_C_839 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110011010");
        state_var_NS <= COMP_LOOP_C_840;
      WHEN COMP_LOOP_C_840 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110011011");
        state_var_NS <= COMP_LOOP_C_841;
      WHEN COMP_LOOP_C_841 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110011100");
        state_var_NS <= COMP_LOOP_C_842;
      WHEN COMP_LOOP_C_842 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110011101");
        state_var_NS <= COMP_LOOP_C_843;
      WHEN COMP_LOOP_C_843 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110011110");
        state_var_NS <= COMP_LOOP_C_844;
      WHEN COMP_LOOP_C_844 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110011111");
        state_var_NS <= COMP_LOOP_C_845;
      WHEN COMP_LOOP_C_845 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110100000");
        state_var_NS <= COMP_LOOP_C_846;
      WHEN COMP_LOOP_C_846 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110100001");
        state_var_NS <= COMP_LOOP_C_847;
      WHEN COMP_LOOP_C_847 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110100010");
        state_var_NS <= COMP_LOOP_C_848;
      WHEN COMP_LOOP_C_848 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110100011");
        state_var_NS <= COMP_LOOP_C_849;
      WHEN COMP_LOOP_C_849 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110100100");
        state_var_NS <= COMP_LOOP_C_850;
      WHEN COMP_LOOP_C_850 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110100101");
        state_var_NS <= COMP_LOOP_C_851;
      WHEN COMP_LOOP_C_851 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110100110");
        state_var_NS <= COMP_LOOP_C_852;
      WHEN COMP_LOOP_C_852 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110100111");
        state_var_NS <= COMP_LOOP_C_853;
      WHEN COMP_LOOP_C_853 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110101000");
        state_var_NS <= COMP_LOOP_C_854;
      WHEN COMP_LOOP_C_854 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110101001");
        state_var_NS <= COMP_LOOP_C_855;
      WHEN COMP_LOOP_C_855 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110101010");
        state_var_NS <= COMP_LOOP_C_856;
      WHEN COMP_LOOP_C_856 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110101011");
        state_var_NS <= COMP_LOOP_C_857;
      WHEN COMP_LOOP_C_857 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110101100");
        state_var_NS <= COMP_LOOP_C_858;
      WHEN COMP_LOOP_C_858 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110101101");
        state_var_NS <= COMP_LOOP_C_859;
      WHEN COMP_LOOP_C_859 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110101110");
        state_var_NS <= COMP_LOOP_C_860;
      WHEN COMP_LOOP_C_860 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110101111");
        state_var_NS <= COMP_LOOP_C_861;
      WHEN COMP_LOOP_C_861 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110110000");
        state_var_NS <= COMP_LOOP_C_862;
      WHEN COMP_LOOP_C_862 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110110001");
        state_var_NS <= COMP_LOOP_C_863;
      WHEN COMP_LOOP_C_863 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110110010");
        state_var_NS <= COMP_LOOP_C_864;
      WHEN COMP_LOOP_C_864 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110110011");
        state_var_NS <= COMP_LOOP_C_865;
      WHEN COMP_LOOP_C_865 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110110100");
        state_var_NS <= COMP_LOOP_C_866;
      WHEN COMP_LOOP_C_866 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110110101");
        state_var_NS <= COMP_LOOP_C_867;
      WHEN COMP_LOOP_C_867 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110110110");
        state_var_NS <= COMP_LOOP_C_868;
      WHEN COMP_LOOP_C_868 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110110111");
        state_var_NS <= COMP_LOOP_C_869;
      WHEN COMP_LOOP_C_869 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110111000");
        state_var_NS <= COMP_LOOP_C_870;
      WHEN COMP_LOOP_C_870 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110111001");
        state_var_NS <= COMP_LOOP_C_871;
      WHEN COMP_LOOP_C_871 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110111010");
        state_var_NS <= COMP_LOOP_C_872;
      WHEN COMP_LOOP_C_872 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110111011");
        state_var_NS <= COMP_LOOP_C_873;
      WHEN COMP_LOOP_C_873 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110111100");
        state_var_NS <= COMP_LOOP_C_874;
      WHEN COMP_LOOP_C_874 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110111101");
        state_var_NS <= COMP_LOOP_C_875;
      WHEN COMP_LOOP_C_875 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110111110");
        state_var_NS <= COMP_LOOP_C_876;
      WHEN COMP_LOOP_C_876 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110111111");
        state_var_NS <= COMP_LOOP_C_877;
      WHEN COMP_LOOP_C_877 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111000000");
        state_var_NS <= COMP_LOOP_C_878;
      WHEN COMP_LOOP_C_878 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111000001");
        state_var_NS <= COMP_LOOP_C_879;
      WHEN COMP_LOOP_C_879 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111000010");
        state_var_NS <= COMP_LOOP_C_880;
      WHEN COMP_LOOP_C_880 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111000011");
        state_var_NS <= COMP_LOOP_C_881;
      WHEN COMP_LOOP_C_881 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111000100");
        state_var_NS <= COMP_LOOP_C_882;
      WHEN COMP_LOOP_C_882 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111000101");
        state_var_NS <= COMP_LOOP_C_883;
      WHEN COMP_LOOP_C_883 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111000110");
        state_var_NS <= COMP_LOOP_C_884;
      WHEN COMP_LOOP_C_884 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111000111");
        state_var_NS <= COMP_LOOP_C_885;
      WHEN COMP_LOOP_C_885 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111001000");
        state_var_NS <= COMP_LOOP_C_886;
      WHEN COMP_LOOP_C_886 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111001001");
        state_var_NS <= COMP_LOOP_C_887;
      WHEN COMP_LOOP_C_887 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111001010");
        state_var_NS <= COMP_LOOP_C_888;
      WHEN COMP_LOOP_C_888 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111001011");
        state_var_NS <= COMP_LOOP_C_889;
      WHEN COMP_LOOP_C_889 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111001100");
        state_var_NS <= COMP_LOOP_C_890;
      WHEN COMP_LOOP_C_890 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111001101");
        state_var_NS <= COMP_LOOP_C_891;
      WHEN COMP_LOOP_C_891 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111001110");
        state_var_NS <= COMP_LOOP_C_892;
      WHEN COMP_LOOP_C_892 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111001111");
        state_var_NS <= COMP_LOOP_C_893;
      WHEN COMP_LOOP_C_893 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111010000");
        state_var_NS <= COMP_LOOP_C_894;
      WHEN COMP_LOOP_C_894 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111010001");
        state_var_NS <= COMP_LOOP_C_895;
      WHEN COMP_LOOP_C_895 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111010010");
        state_var_NS <= COMP_LOOP_C_896;
      WHEN COMP_LOOP_C_896 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111010011");
        IF ( COMP_LOOP_C_896_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_897;
        END IF;
      WHEN COMP_LOOP_C_897 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111010100");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_0;
      WHEN COMP_LOOP_15_modExp_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111010101");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_1;
      WHEN COMP_LOOP_15_modExp_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111010110");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_2;
      WHEN COMP_LOOP_15_modExp_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111010111");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_3;
      WHEN COMP_LOOP_15_modExp_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111011000");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_4;
      WHEN COMP_LOOP_15_modExp_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111011001");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_5;
      WHEN COMP_LOOP_15_modExp_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111011010");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_6;
      WHEN COMP_LOOP_15_modExp_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111011011");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_7;
      WHEN COMP_LOOP_15_modExp_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111011100");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_8;
      WHEN COMP_LOOP_15_modExp_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111011101");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_9;
      WHEN COMP_LOOP_15_modExp_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111011110");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_10;
      WHEN COMP_LOOP_15_modExp_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111011111");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_11;
      WHEN COMP_LOOP_15_modExp_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111100000");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_12;
      WHEN COMP_LOOP_15_modExp_1_while_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111100001");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_13;
      WHEN COMP_LOOP_15_modExp_1_while_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111100010");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_14;
      WHEN COMP_LOOP_15_modExp_1_while_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111100011");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_15;
      WHEN COMP_LOOP_15_modExp_1_while_C_15 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111100100");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_16;
      WHEN COMP_LOOP_15_modExp_1_while_C_16 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111100101");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_17;
      WHEN COMP_LOOP_15_modExp_1_while_C_17 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111100110");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_18;
      WHEN COMP_LOOP_15_modExp_1_while_C_18 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111100111");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_19;
      WHEN COMP_LOOP_15_modExp_1_while_C_19 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111101000");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_20;
      WHEN COMP_LOOP_15_modExp_1_while_C_20 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111101001");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_21;
      WHEN COMP_LOOP_15_modExp_1_while_C_21 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111101010");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_22;
      WHEN COMP_LOOP_15_modExp_1_while_C_22 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111101011");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_23;
      WHEN COMP_LOOP_15_modExp_1_while_C_23 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111101100");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_24;
      WHEN COMP_LOOP_15_modExp_1_while_C_24 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111101101");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_25;
      WHEN COMP_LOOP_15_modExp_1_while_C_25 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111101110");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_26;
      WHEN COMP_LOOP_15_modExp_1_while_C_26 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111101111");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_27;
      WHEN COMP_LOOP_15_modExp_1_while_C_27 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111110000");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_28;
      WHEN COMP_LOOP_15_modExp_1_while_C_28 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111110001");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_29;
      WHEN COMP_LOOP_15_modExp_1_while_C_29 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111110010");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_30;
      WHEN COMP_LOOP_15_modExp_1_while_C_30 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111110011");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_31;
      WHEN COMP_LOOP_15_modExp_1_while_C_31 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111110100");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_32;
      WHEN COMP_LOOP_15_modExp_1_while_C_32 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111110101");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_33;
      WHEN COMP_LOOP_15_modExp_1_while_C_33 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111110110");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_34;
      WHEN COMP_LOOP_15_modExp_1_while_C_34 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111110111");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_35;
      WHEN COMP_LOOP_15_modExp_1_while_C_35 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111111000");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_36;
      WHEN COMP_LOOP_15_modExp_1_while_C_36 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111111001");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_37;
      WHEN COMP_LOOP_15_modExp_1_while_C_37 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111111010");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_38;
      WHEN COMP_LOOP_15_modExp_1_while_C_38 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111111011");
        IF ( COMP_LOOP_15_modExp_1_while_C_38_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_898;
        ELSE
          state_var_NS <= COMP_LOOP_15_modExp_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_898 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111111100");
        state_var_NS <= COMP_LOOP_C_899;
      WHEN COMP_LOOP_C_899 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111111101");
        state_var_NS <= COMP_LOOP_C_900;
      WHEN COMP_LOOP_C_900 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111111110");
        state_var_NS <= COMP_LOOP_C_901;
      WHEN COMP_LOOP_C_901 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111111111");
        state_var_NS <= COMP_LOOP_C_902;
      WHEN COMP_LOOP_C_902 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000000000");
        state_var_NS <= COMP_LOOP_C_903;
      WHEN COMP_LOOP_C_903 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000000001");
        state_var_NS <= COMP_LOOP_C_904;
      WHEN COMP_LOOP_C_904 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000000010");
        state_var_NS <= COMP_LOOP_C_905;
      WHEN COMP_LOOP_C_905 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000000011");
        state_var_NS <= COMP_LOOP_C_906;
      WHEN COMP_LOOP_C_906 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000000100");
        state_var_NS <= COMP_LOOP_C_907;
      WHEN COMP_LOOP_C_907 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000000101");
        state_var_NS <= COMP_LOOP_C_908;
      WHEN COMP_LOOP_C_908 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000000110");
        state_var_NS <= COMP_LOOP_C_909;
      WHEN COMP_LOOP_C_909 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000000111");
        state_var_NS <= COMP_LOOP_C_910;
      WHEN COMP_LOOP_C_910 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000001000");
        state_var_NS <= COMP_LOOP_C_911;
      WHEN COMP_LOOP_C_911 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000001001");
        state_var_NS <= COMP_LOOP_C_912;
      WHEN COMP_LOOP_C_912 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000001010");
        state_var_NS <= COMP_LOOP_C_913;
      WHEN COMP_LOOP_C_913 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000001011");
        state_var_NS <= COMP_LOOP_C_914;
      WHEN COMP_LOOP_C_914 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000001100");
        state_var_NS <= COMP_LOOP_C_915;
      WHEN COMP_LOOP_C_915 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000001101");
        state_var_NS <= COMP_LOOP_C_916;
      WHEN COMP_LOOP_C_916 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000001110");
        state_var_NS <= COMP_LOOP_C_917;
      WHEN COMP_LOOP_C_917 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000001111");
        state_var_NS <= COMP_LOOP_C_918;
      WHEN COMP_LOOP_C_918 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000010000");
        state_var_NS <= COMP_LOOP_C_919;
      WHEN COMP_LOOP_C_919 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000010001");
        state_var_NS <= COMP_LOOP_C_920;
      WHEN COMP_LOOP_C_920 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000010010");
        state_var_NS <= COMP_LOOP_C_921;
      WHEN COMP_LOOP_C_921 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000010011");
        state_var_NS <= COMP_LOOP_C_922;
      WHEN COMP_LOOP_C_922 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000010100");
        state_var_NS <= COMP_LOOP_C_923;
      WHEN COMP_LOOP_C_923 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000010101");
        state_var_NS <= COMP_LOOP_C_924;
      WHEN COMP_LOOP_C_924 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000010110");
        state_var_NS <= COMP_LOOP_C_925;
      WHEN COMP_LOOP_C_925 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000010111");
        state_var_NS <= COMP_LOOP_C_926;
      WHEN COMP_LOOP_C_926 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000011000");
        state_var_NS <= COMP_LOOP_C_927;
      WHEN COMP_LOOP_C_927 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000011001");
        state_var_NS <= COMP_LOOP_C_928;
      WHEN COMP_LOOP_C_928 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000011010");
        state_var_NS <= COMP_LOOP_C_929;
      WHEN COMP_LOOP_C_929 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000011011");
        state_var_NS <= COMP_LOOP_C_930;
      WHEN COMP_LOOP_C_930 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000011100");
        state_var_NS <= COMP_LOOP_C_931;
      WHEN COMP_LOOP_C_931 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000011101");
        state_var_NS <= COMP_LOOP_C_932;
      WHEN COMP_LOOP_C_932 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000011110");
        state_var_NS <= COMP_LOOP_C_933;
      WHEN COMP_LOOP_C_933 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000011111");
        state_var_NS <= COMP_LOOP_C_934;
      WHEN COMP_LOOP_C_934 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000100000");
        state_var_NS <= COMP_LOOP_C_935;
      WHEN COMP_LOOP_C_935 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000100001");
        state_var_NS <= COMP_LOOP_C_936;
      WHEN COMP_LOOP_C_936 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000100010");
        state_var_NS <= COMP_LOOP_C_937;
      WHEN COMP_LOOP_C_937 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000100011");
        state_var_NS <= COMP_LOOP_C_938;
      WHEN COMP_LOOP_C_938 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000100100");
        state_var_NS <= COMP_LOOP_C_939;
      WHEN COMP_LOOP_C_939 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000100101");
        state_var_NS <= COMP_LOOP_C_940;
      WHEN COMP_LOOP_C_940 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000100110");
        state_var_NS <= COMP_LOOP_C_941;
      WHEN COMP_LOOP_C_941 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000100111");
        state_var_NS <= COMP_LOOP_C_942;
      WHEN COMP_LOOP_C_942 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000101000");
        state_var_NS <= COMP_LOOP_C_943;
      WHEN COMP_LOOP_C_943 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000101001");
        state_var_NS <= COMP_LOOP_C_944;
      WHEN COMP_LOOP_C_944 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000101010");
        state_var_NS <= COMP_LOOP_C_945;
      WHEN COMP_LOOP_C_945 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000101011");
        state_var_NS <= COMP_LOOP_C_946;
      WHEN COMP_LOOP_C_946 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000101100");
        state_var_NS <= COMP_LOOP_C_947;
      WHEN COMP_LOOP_C_947 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000101101");
        state_var_NS <= COMP_LOOP_C_948;
      WHEN COMP_LOOP_C_948 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000101110");
        state_var_NS <= COMP_LOOP_C_949;
      WHEN COMP_LOOP_C_949 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000101111");
        state_var_NS <= COMP_LOOP_C_950;
      WHEN COMP_LOOP_C_950 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000110000");
        state_var_NS <= COMP_LOOP_C_951;
      WHEN COMP_LOOP_C_951 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000110001");
        state_var_NS <= COMP_LOOP_C_952;
      WHEN COMP_LOOP_C_952 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000110010");
        state_var_NS <= COMP_LOOP_C_953;
      WHEN COMP_LOOP_C_953 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000110011");
        state_var_NS <= COMP_LOOP_C_954;
      WHEN COMP_LOOP_C_954 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000110100");
        state_var_NS <= COMP_LOOP_C_955;
      WHEN COMP_LOOP_C_955 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000110101");
        state_var_NS <= COMP_LOOP_C_956;
      WHEN COMP_LOOP_C_956 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000110110");
        state_var_NS <= COMP_LOOP_C_957;
      WHEN COMP_LOOP_C_957 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000110111");
        state_var_NS <= COMP_LOOP_C_958;
      WHEN COMP_LOOP_C_958 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000111000");
        state_var_NS <= COMP_LOOP_C_959;
      WHEN COMP_LOOP_C_959 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000111001");
        state_var_NS <= COMP_LOOP_C_960;
      WHEN COMP_LOOP_C_960 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000111010");
        IF ( COMP_LOOP_C_960_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_961;
        END IF;
      WHEN COMP_LOOP_C_961 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000111011");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_0;
      WHEN COMP_LOOP_16_modExp_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000111100");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_1;
      WHEN COMP_LOOP_16_modExp_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000111101");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_2;
      WHEN COMP_LOOP_16_modExp_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000111110");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_3;
      WHEN COMP_LOOP_16_modExp_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000111111");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_4;
      WHEN COMP_LOOP_16_modExp_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001000000");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_5;
      WHEN COMP_LOOP_16_modExp_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001000001");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_6;
      WHEN COMP_LOOP_16_modExp_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001000010");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_7;
      WHEN COMP_LOOP_16_modExp_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001000011");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_8;
      WHEN COMP_LOOP_16_modExp_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001000100");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_9;
      WHEN COMP_LOOP_16_modExp_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001000101");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_10;
      WHEN COMP_LOOP_16_modExp_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001000110");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_11;
      WHEN COMP_LOOP_16_modExp_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001000111");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_12;
      WHEN COMP_LOOP_16_modExp_1_while_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001001000");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_13;
      WHEN COMP_LOOP_16_modExp_1_while_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001001001");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_14;
      WHEN COMP_LOOP_16_modExp_1_while_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001001010");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_15;
      WHEN COMP_LOOP_16_modExp_1_while_C_15 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001001011");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_16;
      WHEN COMP_LOOP_16_modExp_1_while_C_16 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001001100");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_17;
      WHEN COMP_LOOP_16_modExp_1_while_C_17 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001001101");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_18;
      WHEN COMP_LOOP_16_modExp_1_while_C_18 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001001110");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_19;
      WHEN COMP_LOOP_16_modExp_1_while_C_19 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001001111");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_20;
      WHEN COMP_LOOP_16_modExp_1_while_C_20 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001010000");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_21;
      WHEN COMP_LOOP_16_modExp_1_while_C_21 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001010001");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_22;
      WHEN COMP_LOOP_16_modExp_1_while_C_22 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001010010");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_23;
      WHEN COMP_LOOP_16_modExp_1_while_C_23 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001010011");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_24;
      WHEN COMP_LOOP_16_modExp_1_while_C_24 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001010100");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_25;
      WHEN COMP_LOOP_16_modExp_1_while_C_25 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001010101");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_26;
      WHEN COMP_LOOP_16_modExp_1_while_C_26 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001010110");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_27;
      WHEN COMP_LOOP_16_modExp_1_while_C_27 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001010111");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_28;
      WHEN COMP_LOOP_16_modExp_1_while_C_28 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001011000");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_29;
      WHEN COMP_LOOP_16_modExp_1_while_C_29 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001011001");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_30;
      WHEN COMP_LOOP_16_modExp_1_while_C_30 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001011010");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_31;
      WHEN COMP_LOOP_16_modExp_1_while_C_31 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001011011");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_32;
      WHEN COMP_LOOP_16_modExp_1_while_C_32 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001011100");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_33;
      WHEN COMP_LOOP_16_modExp_1_while_C_33 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001011101");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_34;
      WHEN COMP_LOOP_16_modExp_1_while_C_34 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001011110");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_35;
      WHEN COMP_LOOP_16_modExp_1_while_C_35 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001011111");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_36;
      WHEN COMP_LOOP_16_modExp_1_while_C_36 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001100000");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_37;
      WHEN COMP_LOOP_16_modExp_1_while_C_37 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001100001");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_38;
      WHEN COMP_LOOP_16_modExp_1_while_C_38 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001100010");
        IF ( COMP_LOOP_16_modExp_1_while_C_38_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_962;
        ELSE
          state_var_NS <= COMP_LOOP_16_modExp_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_962 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001100011");
        state_var_NS <= COMP_LOOP_C_963;
      WHEN COMP_LOOP_C_963 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001100100");
        state_var_NS <= COMP_LOOP_C_964;
      WHEN COMP_LOOP_C_964 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001100101");
        state_var_NS <= COMP_LOOP_C_965;
      WHEN COMP_LOOP_C_965 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001100110");
        state_var_NS <= COMP_LOOP_C_966;
      WHEN COMP_LOOP_C_966 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001100111");
        state_var_NS <= COMP_LOOP_C_967;
      WHEN COMP_LOOP_C_967 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001101000");
        state_var_NS <= COMP_LOOP_C_968;
      WHEN COMP_LOOP_C_968 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001101001");
        state_var_NS <= COMP_LOOP_C_969;
      WHEN COMP_LOOP_C_969 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001101010");
        state_var_NS <= COMP_LOOP_C_970;
      WHEN COMP_LOOP_C_970 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001101011");
        state_var_NS <= COMP_LOOP_C_971;
      WHEN COMP_LOOP_C_971 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001101100");
        state_var_NS <= COMP_LOOP_C_972;
      WHEN COMP_LOOP_C_972 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001101101");
        state_var_NS <= COMP_LOOP_C_973;
      WHEN COMP_LOOP_C_973 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001101110");
        state_var_NS <= COMP_LOOP_C_974;
      WHEN COMP_LOOP_C_974 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001101111");
        state_var_NS <= COMP_LOOP_C_975;
      WHEN COMP_LOOP_C_975 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001110000");
        state_var_NS <= COMP_LOOP_C_976;
      WHEN COMP_LOOP_C_976 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001110001");
        state_var_NS <= COMP_LOOP_C_977;
      WHEN COMP_LOOP_C_977 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001110010");
        state_var_NS <= COMP_LOOP_C_978;
      WHEN COMP_LOOP_C_978 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001110011");
        state_var_NS <= COMP_LOOP_C_979;
      WHEN COMP_LOOP_C_979 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001110100");
        state_var_NS <= COMP_LOOP_C_980;
      WHEN COMP_LOOP_C_980 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001110101");
        state_var_NS <= COMP_LOOP_C_981;
      WHEN COMP_LOOP_C_981 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001110110");
        state_var_NS <= COMP_LOOP_C_982;
      WHEN COMP_LOOP_C_982 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001110111");
        state_var_NS <= COMP_LOOP_C_983;
      WHEN COMP_LOOP_C_983 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001111000");
        state_var_NS <= COMP_LOOP_C_984;
      WHEN COMP_LOOP_C_984 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001111001");
        state_var_NS <= COMP_LOOP_C_985;
      WHEN COMP_LOOP_C_985 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001111010");
        state_var_NS <= COMP_LOOP_C_986;
      WHEN COMP_LOOP_C_986 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001111011");
        state_var_NS <= COMP_LOOP_C_987;
      WHEN COMP_LOOP_C_987 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001111100");
        state_var_NS <= COMP_LOOP_C_988;
      WHEN COMP_LOOP_C_988 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001111101");
        state_var_NS <= COMP_LOOP_C_989;
      WHEN COMP_LOOP_C_989 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001111110");
        state_var_NS <= COMP_LOOP_C_990;
      WHEN COMP_LOOP_C_990 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001111111");
        state_var_NS <= COMP_LOOP_C_991;
      WHEN COMP_LOOP_C_991 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11010000000");
        state_var_NS <= COMP_LOOP_C_992;
      WHEN COMP_LOOP_C_992 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11010000001");
        state_var_NS <= COMP_LOOP_C_993;
      WHEN COMP_LOOP_C_993 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11010000010");
        state_var_NS <= COMP_LOOP_C_994;
      WHEN COMP_LOOP_C_994 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11010000011");
        state_var_NS <= COMP_LOOP_C_995;
      WHEN COMP_LOOP_C_995 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11010000100");
        state_var_NS <= COMP_LOOP_C_996;
      WHEN COMP_LOOP_C_996 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11010000101");
        state_var_NS <= COMP_LOOP_C_997;
      WHEN COMP_LOOP_C_997 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11010000110");
        state_var_NS <= COMP_LOOP_C_998;
      WHEN COMP_LOOP_C_998 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11010000111");
        state_var_NS <= COMP_LOOP_C_999;
      WHEN COMP_LOOP_C_999 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11010001000");
        state_var_NS <= COMP_LOOP_C_1000;
      WHEN COMP_LOOP_C_1000 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11010001001");
        state_var_NS <= COMP_LOOP_C_1001;
      WHEN COMP_LOOP_C_1001 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11010001010");
        state_var_NS <= COMP_LOOP_C_1002;
      WHEN COMP_LOOP_C_1002 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11010001011");
        state_var_NS <= COMP_LOOP_C_1003;
      WHEN COMP_LOOP_C_1003 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11010001100");
        state_var_NS <= COMP_LOOP_C_1004;
      WHEN COMP_LOOP_C_1004 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11010001101");
        state_var_NS <= COMP_LOOP_C_1005;
      WHEN COMP_LOOP_C_1005 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11010001110");
        state_var_NS <= COMP_LOOP_C_1006;
      WHEN COMP_LOOP_C_1006 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11010001111");
        state_var_NS <= COMP_LOOP_C_1007;
      WHEN COMP_LOOP_C_1007 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11010010000");
        state_var_NS <= COMP_LOOP_C_1008;
      WHEN COMP_LOOP_C_1008 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11010010001");
        state_var_NS <= COMP_LOOP_C_1009;
      WHEN COMP_LOOP_C_1009 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11010010010");
        state_var_NS <= COMP_LOOP_C_1010;
      WHEN COMP_LOOP_C_1010 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11010010011");
        state_var_NS <= COMP_LOOP_C_1011;
      WHEN COMP_LOOP_C_1011 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11010010100");
        state_var_NS <= COMP_LOOP_C_1012;
      WHEN COMP_LOOP_C_1012 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11010010101");
        state_var_NS <= COMP_LOOP_C_1013;
      WHEN COMP_LOOP_C_1013 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11010010110");
        state_var_NS <= COMP_LOOP_C_1014;
      WHEN COMP_LOOP_C_1014 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11010010111");
        state_var_NS <= COMP_LOOP_C_1015;
      WHEN COMP_LOOP_C_1015 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11010011000");
        state_var_NS <= COMP_LOOP_C_1016;
      WHEN COMP_LOOP_C_1016 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11010011001");
        state_var_NS <= COMP_LOOP_C_1017;
      WHEN COMP_LOOP_C_1017 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11010011010");
        state_var_NS <= COMP_LOOP_C_1018;
      WHEN COMP_LOOP_C_1018 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11010011011");
        state_var_NS <= COMP_LOOP_C_1019;
      WHEN COMP_LOOP_C_1019 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11010011100");
        state_var_NS <= COMP_LOOP_C_1020;
      WHEN COMP_LOOP_C_1020 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11010011101");
        state_var_NS <= COMP_LOOP_C_1021;
      WHEN COMP_LOOP_C_1021 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11010011110");
        state_var_NS <= COMP_LOOP_C_1022;
      WHEN COMP_LOOP_C_1022 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11010011111");
        state_var_NS <= COMP_LOOP_C_1023;
      WHEN COMP_LOOP_C_1023 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11010100000");
        state_var_NS <= COMP_LOOP_C_1024;
      WHEN COMP_LOOP_C_1024 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11010100001");
        IF ( COMP_LOOP_C_1024_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_0;
        END IF;
      WHEN VEC_LOOP_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11010100010");
        IF ( VEC_LOOP_C_0_tr0 = '1' ) THEN
          state_var_NS <= STAGE_LOOP_C_9;
        ELSE
          state_var_NS <= COMP_LOOP_C_0;
        END IF;
      WHEN STAGE_LOOP_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11010100011");
        IF ( STAGE_LOOP_C_9_tr0 = '1' ) THEN
          state_var_NS <= main_C_1;
        ELSE
          state_var_NS <= STAGE_LOOP_C_0;
        END IF;
      WHEN main_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11010100100");
        state_var_NS <= main_C_0;
      -- main_C_0
      WHEN OTHERS =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000");
        state_var_NS <= STAGE_LOOP_C_0;
    END CASE;
  END PROCESS inPlaceNTT_DIT_core_core_fsm_1;

  inPlaceNTT_DIT_core_core_fsm_1_REG : PROCESS (clk)
  BEGIN
    IF clk'event AND ( clk = '1' ) THEN
      IF ( rst = '1' ) THEN
        state_var <= main_C_0;
      ELSE
        state_var <= state_var_NS;
      END IF;
    END IF;
  END PROCESS inPlaceNTT_DIT_core_core_fsm_1_REG;

END v44;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT_core
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT_core IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    vec_rsc_triosy_0_0_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_1_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_2_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_3_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_4_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_5_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_6_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_7_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_8_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_9_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_10_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_11_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_12_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_13_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_14_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_15_lz : OUT STD_LOGIC;
    p_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    p_rsc_triosy_lz : OUT STD_LOGIC;
    r_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    r_rsc_triosy_lz : OUT STD_LOGIC;
    vec_rsc_0_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_1_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_2_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_3_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_4_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_5_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_6_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_7_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_8_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_9_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_10_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_11_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_12_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_13_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_14_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_15_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_0_i_adra_d_pff : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    vec_rsc_0_0_i_da_d_pff : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_0_i_wea_d_pff : OUT STD_LOGIC;
    vec_rsc_0_1_i_wea_d_pff : OUT STD_LOGIC;
    vec_rsc_0_2_i_wea_d_pff : OUT STD_LOGIC;
    vec_rsc_0_3_i_wea_d_pff : OUT STD_LOGIC;
    vec_rsc_0_4_i_wea_d_pff : OUT STD_LOGIC;
    vec_rsc_0_5_i_wea_d_pff : OUT STD_LOGIC;
    vec_rsc_0_6_i_wea_d_pff : OUT STD_LOGIC;
    vec_rsc_0_7_i_wea_d_pff : OUT STD_LOGIC;
    vec_rsc_0_8_i_wea_d_pff : OUT STD_LOGIC;
    vec_rsc_0_9_i_wea_d_pff : OUT STD_LOGIC;
    vec_rsc_0_10_i_wea_d_pff : OUT STD_LOGIC;
    vec_rsc_0_11_i_wea_d_pff : OUT STD_LOGIC;
    vec_rsc_0_12_i_wea_d_pff : OUT STD_LOGIC;
    vec_rsc_0_13_i_wea_d_pff : OUT STD_LOGIC;
    vec_rsc_0_14_i_wea_d_pff : OUT STD_LOGIC;
    vec_rsc_0_15_i_wea_d_pff : OUT STD_LOGIC
  );
END inPlaceNTT_DIT_core;

ARCHITECTURE v44 OF inPlaceNTT_DIT_core IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL p_rsci_idat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL r_rsci_idat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL modulo_result_rem_cmp_a : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL modulo_result_rem_cmp_b : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL modulo_result_rem_cmp_z : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL operator_66_true_div_cmp_a : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL operator_66_true_div_cmp_z : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL operator_66_true_div_cmp_b_9_0 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL fsm_output : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL nor_tmp_4 : STD_LOGIC;
  SIGNAL mux_tmp_14 : STD_LOGIC;
  SIGNAL not_tmp_39 : STD_LOGIC;
  SIGNAL or_tmp_68 : STD_LOGIC;
  SIGNAL not_tmp_49 : STD_LOGIC;
  SIGNAL mux_tmp_119 : STD_LOGIC;
  SIGNAL or_tmp_88 : STD_LOGIC;
  SIGNAL mux_tmp_130 : STD_LOGIC;
  SIGNAL mux_tmp_131 : STD_LOGIC;
  SIGNAL or_tmp_93 : STD_LOGIC;
  SIGNAL nand_tmp_4 : STD_LOGIC;
  SIGNAL or_tmp_94 : STD_LOGIC;
  SIGNAL mux_tmp_139 : STD_LOGIC;
  SIGNAL mux_tmp_141 : STD_LOGIC;
  SIGNAL or_tmp_96 : STD_LOGIC;
  SIGNAL mux_tmp_165 : STD_LOGIC;
  SIGNAL or_tmp_104 : STD_LOGIC;
  SIGNAL mux_tmp_214 : STD_LOGIC;
  SIGNAL mux_tmp_215 : STD_LOGIC;
  SIGNAL nand_tmp_7 : STD_LOGIC;
  SIGNAL mux_tmp_227 : STD_LOGIC;
  SIGNAL nor_tmp_23 : STD_LOGIC;
  SIGNAL mux_tmp_228 : STD_LOGIC;
  SIGNAL mux_tmp_231 : STD_LOGIC;
  SIGNAL mux_tmp_236 : STD_LOGIC;
  SIGNAL or_tmp_114 : STD_LOGIC;
  SIGNAL and_dcpl_1 : STD_LOGIC;
  SIGNAL and_dcpl_2 : STD_LOGIC;
  SIGNAL and_dcpl_4 : STD_LOGIC;
  SIGNAL and_dcpl_5 : STD_LOGIC;
  SIGNAL and_dcpl_6 : STD_LOGIC;
  SIGNAL not_tmp_90 : STD_LOGIC;
  SIGNAL or_tmp_167 : STD_LOGIC;
  SIGNAL nor_tmp_48 : STD_LOGIC;
  SIGNAL or_tmp_222 : STD_LOGIC;
  SIGNAL not_tmp_133 : STD_LOGIC;
  SIGNAL nor_tmp_82 : STD_LOGIC;
  SIGNAL or_tmp_258 : STD_LOGIC;
  SIGNAL and_dcpl_19 : STD_LOGIC;
  SIGNAL and_dcpl_26 : STD_LOGIC;
  SIGNAL and_dcpl_27 : STD_LOGIC;
  SIGNAL and_dcpl_33 : STD_LOGIC;
  SIGNAL and_dcpl_34 : STD_LOGIC;
  SIGNAL and_dcpl_39 : STD_LOGIC;
  SIGNAL and_dcpl_40 : STD_LOGIC;
  SIGNAL and_dcpl_44 : STD_LOGIC;
  SIGNAL and_dcpl_48 : STD_LOGIC;
  SIGNAL and_dcpl_55 : STD_LOGIC;
  SIGNAL and_dcpl_59 : STD_LOGIC;
  SIGNAL not_tmp_208 : STD_LOGIC;
  SIGNAL and_dcpl_87 : STD_LOGIC;
  SIGNAL and_dcpl_88 : STD_LOGIC;
  SIGNAL and_dcpl_90 : STD_LOGIC;
  SIGNAL and_dcpl_91 : STD_LOGIC;
  SIGNAL and_dcpl_92 : STD_LOGIC;
  SIGNAL and_dcpl_93 : STD_LOGIC;
  SIGNAL and_dcpl_98 : STD_LOGIC;
  SIGNAL and_dcpl_103 : STD_LOGIC;
  SIGNAL and_dcpl_107 : STD_LOGIC;
  SIGNAL and_dcpl_108 : STD_LOGIC;
  SIGNAL and_dcpl_109 : STD_LOGIC;
  SIGNAL and_dcpl_111 : STD_LOGIC;
  SIGNAL and_dcpl_112 : STD_LOGIC;
  SIGNAL and_dcpl_113 : STD_LOGIC;
  SIGNAL and_dcpl_114 : STD_LOGIC;
  SIGNAL and_dcpl_115 : STD_LOGIC;
  SIGNAL and_dcpl_117 : STD_LOGIC;
  SIGNAL and_dcpl_118 : STD_LOGIC;
  SIGNAL or_tmp_453 : STD_LOGIC;
  SIGNAL mux_tmp_1082 : STD_LOGIC;
  SIGNAL and_dcpl_126 : STD_LOGIC;
  SIGNAL and_dcpl_127 : STD_LOGIC;
  SIGNAL and_dcpl_130 : STD_LOGIC;
  SIGNAL and_dcpl_135 : STD_LOGIC;
  SIGNAL and_dcpl_136 : STD_LOGIC;
  SIGNAL and_dcpl_139 : STD_LOGIC;
  SIGNAL and_dcpl_140 : STD_LOGIC;
  SIGNAL and_dcpl_144 : STD_LOGIC;
  SIGNAL and_dcpl_146 : STD_LOGIC;
  SIGNAL and_dcpl_147 : STD_LOGIC;
  SIGNAL and_dcpl_149 : STD_LOGIC;
  SIGNAL and_dcpl_152 : STD_LOGIC;
  SIGNAL and_dcpl_153 : STD_LOGIC;
  SIGNAL and_dcpl_155 : STD_LOGIC;
  SIGNAL and_dcpl_162 : STD_LOGIC;
  SIGNAL and_dcpl_164 : STD_LOGIC;
  SIGNAL and_dcpl_170 : STD_LOGIC;
  SIGNAL and_dcpl_171 : STD_LOGIC;
  SIGNAL and_dcpl_177 : STD_LOGIC;
  SIGNAL and_dcpl_178 : STD_LOGIC;
  SIGNAL and_dcpl_185 : STD_LOGIC;
  SIGNAL and_dcpl_189 : STD_LOGIC;
  SIGNAL and_dcpl_191 : STD_LOGIC;
  SIGNAL and_dcpl_196 : STD_LOGIC;
  SIGNAL and_dcpl_197 : STD_LOGIC;
  SIGNAL and_dcpl_202 : STD_LOGIC;
  SIGNAL and_dcpl_208 : STD_LOGIC;
  SIGNAL and_dcpl_209 : STD_LOGIC;
  SIGNAL and_dcpl_211 : STD_LOGIC;
  SIGNAL and_dcpl_219 : STD_LOGIC;
  SIGNAL and_dcpl_224 : STD_LOGIC;
  SIGNAL and_dcpl_226 : STD_LOGIC;
  SIGNAL and_dcpl_231 : STD_LOGIC;
  SIGNAL not_tmp_248 : STD_LOGIC;
  SIGNAL mux_tmp_1116 : STD_LOGIC;
  SIGNAL or_tmp_532 : STD_LOGIC;
  SIGNAL not_tmp_253 : STD_LOGIC;
  SIGNAL mux_tmp_1180 : STD_LOGIC;
  SIGNAL or_tmp_643 : STD_LOGIC;
  SIGNAL mux_tmp_1244 : STD_LOGIC;
  SIGNAL or_tmp_756 : STD_LOGIC;
  SIGNAL mux_tmp_1308 : STD_LOGIC;
  SIGNAL or_tmp_866 : STD_LOGIC;
  SIGNAL mux_tmp_1372 : STD_LOGIC;
  SIGNAL or_tmp_974 : STD_LOGIC;
  SIGNAL mux_tmp_1436 : STD_LOGIC;
  SIGNAL or_tmp_1085 : STD_LOGIC;
  SIGNAL mux_tmp_1500 : STD_LOGIC;
  SIGNAL or_tmp_1198 : STD_LOGIC;
  SIGNAL mux_tmp_1564 : STD_LOGIC;
  SIGNAL or_tmp_1308 : STD_LOGIC;
  SIGNAL not_tmp_318 : STD_LOGIC;
  SIGNAL mux_tmp_1628 : STD_LOGIC;
  SIGNAL or_tmp_1416 : STD_LOGIC;
  SIGNAL mux_tmp_1692 : STD_LOGIC;
  SIGNAL or_tmp_1527 : STD_LOGIC;
  SIGNAL mux_tmp_1756 : STD_LOGIC;
  SIGNAL or_tmp_1640 : STD_LOGIC;
  SIGNAL mux_tmp_1820 : STD_LOGIC;
  SIGNAL or_tmp_1750 : STD_LOGIC;
  SIGNAL not_tmp_357 : STD_LOGIC;
  SIGNAL mux_tmp_1884 : STD_LOGIC;
  SIGNAL or_tmp_1858 : STD_LOGIC;
  SIGNAL mux_tmp_1948 : STD_LOGIC;
  SIGNAL or_tmp_1969 : STD_LOGIC;
  SIGNAL not_tmp_377 : STD_LOGIC;
  SIGNAL mux_tmp_2012 : STD_LOGIC;
  SIGNAL or_tmp_2082 : STD_LOGIC;
  SIGNAL not_tmp_387 : STD_LOGIC;
  SIGNAL mux_tmp_2076 : STD_LOGIC;
  SIGNAL not_tmp_390 : STD_LOGIC;
  SIGNAL or_tmp_2192 : STD_LOGIC;
  SIGNAL nor_tmp_265 : STD_LOGIC;
  SIGNAL and_dcpl_235 : STD_LOGIC;
  SIGNAL and_dcpl_236 : STD_LOGIC;
  SIGNAL and_dcpl_237 : STD_LOGIC;
  SIGNAL or_tmp_2274 : STD_LOGIC;
  SIGNAL or_tmp_2276 : STD_LOGIC;
  SIGNAL or_tmp_2277 : STD_LOGIC;
  SIGNAL or_tmp_2280 : STD_LOGIC;
  SIGNAL or_tmp_2281 : STD_LOGIC;
  SIGNAL mux_tmp_2159 : STD_LOGIC;
  SIGNAL or_tmp_2294 : STD_LOGIC;
  SIGNAL mux_tmp_2172 : STD_LOGIC;
  SIGNAL or_tmp_2297 : STD_LOGIC;
  SIGNAL mux_tmp_2176 : STD_LOGIC;
  SIGNAL mux_tmp_2178 : STD_LOGIC;
  SIGNAL or_tmp_2302 : STD_LOGIC;
  SIGNAL mux_tmp_2235 : STD_LOGIC;
  SIGNAL mux_tmp_2241 : STD_LOGIC;
  SIGNAL or_tmp_2340 : STD_LOGIC;
  SIGNAL or_tmp_2341 : STD_LOGIC;
  SIGNAL mux_tmp_2262 : STD_LOGIC;
  SIGNAL mux_tmp_2287 : STD_LOGIC;
  SIGNAL mux_tmp_2289 : STD_LOGIC;
  SIGNAL mux_tmp_2293 : STD_LOGIC;
  SIGNAL or_tmp_2360 : STD_LOGIC;
  SIGNAL mux_tmp_2311 : STD_LOGIC;
  SIGNAL or_tmp_2376 : STD_LOGIC;
  SIGNAL or_tmp_2389 : STD_LOGIC;
  SIGNAL mux_tmp_2347 : STD_LOGIC;
  SIGNAL or_tmp_2390 : STD_LOGIC;
  SIGNAL mux_tmp_2348 : STD_LOGIC;
  SIGNAL mux_tmp_2350 : STD_LOGIC;
  SIGNAL not_tmp_431 : STD_LOGIC;
  SIGNAL mux_tmp_2353 : STD_LOGIC;
  SIGNAL or_tmp_2393 : STD_LOGIC;
  SIGNAL or_tmp_2394 : STD_LOGIC;
  SIGNAL mux_tmp_2355 : STD_LOGIC;
  SIGNAL mux_tmp_2356 : STD_LOGIC;
  SIGNAL or_tmp_2396 : STD_LOGIC;
  SIGNAL or_tmp_2397 : STD_LOGIC;
  SIGNAL or_tmp_2399 : STD_LOGIC;
  SIGNAL mux_tmp_2359 : STD_LOGIC;
  SIGNAL mux_tmp_2361 : STD_LOGIC;
  SIGNAL mux_tmp_2363 : STD_LOGIC;
  SIGNAL mux_tmp_2364 : STD_LOGIC;
  SIGNAL or_tmp_2404 : STD_LOGIC;
  SIGNAL mux_tmp_2365 : STD_LOGIC;
  SIGNAL nand_tmp_54 : STD_LOGIC;
  SIGNAL or_tmp_2405 : STD_LOGIC;
  SIGNAL mux_tmp_2369 : STD_LOGIC;
  SIGNAL mux_tmp_2370 : STD_LOGIC;
  SIGNAL mux_tmp_2371 : STD_LOGIC;
  SIGNAL mux_tmp_2376 : STD_LOGIC;
  SIGNAL mux_tmp_2377 : STD_LOGIC;
  SIGNAL mux_tmp_2378 : STD_LOGIC;
  SIGNAL mux_tmp_2382 : STD_LOGIC;
  SIGNAL or_tmp_2407 : STD_LOGIC;
  SIGNAL mux_tmp_2386 : STD_LOGIC;
  SIGNAL mux_tmp_2389 : STD_LOGIC;
  SIGNAL mux_tmp_2424 : STD_LOGIC;
  SIGNAL not_tmp_441 : STD_LOGIC;
  SIGNAL or_tmp_2436 : STD_LOGIC;
  SIGNAL not_tmp_446 : STD_LOGIC;
  SIGNAL and_dcpl_241 : STD_LOGIC;
  SIGNAL and_dcpl_245 : STD_LOGIC;
  SIGNAL and_dcpl_247 : STD_LOGIC;
  SIGNAL nor_tmp_324 : STD_LOGIC;
  SIGNAL or_tmp_2474 : STD_LOGIC;
  SIGNAL mux_tmp_2640 : STD_LOGIC;
  SIGNAL mux_tmp_2659 : STD_LOGIC;
  SIGNAL and_dcpl_256 : STD_LOGIC;
  SIGNAL mux_tmp_2669 : STD_LOGIC;
  SIGNAL mux_tmp_2672 : STD_LOGIC;
  SIGNAL mux_tmp_2675 : STD_LOGIC;
  SIGNAL not_tmp_500 : STD_LOGIC;
  SIGNAL mux_tmp_2682 : STD_LOGIC;
  SIGNAL mux_tmp_2690 : STD_LOGIC;
  SIGNAL mux_tmp_2691 : STD_LOGIC;
  SIGNAL mux_tmp_2693 : STD_LOGIC;
  SIGNAL or_tmp_2603 : STD_LOGIC;
  SIGNAL or_tmp_2604 : STD_LOGIC;
  SIGNAL mux_tmp_2700 : STD_LOGIC;
  SIGNAL mux_tmp_2702 : STD_LOGIC;
  SIGNAL mux_tmp_2703 : STD_LOGIC;
  SIGNAL mux_tmp_2706 : STD_LOGIC;
  SIGNAL mux_tmp_2709 : STD_LOGIC;
  SIGNAL mux_tmp_2715 : STD_LOGIC;
  SIGNAL mux_tmp_2736 : STD_LOGIC;
  SIGNAL and_dcpl_257 : STD_LOGIC;
  SIGNAL and_dcpl_260 : STD_LOGIC;
  SIGNAL and_dcpl_262 : STD_LOGIC;
  SIGNAL and_dcpl_270 : STD_LOGIC;
  SIGNAL and_dcpl_278 : STD_LOGIC;
  SIGNAL and_dcpl_280 : STD_LOGIC;
  SIGNAL mux_tmp_2745 : STD_LOGIC;
  SIGNAL mux_tmp_2760 : STD_LOGIC;
  SIGNAL or_tmp_2651 : STD_LOGIC;
  SIGNAL or_tmp_2682 : STD_LOGIC;
  SIGNAL or_tmp_2683 : STD_LOGIC;
  SIGNAL or_tmp_2690 : STD_LOGIC;
  SIGNAL or_tmp_2693 : STD_LOGIC;
  SIGNAL or_tmp_2696 : STD_LOGIC;
  SIGNAL or_tmp_2697 : STD_LOGIC;
  SIGNAL mux_tmp_2796 : STD_LOGIC;
  SIGNAL or_tmp_2701 : STD_LOGIC;
  SIGNAL or_tmp_2703 : STD_LOGIC;
  SIGNAL or_tmp_2704 : STD_LOGIC;
  SIGNAL or_tmp_2706 : STD_LOGIC;
  SIGNAL or_tmp_2709 : STD_LOGIC;
  SIGNAL or_tmp_2714 : STD_LOGIC;
  SIGNAL mux_tmp_2841 : STD_LOGIC;
  SIGNAL or_tmp_2729 : STD_LOGIC;
  SIGNAL or_tmp_2731 : STD_LOGIC;
  SIGNAL mux_tmp_2843 : STD_LOGIC;
  SIGNAL mux_tmp_2844 : STD_LOGIC;
  SIGNAL or_tmp_2734 : STD_LOGIC;
  SIGNAL mux_tmp_2848 : STD_LOGIC;
  SIGNAL mux_tmp_2850 : STD_LOGIC;
  SIGNAL or_tmp_2736 : STD_LOGIC;
  SIGNAL mux_tmp_2851 : STD_LOGIC;
  SIGNAL mux_tmp_2856 : STD_LOGIC;
  SIGNAL nand_tmp_67 : STD_LOGIC;
  SIGNAL mux_tmp_2862 : STD_LOGIC;
  SIGNAL mux_tmp_2863 : STD_LOGIC;
  SIGNAL or_tmp_2739 : STD_LOGIC;
  SIGNAL mux_tmp_2867 : STD_LOGIC;
  SIGNAL or_tmp_2740 : STD_LOGIC;
  SIGNAL mux_tmp_2876 : STD_LOGIC;
  SIGNAL mux_tmp_2878 : STD_LOGIC;
  SIGNAL mux_tmp_2879 : STD_LOGIC;
  SIGNAL or_tmp_2742 : STD_LOGIC;
  SIGNAL mux_tmp_2880 : STD_LOGIC;
  SIGNAL mux_tmp_2886 : STD_LOGIC;
  SIGNAL mux_tmp_2888 : STD_LOGIC;
  SIGNAL mux_tmp_2890 : STD_LOGIC;
  SIGNAL or_tmp_2743 : STD_LOGIC;
  SIGNAL nand_tmp_68 : STD_LOGIC;
  SIGNAL mux_tmp_2895 : STD_LOGIC;
  SIGNAL or_tmp_2745 : STD_LOGIC;
  SIGNAL or_tmp_2746 : STD_LOGIC;
  SIGNAL nand_tmp_69 : STD_LOGIC;
  SIGNAL mux_tmp_2906 : STD_LOGIC;
  SIGNAL mux_tmp_2910 : STD_LOGIC;
  SIGNAL nand_tmp_70 : STD_LOGIC;
  SIGNAL mux_tmp_2912 : STD_LOGIC;
  SIGNAL nand_tmp_71 : STD_LOGIC;
  SIGNAL mux_tmp_2916 : STD_LOGIC;
  SIGNAL mux_tmp_2920 : STD_LOGIC;
  SIGNAL or_tmp_2749 : STD_LOGIC;
  SIGNAL or_tmp_2774 : STD_LOGIC;
  SIGNAL mux_tmp_2996 : STD_LOGIC;
  SIGNAL not_tmp_557 : STD_LOGIC;
  SIGNAL nor_tmp_405 : STD_LOGIC;
  SIGNAL mux_tmp_3007 : STD_LOGIC;
  SIGNAL mux_tmp_3008 : STD_LOGIC;
  SIGNAL or_tmp_2791 : STD_LOGIC;
  SIGNAL mux_tmp_3014 : STD_LOGIC;
  SIGNAL or_tmp_2795 : STD_LOGIC;
  SIGNAL or_tmp_2802 : STD_LOGIC;
  SIGNAL or_tmp_2803 : STD_LOGIC;
  SIGNAL mux_tmp_3024 : STD_LOGIC;
  SIGNAL mux_tmp_3032 : STD_LOGIC;
  SIGNAL mux_tmp_3049 : STD_LOGIC;
  SIGNAL or_tmp_2814 : STD_LOGIC;
  SIGNAL nor_tmp_410 : STD_LOGIC;
  SIGNAL and_dcpl_304 : STD_LOGIC;
  SIGNAL not_tmp_619 : STD_LOGIC;
  SIGNAL mux_tmp_3329 : STD_LOGIC;
  SIGNAL nor_tmp_457 : STD_LOGIC;
  SIGNAL mux_tmp_3341 : STD_LOGIC;
  SIGNAL mux_tmp_3343 : STD_LOGIC;
  SIGNAL mux_tmp_3361 : STD_LOGIC;
  SIGNAL or_tmp_2988 : STD_LOGIC;
  SIGNAL mux_tmp_3378 : STD_LOGIC;
  SIGNAL not_tmp_647 : STD_LOGIC;
  SIGNAL mux_tmp_3410 : STD_LOGIC;
  SIGNAL mux_tmp_3414 : STD_LOGIC;
  SIGNAL mux_tmp_3415 : STD_LOGIC;
  SIGNAL mux_tmp_3417 : STD_LOGIC;
  SIGNAL or_tmp_3023 : STD_LOGIC;
  SIGNAL mux_tmp_3418 : STD_LOGIC;
  SIGNAL mux_tmp_3420 : STD_LOGIC;
  SIGNAL mux_tmp_3421 : STD_LOGIC;
  SIGNAL mux_tmp_3423 : STD_LOGIC;
  SIGNAL mux_tmp_3424 : STD_LOGIC;
  SIGNAL mux_tmp_3425 : STD_LOGIC;
  SIGNAL not_tmp_663 : STD_LOGIC;
  SIGNAL mux_tmp_3429 : STD_LOGIC;
  SIGNAL mux_tmp_3432 : STD_LOGIC;
  SIGNAL mux_tmp_3434 : STD_LOGIC;
  SIGNAL mux_tmp_3435 : STD_LOGIC;
  SIGNAL not_tmp_665 : STD_LOGIC;
  SIGNAL mux_tmp_3453 : STD_LOGIC;
  SIGNAL mux_tmp_3456 : STD_LOGIC;
  SIGNAL mux_tmp_3457 : STD_LOGIC;
  SIGNAL mux_tmp_3458 : STD_LOGIC;
  SIGNAL mux_tmp_3459 : STD_LOGIC;
  SIGNAL not_tmp_672 : STD_LOGIC;
  SIGNAL mux_tmp_3463 : STD_LOGIC;
  SIGNAL mux_tmp_3464 : STD_LOGIC;
  SIGNAL mux_tmp_3472 : STD_LOGIC;
  SIGNAL mux_tmp_3473 : STD_LOGIC;
  SIGNAL mux_tmp_3474 : STD_LOGIC;
  SIGNAL mux_tmp_3477 : STD_LOGIC;
  SIGNAL mux_tmp_3481 : STD_LOGIC;
  SIGNAL mux_tmp_3491 : STD_LOGIC;
  SIGNAL not_tmp_688 : STD_LOGIC;
  SIGNAL or_tmp_3053 : STD_LOGIC;
  SIGNAL mux_tmp_3529 : STD_LOGIC;
  SIGNAL not_tmp_701 : STD_LOGIC;
  SIGNAL or_tmp_3095 : STD_LOGIC;
  SIGNAL mux_tmp_3547 : STD_LOGIC;
  SIGNAL mux_tmp_3551 : STD_LOGIC;
  SIGNAL mux_tmp_3574 : STD_LOGIC;
  SIGNAL mux_tmp_3576 : STD_LOGIC;
  SIGNAL mux_tmp_3577 : STD_LOGIC;
  SIGNAL mux_tmp_3618 : STD_LOGIC;
  SIGNAL or_tmp_3135 : STD_LOGIC;
  SIGNAL mux_tmp_3632 : STD_LOGIC;
  SIGNAL or_tmp_3176 : STD_LOGIC;
  SIGNAL or_tmp_3190 : STD_LOGIC;
  SIGNAL mux_tmp_3673 : STD_LOGIC;
  SIGNAL mux_tmp_3674 : STD_LOGIC;
  SIGNAL mux_tmp_3679 : STD_LOGIC;
  SIGNAL mux_tmp_3681 : STD_LOGIC;
  SIGNAL and_tmp_28 : STD_LOGIC;
  SIGNAL mux_tmp_3691 : STD_LOGIC;
  SIGNAL or_tmp_3224 : STD_LOGIC;
  SIGNAL mux_tmp_3698 : STD_LOGIC;
  SIGNAL mux_tmp_3701 : STD_LOGIC;
  SIGNAL mux_tmp_3705 : STD_LOGIC;
  SIGNAL mux_tmp_3720 : STD_LOGIC;
  SIGNAL mux_tmp_3724 : STD_LOGIC;
  SIGNAL mux_tmp_3736 : STD_LOGIC;
  SIGNAL mux_tmp_3737 : STD_LOGIC;
  SIGNAL mux_tmp_3739 : STD_LOGIC;
  SIGNAL mux_tmp_3753 : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_137_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_10_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_11_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_acc_1_cse_6_sva_1 : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL VEC_LOOP_j_sva_11_0 : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL COMP_LOOP_k_9_4_sva_4_0 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_acc_10_cse_12_1_1_sva : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_1_cse_14_sva : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_1_cse_2_sva : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_14_psp_sva : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_17_psp_sva : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_1_cse_6_sva : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_1_cse_10_sva : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_11_psp_sva : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_20_psp_sva : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_1_cse_4_sva : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_1_cse_sva : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_19_psp_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_16_psp_sva : STD_LOGIC_VECTOR (8 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_1_cse_8_sva : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_1_cse_12_sva : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_13_psp_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL tmp_10_lpi_4_dfm : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_1_cse_2_sva_1 : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL mux_2771_m1c : STD_LOGIC;
  SIGNAL and_279_m1c : STD_LOGIC;
  SIGNAL and_281_m1c : STD_LOGIC;
  SIGNAL and_284_m1c : STD_LOGIC;
  SIGNAL and_286_m1c : STD_LOGIC;
  SIGNAL and_288_m1c : STD_LOGIC;
  SIGNAL and_291_m1c : STD_LOGIC;
  SIGNAL and_292_m1c : STD_LOGIC;
  SIGNAL and_295_m1c : STD_LOGIC;
  SIGNAL and_297_m1c : STD_LOGIC;
  SIGNAL and_299_m1c : STD_LOGIC;
  SIGNAL and_302_m1c : STD_LOGIC;
  SIGNAL and_304_m1c : STD_LOGIC;
  SIGNAL and_307_m1c : STD_LOGIC;
  SIGNAL and_309_m1c : STD_LOGIC;
  SIGNAL and_311_m1c : STD_LOGIC;
  SIGNAL and_273_m1c : STD_LOGIC;
  SIGNAL nor_1445_cse : STD_LOGIC;
  SIGNAL mux_1157_cse : STD_LOGIC;
  SIGNAL nand_332_cse : STD_LOGIC;
  SIGNAL mux_1413_cse : STD_LOGIC;
  SIGNAL nand_324_cse : STD_LOGIC;
  SIGNAL mux_1669_cse : STD_LOGIC;
  SIGNAL mux_1925_cse : STD_LOGIC;
  SIGNAL reg_vec_rsc_triosy_0_15_obj_ld_cse : STD_LOGIC;
  SIGNAL and_527_cse : STD_LOGIC;
  SIGNAL or_2377_cse : STD_LOGIC;
  SIGNAL or_2368_cse : STD_LOGIC;
  SIGNAL and_529_cse : STD_LOGIC;
  SIGNAL and_526_cse : STD_LOGIC;
  SIGNAL or_3388_cse : STD_LOGIC;
  SIGNAL nor_758_cse : STD_LOGIC;
  SIGNAL nand_196_cse : STD_LOGIC;
  SIGNAL or_2419_cse : STD_LOGIC;
  SIGNAL nor_297_cse : STD_LOGIC;
  SIGNAL nor_303_cse : STD_LOGIC;
  SIGNAL mux_125_cse : STD_LOGIC;
  SIGNAL nand_356_cse : STD_LOGIC;
  SIGNAL or_491_cse : STD_LOGIC;
  SIGNAL nand_357_cse : STD_LOGIC;
  SIGNAL nand_358_cse : STD_LOGIC;
  SIGNAL or_2921_cse : STD_LOGIC;
  SIGNAL or_2918_cse : STD_LOGIC;
  SIGNAL and_536_cse : STD_LOGIC;
  SIGNAL nor_753_cse : STD_LOGIC;
  SIGNAL nand_159_cse : STD_LOGIC;
  SIGNAL or_2387_cse : STD_LOGIC;
  SIGNAL or_2912_cse : STD_LOGIC;
  SIGNAL mux_554_cse : STD_LOGIC;
  SIGNAL or_181_cse : STD_LOGIC;
  SIGNAL and_458_cse : STD_LOGIC;
  SIGNAL and_407_cse : STD_LOGIC;
  SIGNAL or_3039_cse : STD_LOGIC;
  SIGNAL and_459_cse : STD_LOGIC;
  SIGNAL or_2644_cse : STD_LOGIC;
  SIGNAL or_470_cse : STD_LOGIC;
  SIGNAL and_672_cse : STD_LOGIC;
  SIGNAL and_395_cse : STD_LOGIC;
  SIGNAL and_676_cse : STD_LOGIC;
  SIGNAL or_361_cse : STD_LOGIC;
  SIGNAL or_2414_cse : STD_LOGIC;
  SIGNAL or_3063_cse : STD_LOGIC;
  SIGNAL and_756_cse : STD_LOGIC;
  SIGNAL nand_142_cse : STD_LOGIC;
  SIGNAL and_366_cse : STD_LOGIC;
  SIGNAL and_350_cse : STD_LOGIC;
  SIGNAL or_3427_cse : STD_LOGIC;
  SIGNAL or_2991_cse : STD_LOGIC;
  SIGNAL nand_138_cse : STD_LOGIC;
  SIGNAL or_2407_cse : STD_LOGIC;
  SIGNAL or_2998_cse : STD_LOGIC;
  SIGNAL or_469_cse : STD_LOGIC;
  SIGNAL and_757_cse : STD_LOGIC;
  SIGNAL nor_609_cse : STD_LOGIC;
  SIGNAL or_352_cse : STD_LOGIC;
  SIGNAL and_404_cse : STD_LOGIC;
  SIGNAL and_707_cse : STD_LOGIC;
  SIGNAL or_259_cse : STD_LOGIC;
  SIGNAL nor_1580_cse : STD_LOGIC;
  SIGNAL or_586_cse : STD_LOGIC;
  SIGNAL or_591_cse : STD_LOGIC;
  SIGNAL nand_334_cse : STD_LOGIC;
  SIGNAL or_702_cse : STD_LOGIC;
  SIGNAL nor_209_cse : STD_LOGIC;
  SIGNAL nand_337_cse : STD_LOGIC;
  SIGNAL or_1028_cse : STD_LOGIC;
  SIGNAL nor_223_cse : STD_LOGIC;
  SIGNAL or_1470_cse : STD_LOGIC;
  SIGNAL nor_239_cse : STD_LOGIC;
  SIGNAL or_1912_cse : STD_LOGIC;
  SIGNAL and_564_cse : STD_LOGIC;
  SIGNAL mux_2926_cse : STD_LOGIC;
  SIGNAL mux_2486_cse : STD_LOGIC;
  SIGNAL or_2540_cse : STD_LOGIC;
  SIGNAL nor_694_cse : STD_LOGIC;
  SIGNAL or_70_cse : STD_LOGIC;
  SIGNAL or_56_cse : STD_LOGIC;
  SIGNAL nor_657_cse : STD_LOGIC;
  SIGNAL nand_367_cse : STD_LOGIC;
  SIGNAL or_2947_cse : STD_LOGIC;
  SIGNAL or_2905_cse : STD_LOGIC;
  SIGNAL or_3079_cse : STD_LOGIC;
  SIGNAL and_524_cse : STD_LOGIC;
  SIGNAL or_3074_cse : STD_LOGIC;
  SIGNAL nand_183_cse : STD_LOGIC;
  SIGNAL nor_667_cse : STD_LOGIC;
  SIGNAL or_163_cse : STD_LOGIC;
  SIGNAL or_3417_cse : STD_LOGIC;
  SIGNAL and_465_cse : STD_LOGIC;
  SIGNAL mux_1149_cse : STD_LOGIC;
  SIGNAL mux_1277_cse : STD_LOGIC;
  SIGNAL mux_1405_cse : STD_LOGIC;
  SIGNAL mux_1533_cse : STD_LOGIC;
  SIGNAL mux_1661_cse : STD_LOGIC;
  SIGNAL mux_1789_cse : STD_LOGIC;
  SIGNAL mux_1917_cse : STD_LOGIC;
  SIGNAL mux_2045_cse : STD_LOGIC;
  SIGNAL nor_697_cse : STD_LOGIC;
  SIGNAL nor_653_cse : STD_LOGIC;
  SIGNAL mux_3254_cse : STD_LOGIC;
  SIGNAL mux_3555_cse : STD_LOGIC;
  SIGNAL or_3008_cse : STD_LOGIC;
  SIGNAL mux_155_cse : STD_LOGIC;
  SIGNAL mux_171_cse : STD_LOGIC;
  SIGNAL mux_1036_cse : STD_LOGIC;
  SIGNAL mux_981_cse : STD_LOGIC;
  SIGNAL nand_386_cse : STD_LOGIC;
  SIGNAL mux_2465_cse : STD_LOGIC;
  SIGNAL or_2528_cse : STD_LOGIC;
  SIGNAL or_2534_cse : STD_LOGIC;
  SIGNAL nand_173_cse : STD_LOGIC;
  SIGNAL or_2541_cse : STD_LOGIC;
  SIGNAL mux_2516_cse : STD_LOGIC;
  SIGNAL mux_2494_cse : STD_LOGIC;
  SIGNAL mux_2515_cse : STD_LOGIC;
  SIGNAL mux_544_cse : STD_LOGIC;
  SIGNAL mux_2171_cse : STD_LOGIC;
  SIGNAL mux_2203_cse : STD_LOGIC;
  SIGNAL mux_3281_cse : STD_LOGIC;
  SIGNAL mux_648_cse : STD_LOGIC;
  SIGNAL mux_2998_cse : STD_LOGIC;
  SIGNAL or_2835_cse : STD_LOGIC;
  SIGNAL mux_259_cse : STD_LOGIC;
  SIGNAL mux_3245_cse : STD_LOGIC;
  SIGNAL mux_498_cse : STD_LOGIC;
  SIGNAL mux_161_cse : STD_LOGIC;
  SIGNAL mux_340_cse : STD_LOGIC;
  SIGNAL mux_375_cse : STD_LOGIC;
  SIGNAL mux_2643_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_acc_psp_sva_1 : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_psp_sva : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL COMP_LOOP_10_mul_mut : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mux_2698_itm : STD_LOGIC;
  SIGNAL mux_2757_itm : STD_LOGIC;
  SIGNAL mux_2840_itm : STD_LOGIC;
  SIGNAL mux_3485_itm : STD_LOGIC;
  SIGNAL mux_3494_itm : STD_LOGIC;
  SIGNAL and_dcpl_332 : STD_LOGIC;
  SIGNAL z_out : STD_LOGIC_VECTOR (12 DOWNTO 0);
  SIGNAL and_dcpl_333 : STD_LOGIC;
  SIGNAL and_dcpl_338 : STD_LOGIC;
  SIGNAL and_dcpl_340 : STD_LOGIC;
  SIGNAL and_dcpl_342 : STD_LOGIC;
  SIGNAL and_dcpl_344 : STD_LOGIC;
  SIGNAL and_dcpl_345 : STD_LOGIC;
  SIGNAL and_dcpl_349 : STD_LOGIC;
  SIGNAL and_dcpl_350 : STD_LOGIC;
  SIGNAL and_dcpl_356 : STD_LOGIC;
  SIGNAL and_dcpl_359 : STD_LOGIC;
  SIGNAL z_out_1 : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL and_dcpl_367 : STD_LOGIC;
  SIGNAL and_dcpl_371 : STD_LOGIC;
  SIGNAL and_dcpl_383 : STD_LOGIC;
  SIGNAL and_dcpl_390 : STD_LOGIC;
  SIGNAL and_dcpl_393 : STD_LOGIC;
  SIGNAL and_dcpl_403 : STD_LOGIC;
  SIGNAL and_dcpl_411 : STD_LOGIC;
  SIGNAL and_dcpl_412 : STD_LOGIC;
  SIGNAL and_dcpl_422 : STD_LOGIC;
  SIGNAL and_dcpl_428 : STD_LOGIC;
  SIGNAL and_dcpl_432 : STD_LOGIC;
  SIGNAL and_dcpl_446 : STD_LOGIC;
  SIGNAL and_dcpl_453 : STD_LOGIC;
  SIGNAL and_dcpl_460 : STD_LOGIC;
  SIGNAL and_dcpl_468 : STD_LOGIC;
  SIGNAL and_dcpl_472 : STD_LOGIC;
  SIGNAL and_dcpl_473 : STD_LOGIC;
  SIGNAL and_dcpl_475 : STD_LOGIC;
  SIGNAL and_dcpl_481 : STD_LOGIC;
  SIGNAL and_dcpl_486 : STD_LOGIC;
  SIGNAL and_dcpl_488 : STD_LOGIC;
  SIGNAL and_dcpl_493 : STD_LOGIC;
  SIGNAL and_dcpl_494 : STD_LOGIC;
  SIGNAL and_dcpl_495 : STD_LOGIC;
  SIGNAL and_dcpl_500 : STD_LOGIC;
  SIGNAL and_dcpl_503 : STD_LOGIC;
  SIGNAL and_dcpl_505 : STD_LOGIC;
  SIGNAL and_dcpl_507 : STD_LOGIC;
  SIGNAL and_dcpl_510 : STD_LOGIC;
  SIGNAL and_dcpl_513 : STD_LOGIC;
  SIGNAL z_out_3 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL and_dcpl_531 : STD_LOGIC;
  SIGNAL and_dcpl_539 : STD_LOGIC;
  SIGNAL and_dcpl_540 : STD_LOGIC;
  SIGNAL and_dcpl_544 : STD_LOGIC;
  SIGNAL and_dcpl_551 : STD_LOGIC;
  SIGNAL and_dcpl_553 : STD_LOGIC;
  SIGNAL and_dcpl_557 : STD_LOGIC;
  SIGNAL and_dcpl_561 : STD_LOGIC;
  SIGNAL z_out_4 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL and_dcpl_567 : STD_LOGIC;
  SIGNAL and_dcpl_568 : STD_LOGIC;
  SIGNAL and_dcpl_569 : STD_LOGIC;
  SIGNAL and_dcpl_594 : STD_LOGIC;
  SIGNAL z_out_5 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL and_dcpl_627 : STD_LOGIC;
  SIGNAL and_dcpl_628 : STD_LOGIC;
  SIGNAL and_dcpl_631 : STD_LOGIC;
  SIGNAL and_dcpl_636 : STD_LOGIC;
  SIGNAL and_dcpl_642 : STD_LOGIC;
  SIGNAL or_tmp_3282 : STD_LOGIC;
  SIGNAL not_tmp_834 : STD_LOGIC;
  SIGNAL not_tmp_835 : STD_LOGIC;
  SIGNAL not_tmp_838 : STD_LOGIC;
  SIGNAL and_dcpl_647 : STD_LOGIC;
  SIGNAL and_dcpl_650 : STD_LOGIC;
  SIGNAL z_out_6 : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL and_dcpl_660 : STD_LOGIC;
  SIGNAL and_dcpl_669 : STD_LOGIC;
  SIGNAL and_dcpl_678 : STD_LOGIC;
  SIGNAL and_dcpl_686 : STD_LOGIC;
  SIGNAL z_out_7 : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL or_tmp_3307 : STD_LOGIC;
  SIGNAL or_tmp_3312 : STD_LOGIC;
  SIGNAL or_tmp_3326 : STD_LOGIC;
  SIGNAL z_out_8 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL p_sva : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL r_sva : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL STAGE_LOOP_i_3_0_sva : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL STAGE_LOOP_lshift_psp_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL modExp_result_sva : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL modExp_exp_1_7_1_sva : STD_LOGIC;
  SIGNAL modExp_exp_1_6_1_sva : STD_LOGIC;
  SIGNAL modExp_exp_1_5_1_sva : STD_LOGIC;
  SIGNAL modExp_exp_1_4_1_sva : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_nor_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_2_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_4_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_5_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_6_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_8_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_9_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_11_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_12_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_13_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_14_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_nor_1_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_12_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_62_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_64_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_68_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_139_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_140_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_141_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_143_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_144_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_145_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_146_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_147_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_148_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_149_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_134_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_137_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_305_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_10_acc_8_itm : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL STAGE_LOOP_i_3_0_sva_mx0c1 : STD_LOGIC;
  SIGNAL STAGE_LOOP_i_3_0_sva_2 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL COMP_LOOP_1_acc_5_mut_mx0w5 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_1_modExp_1_while_if_mul_mut_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL STAGE_LOOP_lshift_psp_sva_mx0w0 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL VEC_LOOP_j_sva_11_0_mx0c1 : STD_LOGIC;
  SIGNAL modExp_result_sva_mx0c0 : STD_LOGIC;
  SIGNAL operator_64_false_slc_modExp_exp_63_1_3 : STD_LOGIC_VECTOR (62 DOWNTO 0);
  SIGNAL modulo_qr_sva_1_mx0w6 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL modExp_while_and_3 : STD_LOGIC;
  SIGNAL modExp_while_and_5 : STD_LOGIC;
  SIGNAL and_317_m1c : STD_LOGIC;
  SIGNAL modExp_result_and_rgt : STD_LOGIC;
  SIGNAL modExp_result_and_1_rgt : STD_LOGIC;
  SIGNAL and_978_ssc : STD_LOGIC;
  SIGNAL COMP_LOOP_or_32_cse : STD_LOGIC;
  SIGNAL or_80_cse : STD_LOGIC;
  SIGNAL and_816_cse : STD_LOGIC;
  SIGNAL and_815_cse : STD_LOGIC;
  SIGNAL and_825_cse : STD_LOGIC;
  SIGNAL nor_1670_cse : STD_LOGIC;
  SIGNAL and_824_ssc : STD_LOGIC;
  SIGNAL COMP_LOOP_or_54_ssc : STD_LOGIC;
  SIGNAL COMP_LOOP_or_55_ssc : STD_LOGIC;
  SIGNAL and_872_ssc : STD_LOGIC;
  SIGNAL and_820_cse : STD_LOGIC;
  SIGNAL and_830_cse : STD_LOGIC;
  SIGNAL and_842_cse : STD_LOGIC;
  SIGNAL and_849_cse : STD_LOGIC;
  SIGNAL and_870_cse : STD_LOGIC;
  SIGNAL and_873_cse : STD_LOGIC;
  SIGNAL and_827_cse : STD_LOGIC;
  SIGNAL and_835_cse : STD_LOGIC;
  SIGNAL mux_tmp_3828 : STD_LOGIC;
  SIGNAL mux_tmp_3830 : STD_LOGIC;
  SIGNAL nor_tmp_549 : STD_LOGIC;
  SIGNAL or_tmp_3337 : STD_LOGIC;
  SIGNAL or_tmp_3339 : STD_LOGIC;
  SIGNAL mux_tmp_3839 : STD_LOGIC;
  SIGNAL mux_tmp_3841 : STD_LOGIC;
  SIGNAL or_tmp_3344 : STD_LOGIC;
  SIGNAL nor_tmp_552 : STD_LOGIC;
  SIGNAL or_tmp_3347 : STD_LOGIC;
  SIGNAL mux_tmp_3848 : STD_LOGIC;
  SIGNAL nor_tmp_554 : STD_LOGIC;
  SIGNAL or_tmp_3352 : STD_LOGIC;
  SIGNAL mux_tmp_3856 : STD_LOGIC;
  SIGNAL mux_tmp_3864 : STD_LOGIC;
  SIGNAL or_tmp_3357 : STD_LOGIC;
  SIGNAL or_tmp_3381 : STD_LOGIC;
  SIGNAL or_tmp_3382 : STD_LOGIC;
  SIGNAL or_tmp_3384 : STD_LOGIC;
  SIGNAL mux_tmp_3892 : STD_LOGIC;
  SIGNAL not_tmp_882 : STD_LOGIC;
  SIGNAL not_tmp_883 : STD_LOGIC;
  SIGNAL or_tmp_3402 : STD_LOGIC;
  SIGNAL mux_tmp_3903 : STD_LOGIC;
  SIGNAL or_tmp_3403 : STD_LOGIC;
  SIGNAL mux_tmp_3906 : STD_LOGIC;
  SIGNAL mux_tmp_3907 : STD_LOGIC;
  SIGNAL or_tmp_3409 : STD_LOGIC;
  SIGNAL operator_64_false_mux1h_2_rgt : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL operator_64_false_acc_mut_64 : STD_LOGIC;
  SIGNAL operator_64_false_acc_mut_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL or_2914_cse : STD_LOGIC;
  SIGNAL or_2400_cse : STD_LOGIC;
  SIGNAL and_521_cse : STD_LOGIC;
  SIGNAL nor_1704_cse : STD_LOGIC;
  SIGNAL or_2855_cse : STD_LOGIC;
  SIGNAL or_2965_cse : STD_LOGIC;
  SIGNAL mux_3935_cse : STD_LOGIC;
  SIGNAL or_3532_cse : STD_LOGIC;
  SIGNAL or_2421_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_or_61_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_or_24_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_633_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_685_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_or_65_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_687_itm : STD_LOGIC;
  SIGNAL STAGE_LOOP_acc_itm_2_1 : STD_LOGIC;
  SIGNAL z_out_2_12_1 : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL nor_1657_cse : STD_LOGIC;

  SIGNAL or_651_nl : STD_LOGIC;
  SIGNAL or_650_nl : STD_LOGIC;
  SIGNAL or_638_nl : STD_LOGIC;
  SIGNAL or_637_nl : STD_LOGIC;
  SIGNAL or_859_nl : STD_LOGIC;
  SIGNAL or_858_nl : STD_LOGIC;
  SIGNAL or_1093_nl : STD_LOGIC;
  SIGNAL or_1092_nl : STD_LOGIC;
  SIGNAL or_1080_nl : STD_LOGIC;
  SIGNAL or_1079_nl : STD_LOGIC;
  SIGNAL or_1301_nl : STD_LOGIC;
  SIGNAL or_1300_nl : STD_LOGIC;
  SIGNAL or_1535_nl : STD_LOGIC;
  SIGNAL or_1534_nl : STD_LOGIC;
  SIGNAL or_1522_nl : STD_LOGIC;
  SIGNAL or_1521_nl : STD_LOGIC;
  SIGNAL or_1743_nl : STD_LOGIC;
  SIGNAL or_1742_nl : STD_LOGIC;
  SIGNAL nand_259_nl : STD_LOGIC;
  SIGNAL or_1976_nl : STD_LOGIC;
  SIGNAL or_1964_nl : STD_LOGIC;
  SIGNAL or_1963_nl : STD_LOGIC;
  SIGNAL nand_231_nl : STD_LOGIC;
  SIGNAL or_2184_nl : STD_LOGIC;
  SIGNAL nor_1584_nl : STD_LOGIC;
  SIGNAL and_739_nl : STD_LOGIC;
  SIGNAL modulo_result_or_nl : STD_LOGIC;
  SIGNAL mux_2231_nl : STD_LOGIC;
  SIGNAL mux_2230_nl : STD_LOGIC;
  SIGNAL mux_2229_nl : STD_LOGIC;
  SIGNAL mux_2228_nl : STD_LOGIC;
  SIGNAL mux_2227_nl : STD_LOGIC;
  SIGNAL mux_2226_nl : STD_LOGIC;
  SIGNAL mux_2225_nl : STD_LOGIC;
  SIGNAL mux_2224_nl : STD_LOGIC;
  SIGNAL nand_195_nl : STD_LOGIC;
  SIGNAL mux_2223_nl : STD_LOGIC;
  SIGNAL mux_2222_nl : STD_LOGIC;
  SIGNAL mux_2221_nl : STD_LOGIC;
  SIGNAL or_2375_nl : STD_LOGIC;
  SIGNAL mux_2220_nl : STD_LOGIC;
  SIGNAL mux_2219_nl : STD_LOGIC;
  SIGNAL mux_2218_nl : STD_LOGIC;
  SIGNAL mux_2217_nl : STD_LOGIC;
  SIGNAL mux_2216_nl : STD_LOGIC;
  SIGNAL or_2373_nl : STD_LOGIC;
  SIGNAL or_2371_nl : STD_LOGIC;
  SIGNAL mux_2215_nl : STD_LOGIC;
  SIGNAL mux_2214_nl : STD_LOGIC;
  SIGNAL mux_2213_nl : STD_LOGIC;
  SIGNAL mux_2212_nl : STD_LOGIC;
  SIGNAL mux_2211_nl : STD_LOGIC;
  SIGNAL mux_2210_nl : STD_LOGIC;
  SIGNAL mux_2209_nl : STD_LOGIC;
  SIGNAL or_2367_nl : STD_LOGIC;
  SIGNAL mux_2208_nl : STD_LOGIC;
  SIGNAL mux_2207_nl : STD_LOGIC;
  SIGNAL mux_2206_nl : STD_LOGIC;
  SIGNAL mux_2205_nl : STD_LOGIC;
  SIGNAL mux_2204_nl : STD_LOGIC;
  SIGNAL mux_2202_nl : STD_LOGIC;
  SIGNAL mux_2201_nl : STD_LOGIC;
  SIGNAL mux_2200_nl : STD_LOGIC;
  SIGNAL or_2364_nl : STD_LOGIC;
  SIGNAL mux_2199_nl : STD_LOGIC;
  SIGNAL mux_2198_nl : STD_LOGIC;
  SIGNAL mux_2197_nl : STD_LOGIC;
  SIGNAL or_2362_nl : STD_LOGIC;
  SIGNAL or_2360_nl : STD_LOGIC;
  SIGNAL mux_2196_nl : STD_LOGIC;
  SIGNAL mux_2195_nl : STD_LOGIC;
  SIGNAL mux_2194_nl : STD_LOGIC;
  SIGNAL mux_2193_nl : STD_LOGIC;
  SIGNAL mux_2192_nl : STD_LOGIC;
  SIGNAL mux_2191_nl : STD_LOGIC;
  SIGNAL mux_2190_nl : STD_LOGIC;
  SIGNAL mux_2189_nl : STD_LOGIC;
  SIGNAL mux_2188_nl : STD_LOGIC;
  SIGNAL mux_2187_nl : STD_LOGIC;
  SIGNAL mux_2186_nl : STD_LOGIC;
  SIGNAL mux_2185_nl : STD_LOGIC;
  SIGNAL mux_2184_nl : STD_LOGIC;
  SIGNAL mux_2183_nl : STD_LOGIC;
  SIGNAL mux_2182_nl : STD_LOGIC;
  SIGNAL mux_2181_nl : STD_LOGIC;
  SIGNAL mux_2180_nl : STD_LOGIC;
  SIGNAL mux_2179_nl : STD_LOGIC;
  SIGNAL or_2357_nl : STD_LOGIC;
  SIGNAL mux_2177_nl : STD_LOGIC;
  SIGNAL or_2355_nl : STD_LOGIC;
  SIGNAL mux_2174_nl : STD_LOGIC;
  SIGNAL mux_2173_nl : STD_LOGIC;
  SIGNAL mux_2170_nl : STD_LOGIC;
  SIGNAL mux_2169_nl : STD_LOGIC;
  SIGNAL or_2351_nl : STD_LOGIC;
  SIGNAL mux_2168_nl : STD_LOGIC;
  SIGNAL mux_2167_nl : STD_LOGIC;
  SIGNAL or_2347_nl : STD_LOGIC;
  SIGNAL mux_2166_nl : STD_LOGIC;
  SIGNAL mux_2165_nl : STD_LOGIC;
  SIGNAL mux_2164_nl : STD_LOGIC;
  SIGNAL mux_2163_nl : STD_LOGIC;
  SIGNAL mux_2162_nl : STD_LOGIC;
  SIGNAL mux_2161_nl : STD_LOGIC;
  SIGNAL mux_2160_nl : STD_LOGIC;
  SIGNAL or_2343_nl : STD_LOGIC;
  SIGNAL mux_2158_nl : STD_LOGIC;
  SIGNAL mux_2157_nl : STD_LOGIC;
  SIGNAL mux_2156_nl : STD_LOGIC;
  SIGNAL mux_2155_nl : STD_LOGIC;
  SIGNAL mux_2154_nl : STD_LOGIC;
  SIGNAL mux_2153_nl : STD_LOGIC;
  SIGNAL mux_2152_nl : STD_LOGIC;
  SIGNAL mux_2151_nl : STD_LOGIC;
  SIGNAL mux_2150_nl : STD_LOGIC;
  SIGNAL mux_2149_nl : STD_LOGIC;
  SIGNAL mux_2148_nl : STD_LOGIC;
  SIGNAL mux_2147_nl : STD_LOGIC;
  SIGNAL mux_2146_nl : STD_LOGIC;
  SIGNAL or_2339_nl : STD_LOGIC;
  SIGNAL mux_2144_nl : STD_LOGIC;
  SIGNAL mux_2143_nl : STD_LOGIC;
  SIGNAL mux_2142_nl : STD_LOGIC;
  SIGNAL mux_2141_nl : STD_LOGIC;
  SIGNAL mux_2140_nl : STD_LOGIC;
  SIGNAL mux_2139_nl : STD_LOGIC;
  SIGNAL or_2335_nl : STD_LOGIC;
  SIGNAL mux_2138_nl : STD_LOGIC;
  SIGNAL mux_2137_nl : STD_LOGIC;
  SIGNAL mux_2136_nl : STD_LOGIC;
  SIGNAL nand_197_nl : STD_LOGIC;
  SIGNAL mux_2135_nl : STD_LOGIC;
  SIGNAL mux_2134_nl : STD_LOGIC;
  SIGNAL mux_2133_nl : STD_LOGIC;
  SIGNAL mux_2331_nl : STD_LOGIC;
  SIGNAL mux_2330_nl : STD_LOGIC;
  SIGNAL mux_2329_nl : STD_LOGIC;
  SIGNAL mux_2328_nl : STD_LOGIC;
  SIGNAL mux_2327_nl : STD_LOGIC;
  SIGNAL mux_2326_nl : STD_LOGIC;
  SIGNAL mux_2325_nl : STD_LOGIC;
  SIGNAL mux_2324_nl : STD_LOGIC;
  SIGNAL mux_2323_nl : STD_LOGIC;
  SIGNAL mux_2322_nl : STD_LOGIC;
  SIGNAL and_519_nl : STD_LOGIC;
  SIGNAL mux_2321_nl : STD_LOGIC;
  SIGNAL mux_2320_nl : STD_LOGIC;
  SIGNAL mux_2319_nl : STD_LOGIC;
  SIGNAL mux_2318_nl : STD_LOGIC;
  SIGNAL mux_2317_nl : STD_LOGIC;
  SIGNAL mux_2316_nl : STD_LOGIC;
  SIGNAL mux_2315_nl : STD_LOGIC;
  SIGNAL mux_2314_nl : STD_LOGIC;
  SIGNAL mux_2313_nl : STD_LOGIC;
  SIGNAL mux_2312_nl : STD_LOGIC;
  SIGNAL mux_2310_nl : STD_LOGIC;
  SIGNAL mux_2309_nl : STD_LOGIC;
  SIGNAL or_2418_nl : STD_LOGIC;
  SIGNAL mux_2308_nl : STD_LOGIC;
  SIGNAL mux_2307_nl : STD_LOGIC;
  SIGNAL mux_2306_nl : STD_LOGIC;
  SIGNAL mux_2305_nl : STD_LOGIC;
  SIGNAL mux_2304_nl : STD_LOGIC;
  SIGNAL mux_2303_nl : STD_LOGIC;
  SIGNAL mux_2302_nl : STD_LOGIC;
  SIGNAL mux_2301_nl : STD_LOGIC;
  SIGNAL mux_2300_nl : STD_LOGIC;
  SIGNAL mux_2299_nl : STD_LOGIC;
  SIGNAL mux_2298_nl : STD_LOGIC;
  SIGNAL mux_2297_nl : STD_LOGIC;
  SIGNAL mux_2296_nl : STD_LOGIC;
  SIGNAL mux_2295_nl : STD_LOGIC;
  SIGNAL mux_2294_nl : STD_LOGIC;
  SIGNAL or_2408_nl : STD_LOGIC;
  SIGNAL mux_2292_nl : STD_LOGIC;
  SIGNAL mux_2291_nl : STD_LOGIC;
  SIGNAL mux_2290_nl : STD_LOGIC;
  SIGNAL mux_2288_nl : STD_LOGIC;
  SIGNAL mux_2286_nl : STD_LOGIC;
  SIGNAL mux_2285_nl : STD_LOGIC;
  SIGNAL or_2406_nl : STD_LOGIC;
  SIGNAL or_2404_nl : STD_LOGIC;
  SIGNAL mux_2284_nl : STD_LOGIC;
  SIGNAL mux_2283_nl : STD_LOGIC;
  SIGNAL mux_2282_nl : STD_LOGIC;
  SIGNAL mux_2281_nl : STD_LOGIC;
  SIGNAL mux_2280_nl : STD_LOGIC;
  SIGNAL or_2403_nl : STD_LOGIC;
  SIGNAL mux_2279_nl : STD_LOGIC;
  SIGNAL mux_2278_nl : STD_LOGIC;
  SIGNAL or_2402_nl : STD_LOGIC;
  SIGNAL mux_2277_nl : STD_LOGIC;
  SIGNAL mux_2276_nl : STD_LOGIC;
  SIGNAL mux_2275_nl : STD_LOGIC;
  SIGNAL mux_2274_nl : STD_LOGIC;
  SIGNAL mux_2273_nl : STD_LOGIC;
  SIGNAL mux_2272_nl : STD_LOGIC;
  SIGNAL nor_295_nl : STD_LOGIC;
  SIGNAL mux_2271_nl : STD_LOGIC;
  SIGNAL mux_2270_nl : STD_LOGIC;
  SIGNAL mux_2269_nl : STD_LOGIC;
  SIGNAL mux_2268_nl : STD_LOGIC;
  SIGNAL mux_2267_nl : STD_LOGIC;
  SIGNAL or_2398_nl : STD_LOGIC;
  SIGNAL mux_2266_nl : STD_LOGIC;
  SIGNAL mux_2265_nl : STD_LOGIC;
  SIGNAL mux_2264_nl : STD_LOGIC;
  SIGNAL mux_2263_nl : STD_LOGIC;
  SIGNAL mux_2261_nl : STD_LOGIC;
  SIGNAL mux_2260_nl : STD_LOGIC;
  SIGNAL mux_2259_nl : STD_LOGIC;
  SIGNAL or_2395_nl : STD_LOGIC;
  SIGNAL mux_2257_nl : STD_LOGIC;
  SIGNAL mux_2256_nl : STD_LOGIC;
  SIGNAL mux_2255_nl : STD_LOGIC;
  SIGNAL mux_2254_nl : STD_LOGIC;
  SIGNAL mux_2253_nl : STD_LOGIC;
  SIGNAL mux_2251_nl : STD_LOGIC;
  SIGNAL mux_2250_nl : STD_LOGIC;
  SIGNAL mux_2249_nl : STD_LOGIC;
  SIGNAL or_2392_nl : STD_LOGIC;
  SIGNAL mux_2248_nl : STD_LOGIC;
  SIGNAL mux_2247_nl : STD_LOGIC;
  SIGNAL mux_2246_nl : STD_LOGIC;
  SIGNAL mux_2245_nl : STD_LOGIC;
  SIGNAL or_2390_nl : STD_LOGIC;
  SIGNAL mux_2244_nl : STD_LOGIC;
  SIGNAL or_2385_nl : STD_LOGIC;
  SIGNAL mux_2243_nl : STD_LOGIC;
  SIGNAL mux_2237_nl : STD_LOGIC;
  SIGNAL nand_51_nl : STD_LOGIC;
  SIGNAL mux_2236_nl : STD_LOGIC;
  SIGNAL mux_2346_nl : STD_LOGIC;
  SIGNAL mux_2345_nl : STD_LOGIC;
  SIGNAL mux_2344_nl : STD_LOGIC;
  SIGNAL nand_189_nl : STD_LOGIC;
  SIGNAL mux_2343_nl : STD_LOGIC;
  SIGNAL and_517_nl : STD_LOGIC;
  SIGNAL nor_752_nl : STD_LOGIC;
  SIGNAL mux_2341_nl : STD_LOGIC;
  SIGNAL or_3386_nl : STD_LOGIC;
  SIGNAL nand_190_nl : STD_LOGIC;
  SIGNAL or_2438_nl : STD_LOGIC;
  SIGNAL mux_2340_nl : STD_LOGIC;
  SIGNAL or_2437_nl : STD_LOGIC;
  SIGNAL mux_2339_nl : STD_LOGIC;
  SIGNAL mux_2338_nl : STD_LOGIC;
  SIGNAL mux_2337_nl : STD_LOGIC;
  SIGNAL mux_2336_nl : STD_LOGIC;
  SIGNAL mux_2335_nl : STD_LOGIC;
  SIGNAL or_2435_nl : STD_LOGIC;
  SIGNAL or_2433_nl : STD_LOGIC;
  SIGNAL or_2431_nl : STD_LOGIC;
  SIGNAL or_2430_nl : STD_LOGIC;
  SIGNAL mux_2334_nl : STD_LOGIC;
  SIGNAL nand_191_nl : STD_LOGIC;
  SIGNAL mux_2333_nl : STD_LOGIC;
  SIGNAL or_2427_nl : STD_LOGIC;
  SIGNAL or_2426_nl : STD_LOGIC;
  SIGNAL mux_2418_nl : STD_LOGIC;
  SIGNAL mux_2417_nl : STD_LOGIC;
  SIGNAL mux_2416_nl : STD_LOGIC;
  SIGNAL mux_2415_nl : STD_LOGIC;
  SIGNAL mux_2414_nl : STD_LOGIC;
  SIGNAL mux_2413_nl : STD_LOGIC;
  SIGNAL mux_2412_nl : STD_LOGIC;
  SIGNAL mux_2411_nl : STD_LOGIC;
  SIGNAL mux_2410_nl : STD_LOGIC;
  SIGNAL mux_2409_nl : STD_LOGIC;
  SIGNAL mux_2408_nl : STD_LOGIC;
  SIGNAL mux_2407_nl : STD_LOGIC;
  SIGNAL mux_2406_nl : STD_LOGIC;
  SIGNAL mux_2405_nl : STD_LOGIC;
  SIGNAL mux_2404_nl : STD_LOGIC;
  SIGNAL mux_2403_nl : STD_LOGIC;
  SIGNAL mux_2402_nl : STD_LOGIC;
  SIGNAL mux_2401_nl : STD_LOGIC;
  SIGNAL mux_2400_nl : STD_LOGIC;
  SIGNAL mux_2399_nl : STD_LOGIC;
  SIGNAL mux_2398_nl : STD_LOGIC;
  SIGNAL mux_2397_nl : STD_LOGIC;
  SIGNAL mux_2396_nl : STD_LOGIC;
  SIGNAL mux_2395_nl : STD_LOGIC;
  SIGNAL mux_2394_nl : STD_LOGIC;
  SIGNAL mux_2393_nl : STD_LOGIC;
  SIGNAL mux_2392_nl : STD_LOGIC;
  SIGNAL mux_2391_nl : STD_LOGIC;
  SIGNAL mux_2390_nl : STD_LOGIC;
  SIGNAL mux_2384_nl : STD_LOGIC;
  SIGNAL mux_2383_nl : STD_LOGIC;
  SIGNAL mux_2381_nl : STD_LOGIC;
  SIGNAL mux_2380_nl : STD_LOGIC;
  SIGNAL mux_2379_nl : STD_LOGIC;
  SIGNAL mux_2374_nl : STD_LOGIC;
  SIGNAL mux_2373_nl : STD_LOGIC;
  SIGNAL mux_2372_nl : STD_LOGIC;
  SIGNAL mux_2368_nl : STD_LOGIC;
  SIGNAL mux_2367_nl : STD_LOGIC;
  SIGNAL mux_2366_nl : STD_LOGIC;
  SIGNAL mux_2362_nl : STD_LOGIC;
  SIGNAL mux_2360_nl : STD_LOGIC;
  SIGNAL mux_2358_nl : STD_LOGIC;
  SIGNAL mux_2357_nl : STD_LOGIC;
  SIGNAL mux_2354_nl : STD_LOGIC;
  SIGNAL mux_2351_nl : STD_LOGIC;
  SIGNAL mux_2349_nl : STD_LOGIC;
  SIGNAL mux_2452_nl : STD_LOGIC;
  SIGNAL mux_2451_nl : STD_LOGIC;
  SIGNAL mux_2450_nl : STD_LOGIC;
  SIGNAL mux_2449_nl : STD_LOGIC;
  SIGNAL or_3396_nl : STD_LOGIC;
  SIGNAL nand_175_nl : STD_LOGIC;
  SIGNAL modExp_while_if_mux1h_nl : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL and_323_nl : STD_LOGIC;
  SIGNAL mux_3257_nl : STD_LOGIC;
  SIGNAL mux_3256_nl : STD_LOGIC;
  SIGNAL nor_640_nl : STD_LOGIC;
  SIGNAL mux_3255_nl : STD_LOGIC;
  SIGNAL or_2920_nl : STD_LOGIC;
  SIGNAL mux_3253_nl : STD_LOGIC;
  SIGNAL and_421_nl : STD_LOGIC;
  SIGNAL mux_3252_nl : STD_LOGIC;
  SIGNAL nor_641_nl : STD_LOGIC;
  SIGNAL mux_3251_nl : STD_LOGIC;
  SIGNAL nand_85_nl : STD_LOGIC;
  SIGNAL mux_3250_nl : STD_LOGIC;
  SIGNAL nor_642_nl : STD_LOGIC;
  SIGNAL nor_643_nl : STD_LOGIC;
  SIGNAL mux_3249_nl : STD_LOGIC;
  SIGNAL mux_3248_nl : STD_LOGIC;
  SIGNAL and_422_nl : STD_LOGIC;
  SIGNAL mux_3247_nl : STD_LOGIC;
  SIGNAL and_423_nl : STD_LOGIC;
  SIGNAL mux_3246_nl : STD_LOGIC;
  SIGNAL or_2910_nl : STD_LOGIC;
  SIGNAL nor_644_nl : STD_LOGIC;
  SIGNAL nor_645_nl : STD_LOGIC;
  SIGNAL modExp_while_if_and_nl : STD_LOGIC;
  SIGNAL modExp_while_if_and_1_nl : STD_LOGIC;
  SIGNAL and_261_nl : STD_LOGIC;
  SIGNAL mux_2545_nl : STD_LOGIC;
  SIGNAL mux_2544_nl : STD_LOGIC;
  SIGNAL mux_2543_nl : STD_LOGIC;
  SIGNAL mux_2542_nl : STD_LOGIC;
  SIGNAL mux_2541_nl : STD_LOGIC;
  SIGNAL mux_2540_nl : STD_LOGIC;
  SIGNAL or_2578_nl : STD_LOGIC;
  SIGNAL mux_2630_nl : STD_LOGIC;
  SIGNAL mux_2629_nl : STD_LOGIC;
  SIGNAL mux_2628_nl : STD_LOGIC;
  SIGNAL mux_2610_nl : STD_LOGIC;
  SIGNAL mux_2609_nl : STD_LOGIC;
  SIGNAL or_2624_nl : STD_LOGIC;
  SIGNAL mux_2608_nl : STD_LOGIC;
  SIGNAL mux_2607_nl : STD_LOGIC;
  SIGNAL or_2622_nl : STD_LOGIC;
  SIGNAL mux_2532_nl : STD_LOGIC;
  SIGNAL mux_2617_nl : STD_LOGIC;
  SIGNAL mux_2616_nl : STD_LOGIC;
  SIGNAL mux_2615_nl : STD_LOGIC;
  SIGNAL mux_2614_nl : STD_LOGIC;
  SIGNAL nor_696_nl : STD_LOGIC;
  SIGNAL or_2627_nl : STD_LOGIC;
  SIGNAL mux_2600_nl : STD_LOGIC;
  SIGNAL mux_2599_nl : STD_LOGIC;
  SIGNAL mux_2598_nl : STD_LOGIC;
  SIGNAL mux_2524_nl : STD_LOGIC;
  SIGNAL mux_2523_nl : STD_LOGIC;
  SIGNAL mux_2522_nl : STD_LOGIC;
  SIGNAL mux_2521_nl : STD_LOGIC;
  SIGNAL mux_2520_nl : STD_LOGIC;
  SIGNAL mux_2624_nl : STD_LOGIC;
  SIGNAL mux_2623_nl : STD_LOGIC;
  SIGNAL mux_2622_nl : STD_LOGIC;
  SIGNAL mux_2620_nl : STD_LOGIC;
  SIGNAL mux_2619_nl : STD_LOGIC;
  SIGNAL mux_2604_nl : STD_LOGIC;
  SIGNAL mux_2603_nl : STD_LOGIC;
  SIGNAL mux_2602_nl : STD_LOGIC;
  SIGNAL mux_2586_nl : STD_LOGIC;
  SIGNAL or_2620_nl : STD_LOGIC;
  SIGNAL mux_2508_nl : STD_LOGIC;
  SIGNAL mux_2613_nl : STD_LOGIC;
  SIGNAL or_2625_nl : STD_LOGIC;
  SIGNAL mux_2597_nl : STD_LOGIC;
  SIGNAL mux_2596_nl : STD_LOGIC;
  SIGNAL mux_2595_nl : STD_LOGIC;
  SIGNAL mux_2594_nl : STD_LOGIC;
  SIGNAL or_2616_nl : STD_LOGIC;
  SIGNAL mux_2593_nl : STD_LOGIC;
  SIGNAL nor_704_nl : STD_LOGIC;
  SIGNAL or_2612_nl : STD_LOGIC;
  SIGNAL mux_2501_nl : STD_LOGIC;
  SIGNAL mux_2500_nl : STD_LOGIC;
  SIGNAL mux_2499_nl : STD_LOGIC;
  SIGNAL mux_2498_nl : STD_LOGIC;
  SIGNAL mux_2497_nl : STD_LOGIC;
  SIGNAL mux_2496_nl : STD_LOGIC;
  SIGNAL mux_2495_nl : STD_LOGIC;
  SIGNAL mux_2561_nl : STD_LOGIC;
  SIGNAL mux_2560_nl : STD_LOGIC;
  SIGNAL nor_707_nl : STD_LOGIC;
  SIGNAL or_2591_nl : STD_LOGIC;
  SIGNAL mux_2559_nl : STD_LOGIC;
  SIGNAL or_2589_nl : STD_LOGIC;
  SIGNAL mux_2490_nl : STD_LOGIC;
  SIGNAL mux_2576_nl : STD_LOGIC;
  SIGNAL mux_2575_nl : STD_LOGIC;
  SIGNAL mux_2574_nl : STD_LOGIC;
  SIGNAL mux_2572_nl : STD_LOGIC;
  SIGNAL mux_2571_nl : STD_LOGIC;
  SIGNAL mux_2570_nl : STD_LOGIC;
  SIGNAL or_2602_nl : STD_LOGIC;
  SIGNAL mux_2553_nl : STD_LOGIC;
  SIGNAL mux_2552_nl : STD_LOGIC;
  SIGNAL nor_709_nl : STD_LOGIC;
  SIGNAL mux_2551_nl : STD_LOGIC;
  SIGNAL mux_2550_nl : STD_LOGIC;
  SIGNAL mux_2478_nl : STD_LOGIC;
  SIGNAL mux_2477_nl : STD_LOGIC;
  SIGNAL mux_2585_nl : STD_LOGIC;
  SIGNAL mux_2584_nl : STD_LOGIC;
  SIGNAL mux_2583_nl : STD_LOGIC;
  SIGNAL mux_2582_nl : STD_LOGIC;
  SIGNAL mux_2581_nl : STD_LOGIC;
  SIGNAL mux_2580_nl : STD_LOGIC;
  SIGNAL mux_2579_nl : STD_LOGIC;
  SIGNAL mux_2578_nl : STD_LOGIC;
  SIGNAL or_2608_nl : STD_LOGIC;
  SIGNAL or_2606_nl : STD_LOGIC;
  SIGNAL mux_2558_nl : STD_LOGIC;
  SIGNAL mux_2557_nl : STD_LOGIC;
  SIGNAL mux_2556_nl : STD_LOGIC;
  SIGNAL mux_2464_nl : STD_LOGIC;
  SIGNAL mux_2569_nl : STD_LOGIC;
  SIGNAL mux_2568_nl : STD_LOGIC;
  SIGNAL mux_2567_nl : STD_LOGIC;
  SIGNAL mux_2566_nl : STD_LOGIC;
  SIGNAL or_2598_nl : STD_LOGIC;
  SIGNAL mux_2565_nl : STD_LOGIC;
  SIGNAL mux_2564_nl : STD_LOGIC;
  SIGNAL mux_2549_nl : STD_LOGIC;
  SIGNAL mux_2548_nl : STD_LOGIC;
  SIGNAL or_2582_nl : STD_LOGIC;
  SIGNAL mux_2547_nl : STD_LOGIC;
  SIGNAL mux_2546_nl : STD_LOGIC;
  SIGNAL or_2580_nl : STD_LOGIC;
  SIGNAL mux_3889_nl : STD_LOGIC;
  SIGNAL mux_3888_nl : STD_LOGIC;
  SIGNAL mux_3887_nl : STD_LOGIC;
  SIGNAL mux_3886_nl : STD_LOGIC;
  SIGNAL nor_1705_nl : STD_LOGIC;
  SIGNAL mux_3885_nl : STD_LOGIC;
  SIGNAL or_3549_nl : STD_LOGIC;
  SIGNAL mux_3884_nl : STD_LOGIC;
  SIGNAL mux_3883_nl : STD_LOGIC;
  SIGNAL nor_1706_nl : STD_LOGIC;
  SIGNAL and_1165_nl : STD_LOGIC;
  SIGNAL and_1166_nl : STD_LOGIC;
  SIGNAL mux_3882_nl : STD_LOGIC;
  SIGNAL mux_3881_nl : STD_LOGIC;
  SIGNAL or_3619_nl : STD_LOGIC;
  SIGNAL or_3620_nl : STD_LOGIC;
  SIGNAL mux_3880_nl : STD_LOGIC;
  SIGNAL or_3543_nl : STD_LOGIC;
  SIGNAL mux_3879_nl : STD_LOGIC;
  SIGNAL mux_3878_nl : STD_LOGIC;
  SIGNAL mux_3877_nl : STD_LOGIC;
  SIGNAL or_3541_nl : STD_LOGIC;
  SIGNAL mux_3876_nl : STD_LOGIC;
  SIGNAL nor_1708_nl : STD_LOGIC;
  SIGNAL mux_3875_nl : STD_LOGIC;
  SIGNAL mux_3874_nl : STD_LOGIC;
  SIGNAL mux_3873_nl : STD_LOGIC;
  SIGNAL mux_3872_nl : STD_LOGIC;
  SIGNAL mux_3871_nl : STD_LOGIC;
  SIGNAL or_3537_nl : STD_LOGIC;
  SIGNAL mux_3870_nl : STD_LOGIC;
  SIGNAL mux_3869_nl : STD_LOGIC;
  SIGNAL mux_3868_nl : STD_LOGIC;
  SIGNAL or_3534_nl : STD_LOGIC;
  SIGNAL mux_3867_nl : STD_LOGIC;
  SIGNAL nand_417_nl : STD_LOGIC;
  SIGNAL mux_3865_nl : STD_LOGIC;
  SIGNAL mux_3864_nl : STD_LOGIC;
  SIGNAL and_1168_nl : STD_LOGIC;
  SIGNAL mux_3863_nl : STD_LOGIC;
  SIGNAL mux_3862_nl : STD_LOGIC;
  SIGNAL mux_3861_nl : STD_LOGIC;
  SIGNAL mux_3860_nl : STD_LOGIC;
  SIGNAL mux_3859_nl : STD_LOGIC;
  SIGNAL mux_3857_nl : STD_LOGIC;
  SIGNAL or_3529_nl : STD_LOGIC;
  SIGNAL mux_3856_nl : STD_LOGIC;
  SIGNAL mux_3855_nl : STD_LOGIC;
  SIGNAL mux_3854_nl : STD_LOGIC;
  SIGNAL mux_3853_nl : STD_LOGIC;
  SIGNAL mux_3852_nl : STD_LOGIC;
  SIGNAL mux_3851_nl : STD_LOGIC;
  SIGNAL mux_3848_nl : STD_LOGIC;
  SIGNAL mux_3847_nl : STD_LOGIC;
  SIGNAL mux_3846_nl : STD_LOGIC;
  SIGNAL mux_3845_nl : STD_LOGIC;
  SIGNAL mux_3844_nl : STD_LOGIC;
  SIGNAL or_3522_nl : STD_LOGIC;
  SIGNAL mux_3840_nl : STD_LOGIC;
  SIGNAL mux_3839_nl : STD_LOGIC;
  SIGNAL mux_3838_nl : STD_LOGIC;
  SIGNAL nand_416_nl : STD_LOGIC;
  SIGNAL mux_3837_nl : STD_LOGIC;
  SIGNAL mux_3836_nl : STD_LOGIC;
  SIGNAL mux_3835_nl : STD_LOGIC;
  SIGNAL mux_3834_nl : STD_LOGIC;
  SIGNAL mux_3833_nl : STD_LOGIC;
  SIGNAL or_3513_nl : STD_LOGIC;
  SIGNAL mux_3831_nl : STD_LOGIC;
  SIGNAL or_3609_nl : STD_LOGIC;
  SIGNAL mux_3943_nl : STD_LOGIC;
  SIGNAL mux_3942_nl : STD_LOGIC;
  SIGNAL mux_3941_nl : STD_LOGIC;
  SIGNAL mux_3940_nl : STD_LOGIC;
  SIGNAL mux_3939_nl : STD_LOGIC;
  SIGNAL mux_3938_nl : STD_LOGIC;
  SIGNAL or_3612_nl : STD_LOGIC;
  SIGNAL or_3611_nl : STD_LOGIC;
  SIGNAL mux_3937_nl : STD_LOGIC;
  SIGNAL mux_3936_nl : STD_LOGIC;
  SIGNAL or_3608_nl : STD_LOGIC;
  SIGNAL mux_3934_nl : STD_LOGIC;
  SIGNAL mux_3933_nl : STD_LOGIC;
  SIGNAL or_3606_nl : STD_LOGIC;
  SIGNAL mux_3932_nl : STD_LOGIC;
  SIGNAL or_3604_nl : STD_LOGIC;
  SIGNAL nand_423_nl : STD_LOGIC;
  SIGNAL mux_3931_nl : STD_LOGIC;
  SIGNAL mux_3930_nl : STD_LOGIC;
  SIGNAL mux_3929_nl : STD_LOGIC;
  SIGNAL or_3601_nl : STD_LOGIC;
  SIGNAL mux_3928_nl : STD_LOGIC;
  SIGNAL or_3600_nl : STD_LOGIC;
  SIGNAL mux_3927_nl : STD_LOGIC;
  SIGNAL mux_3926_nl : STD_LOGIC;
  SIGNAL mux_3925_nl : STD_LOGIC;
  SIGNAL mux_3924_nl : STD_LOGIC;
  SIGNAL mux_3923_nl : STD_LOGIC;
  SIGNAL or_3599_nl : STD_LOGIC;
  SIGNAL or_3598_nl : STD_LOGIC;
  SIGNAL mux_3922_nl : STD_LOGIC;
  SIGNAL nand_420_nl : STD_LOGIC;
  SIGNAL or_3597_nl : STD_LOGIC;
  SIGNAL mux_3921_nl : STD_LOGIC;
  SIGNAL mux_3920_nl : STD_LOGIC;
  SIGNAL or_3595_nl : STD_LOGIC;
  SIGNAL mux_3919_nl : STD_LOGIC;
  SIGNAL mux_3918_nl : STD_LOGIC;
  SIGNAL or_3594_nl : STD_LOGIC;
  SIGNAL or_3593_nl : STD_LOGIC;
  SIGNAL or_3591_nl : STD_LOGIC;
  SIGNAL or_3590_nl : STD_LOGIC;
  SIGNAL mux_3917_nl : STD_LOGIC;
  SIGNAL or_3589_nl : STD_LOGIC;
  SIGNAL mux_3916_nl : STD_LOGIC;
  SIGNAL mux_3915_nl : STD_LOGIC;
  SIGNAL mux_3914_nl : STD_LOGIC;
  SIGNAL mux_3913_nl : STD_LOGIC;
  SIGNAL mux_3912_nl : STD_LOGIC;
  SIGNAL mux_3911_nl : STD_LOGIC;
  SIGNAL mux_3910_nl : STD_LOGIC;
  SIGNAL mux_3906_nl : STD_LOGIC;
  SIGNAL or_3578_nl : STD_LOGIC;
  SIGNAL or_3576_nl : STD_LOGIC;
  SIGNAL mux_3903_nl : STD_LOGIC;
  SIGNAL or_3575_nl : STD_LOGIC;
  SIGNAL mux_3902_nl : STD_LOGIC;
  SIGNAL mux_3901_nl : STD_LOGIC;
  SIGNAL or_3573_nl : STD_LOGIC;
  SIGNAL or_3572_nl : STD_LOGIC;
  SIGNAL mux_3900_nl : STD_LOGIC;
  SIGNAL mux_3899_nl : STD_LOGIC;
  SIGNAL or_3571_nl : STD_LOGIC;
  SIGNAL mux_3898_nl : STD_LOGIC;
  SIGNAL or_3569_nl : STD_LOGIC;
  SIGNAL mux_3897_nl : STD_LOGIC;
  SIGNAL or_3568_nl : STD_LOGIC;
  SIGNAL mux_3896_nl : STD_LOGIC;
  SIGNAL or_3565_nl : STD_LOGIC;
  SIGNAL mux_3895_nl : STD_LOGIC;
  SIGNAL mux_3892_nl : STD_LOGIC;
  SIGNAL or_3556_nl : STD_LOGIC;
  SIGNAL mux_3891_nl : STD_LOGIC;
  SIGNAL or_3554_nl : STD_LOGIC;
  SIGNAL mux_3890_nl : STD_LOGIC;
  SIGNAL or_3553_nl : STD_LOGIC;
  SIGNAL or_3551_nl : STD_LOGIC;
  SIGNAL or_3508_nl : STD_LOGIC;
  SIGNAL mux_2639_nl : STD_LOGIC;
  SIGNAL or_2642_nl : STD_LOGIC;
  SIGNAL mux_2638_nl : STD_LOGIC;
  SIGNAL or_2641_nl : STD_LOGIC;
  SIGNAL or_2640_nl : STD_LOGIC;
  SIGNAL or_2638_nl : STD_LOGIC;
  SIGNAL mux_3946_nl : STD_LOGIC;
  SIGNAL nor_1700_nl : STD_LOGIC;
  SIGNAL nor_1701_nl : STD_LOGIC;
  SIGNAL mux_3945_nl : STD_LOGIC;
  SIGNAL mux_3944_nl : STD_LOGIC;
  SIGNAL or_3616_nl : STD_LOGIC;
  SIGNAL or_3615_nl : STD_LOGIC;
  SIGNAL or_3613_nl : STD_LOGIC;
  SIGNAL mux_2668_nl : STD_LOGIC;
  SIGNAL mux_2667_nl : STD_LOGIC;
  SIGNAL mux_2666_nl : STD_LOGIC;
  SIGNAL mux_2665_nl : STD_LOGIC;
  SIGNAL mux_2664_nl : STD_LOGIC;
  SIGNAL mux_2663_nl : STD_LOGIC;
  SIGNAL nor_690_nl : STD_LOGIC;
  SIGNAL mux_2662_nl : STD_LOGIC;
  SIGNAL mux_2661_nl : STD_LOGIC;
  SIGNAL mux_2660_nl : STD_LOGIC;
  SIGNAL nand_170_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_8_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_9_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_10_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_11_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_12_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_13_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_14_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_15_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_16_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_17_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_18_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_19_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_20_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_21_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_22_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_23_nl : STD_LOGIC;
  SIGNAL mux_2741_nl : STD_LOGIC;
  SIGNAL mux_2740_nl : STD_LOGIC;
  SIGNAL mux_2739_nl : STD_LOGIC;
  SIGNAL mux_2738_nl : STD_LOGIC;
  SIGNAL mux_2737_nl : STD_LOGIC;
  SIGNAL and_276_nl : STD_LOGIC;
  SIGNAL mux_2735_nl : STD_LOGIC;
  SIGNAL mux_2734_nl : STD_LOGIC;
  SIGNAL nor_687_nl : STD_LOGIC;
  SIGNAL mux_2733_nl : STD_LOGIC;
  SIGNAL mux_2732_nl : STD_LOGIC;
  SIGNAL mux_2731_nl : STD_LOGIC;
  SIGNAL mux_2730_nl : STD_LOGIC;
  SIGNAL mux_2729_nl : STD_LOGIC;
  SIGNAL mux_2728_nl : STD_LOGIC;
  SIGNAL or_2666_nl : STD_LOGIC;
  SIGNAL mux_2727_nl : STD_LOGIC;
  SIGNAL and_454_nl : STD_LOGIC;
  SIGNAL mux_2726_nl : STD_LOGIC;
  SIGNAL mux_2725_nl : STD_LOGIC;
  SIGNAL mux_2724_nl : STD_LOGIC;
  SIGNAL mux_2723_nl : STD_LOGIC;
  SIGNAL mux_2722_nl : STD_LOGIC;
  SIGNAL mux_2721_nl : STD_LOGIC;
  SIGNAL mux_2720_nl : STD_LOGIC;
  SIGNAL mux_2719_nl : STD_LOGIC;
  SIGNAL mux_2718_nl : STD_LOGIC;
  SIGNAL mux_2717_nl : STD_LOGIC;
  SIGNAL mux_2716_nl : STD_LOGIC;
  SIGNAL mux_2714_nl : STD_LOGIC;
  SIGNAL mux_2713_nl : STD_LOGIC;
  SIGNAL mux_2712_nl : STD_LOGIC;
  SIGNAL mux_2711_nl : STD_LOGIC;
  SIGNAL mux_2710_nl : STD_LOGIC;
  SIGNAL mux_2707_nl : STD_LOGIC;
  SIGNAL mux_2705_nl : STD_LOGIC;
  SIGNAL mux_2704_nl : STD_LOGIC;
  SIGNAL mux_2701_nl : STD_LOGIC;
  SIGNAL mux_2699_nl : STD_LOGIC;
  SIGNAL mux_2697_nl : STD_LOGIC;
  SIGNAL mux_2696_nl : STD_LOGIC;
  SIGNAL mux_2695_nl : STD_LOGIC;
  SIGNAL mux_2694_nl : STD_LOGIC;
  SIGNAL mux_2692_nl : STD_LOGIC;
  SIGNAL mux_2689_nl : STD_LOGIC;
  SIGNAL mux_2688_nl : STD_LOGIC;
  SIGNAL mux_2687_nl : STD_LOGIC;
  SIGNAL mux_2686_nl : STD_LOGIC;
  SIGNAL mux_2685_nl : STD_LOGIC;
  SIGNAL mux_2684_nl : STD_LOGIC;
  SIGNAL mux_2683_nl : STD_LOGIC;
  SIGNAL mux_2680_nl : STD_LOGIC;
  SIGNAL mux_2679_nl : STD_LOGIC;
  SIGNAL mux_2678_nl : STD_LOGIC;
  SIGNAL or_2658_nl : STD_LOGIC;
  SIGNAL mux_2674_nl : STD_LOGIC;
  SIGNAL mux_2673_nl : STD_LOGIC;
  SIGNAL mux_2671_nl : STD_LOGIC;
  SIGNAL mux_2770_nl : STD_LOGIC;
  SIGNAL nor_678_nl : STD_LOGIC;
  SIGNAL mux_2769_nl : STD_LOGIC;
  SIGNAL nand_166_nl : STD_LOGIC;
  SIGNAL nor_679_nl : STD_LOGIC;
  SIGNAL mux_2768_nl : STD_LOGIC;
  SIGNAL or_2717_nl : STD_LOGIC;
  SIGNAL mux_2767_nl : STD_LOGIC;
  SIGNAL or_2716_nl : STD_LOGIC;
  SIGNAL or_2714_nl : STD_LOGIC;
  SIGNAL nand_58_nl : STD_LOGIC;
  SIGNAL mux_2766_nl : STD_LOGIC;
  SIGNAL mux_2765_nl : STD_LOGIC;
  SIGNAL mux_2764_nl : STD_LOGIC;
  SIGNAL nor_680_nl : STD_LOGIC;
  SIGNAL mux_2763_nl : STD_LOGIC;
  SIGNAL mux_2762_nl : STD_LOGIC;
  SIGNAL or_2708_nl : STD_LOGIC;
  SIGNAL nor_681_nl : STD_LOGIC;
  SIGNAL mux_2761_nl : STD_LOGIC;
  SIGNAL or_2702_nl : STD_LOGIC;
  SIGNAL and_451_nl : STD_LOGIC;
  SIGNAL mux_2759_nl : STD_LOGIC;
  SIGNAL nor_682_nl : STD_LOGIC;
  SIGNAL mux_2758_nl : STD_LOGIC;
  SIGNAL nor_683_nl : STD_LOGIC;
  SIGNAL nor_684_nl : STD_LOGIC;
  SIGNAL mux_2743_nl : STD_LOGIC;
  SIGNAL nor_685_nl : STD_LOGIC;
  SIGNAL nor_686_nl : STD_LOGIC;
  SIGNAL and_312_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_29_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_30_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_and_277_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_932_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_934_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_and_1_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_936_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_and_2_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_and_3_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_and_4_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_930_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_and_5_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_and_6_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_and_7_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_and_8_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_and_9_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_and_10_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_and_11_nl : STD_LOGIC;
  SIGNAL mux_129_nl : STD_LOGIC;
  SIGNAL mux_128_nl : STD_LOGIC;
  SIGNAL nand_3_nl : STD_LOGIC;
  SIGNAL mux_127_nl : STD_LOGIC;
  SIGNAL mux_126_nl : STD_LOGIC;
  SIGNAL nand_2_nl : STD_LOGIC;
  SIGNAL or_92_nl : STD_LOGIC;
  SIGNAL mux_124_nl : STD_LOGIC;
  SIGNAL mux_123_nl : STD_LOGIC;
  SIGNAL or_91_nl : STD_LOGIC;
  SIGNAL or_89_nl : STD_LOGIC;
  SIGNAL or_88_nl : STD_LOGIC;
  SIGNAL mux_122_nl : STD_LOGIC;
  SIGNAL mux_121_nl : STD_LOGIC;
  SIGNAL mux_120_nl : STD_LOGIC;
  SIGNAL or_87_nl : STD_LOGIC;
  SIGNAL or_85_nl : STD_LOGIC;
  SIGNAL or_81_nl : STD_LOGIC;
  SIGNAL mux_118_nl : STD_LOGIC;
  SIGNAL mux_117_nl : STD_LOGIC;
  SIGNAL or_79_nl : STD_LOGIC;
  SIGNAL mux_116_nl : STD_LOGIC;
  SIGNAL nand_373_nl : STD_LOGIC;
  SIGNAL mux_2981_nl : STD_LOGIC;
  SIGNAL mux_2980_nl : STD_LOGIC;
  SIGNAL mux_2979_nl : STD_LOGIC;
  SIGNAL mux_2978_nl : STD_LOGIC;
  SIGNAL mux_2977_nl : STD_LOGIC;
  SIGNAL mux_2976_nl : STD_LOGIC;
  SIGNAL mux_2975_nl : STD_LOGIC;
  SIGNAL mux_2974_nl : STD_LOGIC;
  SIGNAL mux_2973_nl : STD_LOGIC;
  SIGNAL mux_2972_nl : STD_LOGIC;
  SIGNAL mux_2971_nl : STD_LOGIC;
  SIGNAL mux_2970_nl : STD_LOGIC;
  SIGNAL mux_2969_nl : STD_LOGIC;
  SIGNAL mux_2968_nl : STD_LOGIC;
  SIGNAL mux_2967_nl : STD_LOGIC;
  SIGNAL mux_2966_nl : STD_LOGIC;
  SIGNAL mux_2965_nl : STD_LOGIC;
  SIGNAL mux_2964_nl : STD_LOGIC;
  SIGNAL mux_2963_nl : STD_LOGIC;
  SIGNAL mux_2962_nl : STD_LOGIC;
  SIGNAL mux_2961_nl : STD_LOGIC;
  SIGNAL mux_2960_nl : STD_LOGIC;
  SIGNAL or_2810_nl : STD_LOGIC;
  SIGNAL mux_2959_nl : STD_LOGIC;
  SIGNAL nand_72_nl : STD_LOGIC;
  SIGNAL mux_2958_nl : STD_LOGIC;
  SIGNAL mux_2957_nl : STD_LOGIC;
  SIGNAL mux_2956_nl : STD_LOGIC;
  SIGNAL mux_2955_nl : STD_LOGIC;
  SIGNAL mux_2954_nl : STD_LOGIC;
  SIGNAL mux_2953_nl : STD_LOGIC;
  SIGNAL mux_2952_nl : STD_LOGIC;
  SIGNAL mux_2951_nl : STD_LOGIC;
  SIGNAL mux_2950_nl : STD_LOGIC;
  SIGNAL mux_2949_nl : STD_LOGIC;
  SIGNAL mux_2948_nl : STD_LOGIC;
  SIGNAL or_2809_nl : STD_LOGIC;
  SIGNAL mux_2947_nl : STD_LOGIC;
  SIGNAL mux_2946_nl : STD_LOGIC;
  SIGNAL mux_2945_nl : STD_LOGIC;
  SIGNAL mux_2944_nl : STD_LOGIC;
  SIGNAL mux_2943_nl : STD_LOGIC;
  SIGNAL mux_2942_nl : STD_LOGIC;
  SIGNAL mux_2941_nl : STD_LOGIC;
  SIGNAL mux_2940_nl : STD_LOGIC;
  SIGNAL mux_2939_nl : STD_LOGIC;
  SIGNAL mux_2938_nl : STD_LOGIC;
  SIGNAL mux_2937_nl : STD_LOGIC;
  SIGNAL mux_2936_nl : STD_LOGIC;
  SIGNAL mux_2935_nl : STD_LOGIC;
  SIGNAL mux_2934_nl : STD_LOGIC;
  SIGNAL mux_2933_nl : STD_LOGIC;
  SIGNAL mux_2932_nl : STD_LOGIC;
  SIGNAL mux_2931_nl : STD_LOGIC;
  SIGNAL mux_2930_nl : STD_LOGIC;
  SIGNAL mux_2929_nl : STD_LOGIC;
  SIGNAL mux_2928_nl : STD_LOGIC;
  SIGNAL or_2807_nl : STD_LOGIC;
  SIGNAL mux_2927_nl : STD_LOGIC;
  SIGNAL mux_2925_nl : STD_LOGIC;
  SIGNAL mux_2924_nl : STD_LOGIC;
  SIGNAL mux_2923_nl : STD_LOGIC;
  SIGNAL mux_2922_nl : STD_LOGIC;
  SIGNAL mux_2921_nl : STD_LOGIC;
  SIGNAL mux_2919_nl : STD_LOGIC;
  SIGNAL mux_2918_nl : STD_LOGIC;
  SIGNAL mux_2917_nl : STD_LOGIC;
  SIGNAL mux_2915_nl : STD_LOGIC;
  SIGNAL mux_2914_nl : STD_LOGIC;
  SIGNAL mux_2913_nl : STD_LOGIC;
  SIGNAL mux_2911_nl : STD_LOGIC;
  SIGNAL mux_2908_nl : STD_LOGIC;
  SIGNAL mux_2907_nl : STD_LOGIC;
  SIGNAL mux_2905_nl : STD_LOGIC;
  SIGNAL mux_2904_nl : STD_LOGIC;
  SIGNAL mux_2903_nl : STD_LOGIC;
  SIGNAL mux_2902_nl : STD_LOGIC;
  SIGNAL mux_2900_nl : STD_LOGIC;
  SIGNAL mux_2899_nl : STD_LOGIC;
  SIGNAL mux_2898_nl : STD_LOGIC;
  SIGNAL mux_2897_nl : STD_LOGIC;
  SIGNAL mux_2896_nl : STD_LOGIC;
  SIGNAL mux_2894_nl : STD_LOGIC;
  SIGNAL mux_2893_nl : STD_LOGIC;
  SIGNAL mux_2892_nl : STD_LOGIC;
  SIGNAL mux_2891_nl : STD_LOGIC;
  SIGNAL mux_2889_nl : STD_LOGIC;
  SIGNAL mux_2887_nl : STD_LOGIC;
  SIGNAL mux_2885_nl : STD_LOGIC;
  SIGNAL mux_2884_nl : STD_LOGIC;
  SIGNAL mux_2883_nl : STD_LOGIC;
  SIGNAL mux_2882_nl : STD_LOGIC;
  SIGNAL mux_2881_nl : STD_LOGIC;
  SIGNAL mux_2877_nl : STD_LOGIC;
  SIGNAL mux_2874_nl : STD_LOGIC;
  SIGNAL mux_2873_nl : STD_LOGIC;
  SIGNAL mux_2872_nl : STD_LOGIC;
  SIGNAL mux_2871_nl : STD_LOGIC;
  SIGNAL mux_2870_nl : STD_LOGIC;
  SIGNAL mux_2869_nl : STD_LOGIC;
  SIGNAL mux_2868_nl : STD_LOGIC;
  SIGNAL mux_2865_nl : STD_LOGIC;
  SIGNAL mux_2864_nl : STD_LOGIC;
  SIGNAL mux_2861_nl : STD_LOGIC;
  SIGNAL mux_2860_nl : STD_LOGIC;
  SIGNAL mux_2859_nl : STD_LOGIC;
  SIGNAL or_2797_nl : STD_LOGIC;
  SIGNAL mux_2857_nl : STD_LOGIC;
  SIGNAL nand_66_nl : STD_LOGIC;
  SIGNAL mux_2855_nl : STD_LOGIC;
  SIGNAL mux_2854_nl : STD_LOGIC;
  SIGNAL mux_2853_nl : STD_LOGIC;
  SIGNAL mux_2852_nl : STD_LOGIC;
  SIGNAL mux_2847_nl : STD_LOGIC;
  SIGNAL mux_2845_nl : STD_LOGIC;
  SIGNAL mux_2842_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_428_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_11_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_and_274_nl : STD_LOGIC;
  SIGNAL mux_3070_nl : STD_LOGIC;
  SIGNAL mux_3069_nl : STD_LOGIC;
  SIGNAL mux_3068_nl : STD_LOGIC;
  SIGNAL mux_3067_nl : STD_LOGIC;
  SIGNAL mux_3066_nl : STD_LOGIC;
  SIGNAL mux_3065_nl : STD_LOGIC;
  SIGNAL or_2881_nl : STD_LOGIC;
  SIGNAL mux_3064_nl : STD_LOGIC;
  SIGNAL mux_3063_nl : STD_LOGIC;
  SIGNAL mux_3062_nl : STD_LOGIC;
  SIGNAL mux_3061_nl : STD_LOGIC;
  SIGNAL mux_3060_nl : STD_LOGIC;
  SIGNAL mux_3059_nl : STD_LOGIC;
  SIGNAL or_449_nl : STD_LOGIC;
  SIGNAL or_2876_nl : STD_LOGIC;
  SIGNAL mux_3058_nl : STD_LOGIC;
  SIGNAL mux_3057_nl : STD_LOGIC;
  SIGNAL mux_3056_nl : STD_LOGIC;
  SIGNAL nor_407_nl : STD_LOGIC;
  SIGNAL mux_3055_nl : STD_LOGIC;
  SIGNAL mux_3054_nl : STD_LOGIC;
  SIGNAL mux_3053_nl : STD_LOGIC;
  SIGNAL mux_3052_nl : STD_LOGIC;
  SIGNAL mux_3051_nl : STD_LOGIC;
  SIGNAL or_439_nl : STD_LOGIC;
  SIGNAL mux_3050_nl : STD_LOGIC;
  SIGNAL mux_3048_nl : STD_LOGIC;
  SIGNAL mux_3047_nl : STD_LOGIC;
  SIGNAL or_2870_nl : STD_LOGIC;
  SIGNAL mux_3046_nl : STD_LOGIC;
  SIGNAL mux_3045_nl : STD_LOGIC;
  SIGNAL mux_3044_nl : STD_LOGIC;
  SIGNAL mux_3043_nl : STD_LOGIC;
  SIGNAL mux_3042_nl : STD_LOGIC;
  SIGNAL mux_3041_nl : STD_LOGIC;
  SIGNAL mux_3040_nl : STD_LOGIC;
  SIGNAL mux_3039_nl : STD_LOGIC;
  SIGNAL mux_3038_nl : STD_LOGIC;
  SIGNAL mux_3036_nl : STD_LOGIC;
  SIGNAL mux_3035_nl : STD_LOGIC;
  SIGNAL mux_3034_nl : STD_LOGIC;
  SIGNAL mux_3033_nl : STD_LOGIC;
  SIGNAL mux_3030_nl : STD_LOGIC;
  SIGNAL or_2866_nl : STD_LOGIC;
  SIGNAL or_2865_nl : STD_LOGIC;
  SIGNAL mux_3029_nl : STD_LOGIC;
  SIGNAL mux_3028_nl : STD_LOGIC;
  SIGNAL mux_3027_nl : STD_LOGIC;
  SIGNAL mux_3026_nl : STD_LOGIC;
  SIGNAL mux_3025_nl : STD_LOGIC;
  SIGNAL mux_3023_nl : STD_LOGIC;
  SIGNAL or_2859_nl : STD_LOGIC;
  SIGNAL mux_3021_nl : STD_LOGIC;
  SIGNAL mux_3020_nl : STD_LOGIC;
  SIGNAL mux_3019_nl : STD_LOGIC;
  SIGNAL mux_3018_nl : STD_LOGIC;
  SIGNAL mux_3017_nl : STD_LOGIC;
  SIGNAL mux_3016_nl : STD_LOGIC;
  SIGNAL mux_3015_nl : STD_LOGIC;
  SIGNAL mux_3013_nl : STD_LOGIC;
  SIGNAL or_2851_nl : STD_LOGIC;
  SIGNAL mux_3012_nl : STD_LOGIC;
  SIGNAL mux_3011_nl : STD_LOGIC;
  SIGNAL mux_3010_nl : STD_LOGIC;
  SIGNAL mux_3009_nl : STD_LOGIC;
  SIGNAL mux_3005_nl : STD_LOGIC;
  SIGNAL or_2846_nl : STD_LOGIC;
  SIGNAL mux_2989_nl : STD_LOGIC;
  SIGNAL or_3440_nl : STD_LOGIC;
  SIGNAL mux_2988_nl : STD_LOGIC;
  SIGNAL or_2821_nl : STD_LOGIC;
  SIGNAL mux_2987_nl : STD_LOGIC;
  SIGNAL nand_74_nl : STD_LOGIC;
  SIGNAL mux_2986_nl : STD_LOGIC;
  SIGNAL nor_671_nl : STD_LOGIC;
  SIGNAL nor_672_nl : STD_LOGIC;
  SIGNAL or_2818_nl : STD_LOGIC;
  SIGNAL mux_2985_nl : STD_LOGIC;
  SIGNAL or_3441_nl : STD_LOGIC;
  SIGNAL or_3442_nl : STD_LOGIC;
  SIGNAL mux_2984_nl : STD_LOGIC;
  SIGNAL nand_73_nl : STD_LOGIC;
  SIGNAL mux_2983_nl : STD_LOGIC;
  SIGNAL and_447_nl : STD_LOGIC;
  SIGNAL nor_675_nl : STD_LOGIC;
  SIGNAL or_2811_nl : STD_LOGIC;
  SIGNAL mux_3077_nl : STD_LOGIC;
  SIGNAL mux_3076_nl : STD_LOGIC;
  SIGNAL nor_646_nl : STD_LOGIC;
  SIGNAL mux_3075_nl : STD_LOGIC;
  SIGNAL nor_647_nl : STD_LOGIC;
  SIGNAL and_439_nl : STD_LOGIC;
  SIGNAL mux_3074_nl : STD_LOGIC;
  SIGNAL nor_648_nl : STD_LOGIC;
  SIGNAL nor_649_nl : STD_LOGIC;
  SIGNAL mux_3073_nl : STD_LOGIC;
  SIGNAL and_440_nl : STD_LOGIC;
  SIGNAL mux_3072_nl : STD_LOGIC;
  SIGNAL nor_650_nl : STD_LOGIC;
  SIGNAL mux_3071_nl : STD_LOGIC;
  SIGNAL nor_651_nl : STD_LOGIC;
  SIGNAL nor_652_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_17_nl : STD_LOGIC;
  SIGNAL or_2962_nl : STD_LOGIC;
  SIGNAL or_2961_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_1_acc_8_nl : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mux_3288_nl : STD_LOGIC;
  SIGNAL mux_3287_nl : STD_LOGIC;
  SIGNAL mux_3286_nl : STD_LOGIC;
  SIGNAL mux_3285_nl : STD_LOGIC;
  SIGNAL nor_631_nl : STD_LOGIC;
  SIGNAL nor_632_nl : STD_LOGIC;
  SIGNAL mux_3284_nl : STD_LOGIC;
  SIGNAL and_417_nl : STD_LOGIC;
  SIGNAL nor_633_nl : STD_LOGIC;
  SIGNAL mux_3280_nl : STD_LOGIC;
  SIGNAL or_2959_nl : STD_LOGIC;
  SIGNAL mux_3279_nl : STD_LOGIC;
  SIGNAL or_2958_nl : STD_LOGIC;
  SIGNAL or_2957_nl : STD_LOGIC;
  SIGNAL mux_3278_nl : STD_LOGIC;
  SIGNAL or_2954_nl : STD_LOGIC;
  SIGNAL mux_3277_nl : STD_LOGIC;
  SIGNAL mux_3276_nl : STD_LOGIC;
  SIGNAL and_418_nl : STD_LOGIC;
  SIGNAL nor_634_nl : STD_LOGIC;
  SIGNAL nor_635_nl : STD_LOGIC;
  SIGNAL mux_3275_nl : STD_LOGIC;
  SIGNAL nand_92_nl : STD_LOGIC;
  SIGNAL or_2945_nl : STD_LOGIC;
  SIGNAL mux_3273_nl : STD_LOGIC;
  SIGNAL or_2943_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_10_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_1_acc_nl : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL mux_3334_nl : STD_LOGIC;
  SIGNAL mux_3333_nl : STD_LOGIC;
  SIGNAL mux_3332_nl : STD_LOGIC;
  SIGNAL mux_3331_nl : STD_LOGIC;
  SIGNAL mux_3330_nl : STD_LOGIC;
  SIGNAL mux_2642_nl : STD_LOGIC;
  SIGNAL or_2647_nl : STD_LOGIC;
  SIGNAL mux_3327_nl : STD_LOGIC;
  SIGNAL mux_3326_nl : STD_LOGIC;
  SIGNAL or_3032_nl : STD_LOGIC;
  SIGNAL and_410_nl : STD_LOGIC;
  SIGNAL mux_3325_nl : STD_LOGIC;
  SIGNAL and_411_nl : STD_LOGIC;
  SIGNAL mux_3340_nl : STD_LOGIC;
  SIGNAL mux_3339_nl : STD_LOGIC;
  SIGNAL mux_3338_nl : STD_LOGIC;
  SIGNAL mux_3337_nl : STD_LOGIC;
  SIGNAL or_3037_nl : STD_LOGIC;
  SIGNAL mux_3336_nl : STD_LOGIC;
  SIGNAL and_408_nl : STD_LOGIC;
  SIGNAL or_3036_nl : STD_LOGIC;
  SIGNAL mux_3350_nl : STD_LOGIC;
  SIGNAL mux_3349_nl : STD_LOGIC;
  SIGNAL mux_3348_nl : STD_LOGIC;
  SIGNAL mux_3347_nl : STD_LOGIC;
  SIGNAL mux_3346_nl : STD_LOGIC;
  SIGNAL mux_3345_nl : STD_LOGIC;
  SIGNAL mux_3344_nl : STD_LOGIC;
  SIGNAL mux_3355_nl : STD_LOGIC;
  SIGNAL mux_3354_nl : STD_LOGIC;
  SIGNAL mux_3353_nl : STD_LOGIC;
  SIGNAL mux_3351_nl : STD_LOGIC;
  SIGNAL nor_623_nl : STD_LOGIC;
  SIGNAL mux_3359_nl : STD_LOGIC;
  SIGNAL mux_3358_nl : STD_LOGIC;
  SIGNAL mux_3357_nl : STD_LOGIC;
  SIGNAL mux_3356_nl : STD_LOGIC;
  SIGNAL and_401_nl : STD_LOGIC;
  SIGNAL and_402_nl : STD_LOGIC;
  SIGNAL mux_3364_nl : STD_LOGIC;
  SIGNAL mux_3363_nl : STD_LOGIC;
  SIGNAL mux_3362_nl : STD_LOGIC;
  SIGNAL or_3045_nl : STD_LOGIC;
  SIGNAL mux_3360_nl : STD_LOGIC;
  SIGNAL mux_3367_nl : STD_LOGIC;
  SIGNAL mux_3366_nl : STD_LOGIC;
  SIGNAL nor_621_nl : STD_LOGIC;
  SIGNAL mux_3365_nl : STD_LOGIC;
  SIGNAL or_3048_nl : STD_LOGIC;
  SIGNAL and_334_nl : STD_LOGIC;
  SIGNAL mux_3372_nl : STD_LOGIC;
  SIGNAL mux_3371_nl : STD_LOGIC;
  SIGNAL mux_3370_nl : STD_LOGIC;
  SIGNAL nor_619_nl : STD_LOGIC;
  SIGNAL nor_620_nl : STD_LOGIC;
  SIGNAL mux_3369_nl : STD_LOGIC;
  SIGNAL and_337_nl : STD_LOGIC;
  SIGNAL mux_3368_nl : STD_LOGIC;
  SIGNAL and_30_nl : STD_LOGIC;
  SIGNAL mux_3375_nl : STD_LOGIC;
  SIGNAL mux_3374_nl : STD_LOGIC;
  SIGNAL nor_1596_nl : STD_LOGIC;
  SIGNAL mux_3373_nl : STD_LOGIC;
  SIGNAL nor_1597_nl : STD_LOGIC;
  SIGNAL and_749_nl : STD_LOGIC;
  SIGNAL and_750_nl : STD_LOGIC;
  SIGNAL mux_3381_nl : STD_LOGIC;
  SIGNAL mux_3380_nl : STD_LOGIC;
  SIGNAL mux_3379_nl : STD_LOGIC;
  SIGNAL or_3060_nl : STD_LOGIC;
  SIGNAL mux_3377_nl : STD_LOGIC;
  SIGNAL mux_3376_nl : STD_LOGIC;
  SIGNAL or_3058_nl : STD_LOGIC;
  SIGNAL mux_3386_nl : STD_LOGIC;
  SIGNAL mux_3385_nl : STD_LOGIC;
  SIGNAL mux_3384_nl : STD_LOGIC;
  SIGNAL or_3065_nl : STD_LOGIC;
  SIGNAL mux_3383_nl : STD_LOGIC;
  SIGNAL and_394_nl : STD_LOGIC;
  SIGNAL mux_3391_nl : STD_LOGIC;
  SIGNAL mux_3390_nl : STD_LOGIC;
  SIGNAL mux_3389_nl : STD_LOGIC;
  SIGNAL mux_3388_nl : STD_LOGIC;
  SIGNAL nor_615_nl : STD_LOGIC;
  SIGNAL and_391_nl : STD_LOGIC;
  SIGNAL mux_3396_nl : STD_LOGIC;
  SIGNAL mux_3395_nl : STD_LOGIC;
  SIGNAL mux_3394_nl : STD_LOGIC;
  SIGNAL nor_613_nl : STD_LOGIC;
  SIGNAL nor_614_nl : STD_LOGIC;
  SIGNAL mux_3393_nl : STD_LOGIC;
  SIGNAL and_388_nl : STD_LOGIC;
  SIGNAL mux_3400_nl : STD_LOGIC;
  SIGNAL mux_3399_nl : STD_LOGIC;
  SIGNAL nor_611_nl : STD_LOGIC;
  SIGNAL mux_3398_nl : STD_LOGIC;
  SIGNAL nor_612_nl : STD_LOGIC;
  SIGNAL and_384_nl : STD_LOGIC;
  SIGNAL and_386_nl : STD_LOGIC;
  SIGNAL nor_1680_nl : STD_LOGIC;
  SIGNAL mux_3403_nl : STD_LOGIC;
  SIGNAL or_3078_nl : STD_LOGIC;
  SIGNAL and_1162_nl : STD_LOGIC;
  SIGNAL mux_3402_nl : STD_LOGIC;
  SIGNAL or_3076_nl : STD_LOGIC;
  SIGNAL mux_3408_nl : STD_LOGIC;
  SIGNAL mux_3407_nl : STD_LOGIC;
  SIGNAL mux_3406_nl : STD_LOGIC;
  SIGNAL nor_610_nl : STD_LOGIC;
  SIGNAL mux_3405_nl : STD_LOGIC;
  SIGNAL and_341_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_464_nl : STD_LOGIC;
  SIGNAL mux_3521_nl : STD_LOGIC;
  SIGNAL mux_3520_nl : STD_LOGIC;
  SIGNAL mux_3519_nl : STD_LOGIC;
  SIGNAL mux_3518_nl : STD_LOGIC;
  SIGNAL or_3501_nl : STD_LOGIC;
  SIGNAL mux_3517_nl : STD_LOGIC;
  SIGNAL or_3502_nl : STD_LOGIC;
  SIGNAL or_3503_nl : STD_LOGIC;
  SIGNAL or_3504_nl : STD_LOGIC;
  SIGNAL mux_3516_nl : STD_LOGIC;
  SIGNAL mux_3515_nl : STD_LOGIC;
  SIGNAL or_3133_nl : STD_LOGIC;
  SIGNAL mux_3514_nl : STD_LOGIC;
  SIGNAL or_3131_nl : STD_LOGIC;
  SIGNAL or_3130_nl : STD_LOGIC;
  SIGNAL mux_3513_nl : STD_LOGIC;
  SIGNAL mux_3512_nl : STD_LOGIC;
  SIGNAL or_3505_nl : STD_LOGIC;
  SIGNAL nand_412_nl : STD_LOGIC;
  SIGNAL mux_3511_nl : STD_LOGIC;
  SIGNAL nor_600_nl : STD_LOGIC;
  SIGNAL nor_601_nl : STD_LOGIC;
  SIGNAL mux_3510_nl : STD_LOGIC;
  SIGNAL or_3506_nl : STD_LOGIC;
  SIGNAL mux_3509_nl : STD_LOGIC;
  SIGNAL or_3124_nl : STD_LOGIC;
  SIGNAL or_3123_nl : STD_LOGIC;
  SIGNAL nand_413_nl : STD_LOGIC;
  SIGNAL mux_3508_nl : STD_LOGIC;
  SIGNAL or_3120_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_474_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_12_nl : STD_LOGIC;
  SIGNAL mux_3616_nl : STD_LOGIC;
  SIGNAL mux_3615_nl : STD_LOGIC;
  SIGNAL mux_3614_nl : STD_LOGIC;
  SIGNAL mux_3613_nl : STD_LOGIC;
  SIGNAL mux_3612_nl : STD_LOGIC;
  SIGNAL mux_3611_nl : STD_LOGIC;
  SIGNAL mux_3610_nl : STD_LOGIC;
  SIGNAL mux_3609_nl : STD_LOGIC;
  SIGNAL mux_3608_nl : STD_LOGIC;
  SIGNAL mux_3607_nl : STD_LOGIC;
  SIGNAL mux_3606_nl : STD_LOGIC;
  SIGNAL mux_3605_nl : STD_LOGIC;
  SIGNAL mux_3604_nl : STD_LOGIC;
  SIGNAL mux_3603_nl : STD_LOGIC;
  SIGNAL mux_3602_nl : STD_LOGIC;
  SIGNAL mux_3601_nl : STD_LOGIC;
  SIGNAL mux_3600_nl : STD_LOGIC;
  SIGNAL mux_3599_nl : STD_LOGIC;
  SIGNAL or_3192_nl : STD_LOGIC;
  SIGNAL mux_3598_nl : STD_LOGIC;
  SIGNAL mux_3597_nl : STD_LOGIC;
  SIGNAL mux_3596_nl : STD_LOGIC;
  SIGNAL mux_3595_nl : STD_LOGIC;
  SIGNAL mux_493_nl : STD_LOGIC;
  SIGNAL mux_3592_nl : STD_LOGIC;
  SIGNAL mux_3591_nl : STD_LOGIC;
  SIGNAL mux_454_nl : STD_LOGIC;
  SIGNAL mux_3588_nl : STD_LOGIC;
  SIGNAL mux_3586_nl : STD_LOGIC;
  SIGNAL mux_3585_nl : STD_LOGIC;
  SIGNAL mux_3584_nl : STD_LOGIC;
  SIGNAL mux_3583_nl : STD_LOGIC;
  SIGNAL and_364_nl : STD_LOGIC;
  SIGNAL mux_3582_nl : STD_LOGIC;
  SIGNAL mux_3581_nl : STD_LOGIC;
  SIGNAL mux_3580_nl : STD_LOGIC;
  SIGNAL mux_3579_nl : STD_LOGIC;
  SIGNAL mux_3578_nl : STD_LOGIC;
  SIGNAL mux_3572_nl : STD_LOGIC;
  SIGNAL mux_3571_nl : STD_LOGIC;
  SIGNAL mux_3570_nl : STD_LOGIC;
  SIGNAL mux_3569_nl : STD_LOGIC;
  SIGNAL mux_481_nl : STD_LOGIC;
  SIGNAL mux_3566_nl : STD_LOGIC;
  SIGNAL mux_3565_nl : STD_LOGIC;
  SIGNAL mux_3563_nl : STD_LOGIC;
  SIGNAL mux_3562_nl : STD_LOGIC;
  SIGNAL mux_3560_nl : STD_LOGIC;
  SIGNAL mux_3559_nl : STD_LOGIC;
  SIGNAL mux_3558_nl : STD_LOGIC;
  SIGNAL mux_3557_nl : STD_LOGIC;
  SIGNAL and_365_nl : STD_LOGIC;
  SIGNAL mux_3556_nl : STD_LOGIC;
  SIGNAL mux_3554_nl : STD_LOGIC;
  SIGNAL mux_3553_nl : STD_LOGIC;
  SIGNAL mux_3552_nl : STD_LOGIC;
  SIGNAL mux_3548_nl : STD_LOGIC;
  SIGNAL mux_3546_nl : STD_LOGIC;
  SIGNAL or_3177_nl : STD_LOGIC;
  SIGNAL mux_3545_nl : STD_LOGIC;
  SIGNAL mux_3630_nl : STD_LOGIC;
  SIGNAL mux_3629_nl : STD_LOGIC;
  SIGNAL mux_3628_nl : STD_LOGIC;
  SIGNAL nor_565_nl : STD_LOGIC;
  SIGNAL mux_3627_nl : STD_LOGIC;
  SIGNAL nor_566_nl : STD_LOGIC;
  SIGNAL mux_3626_nl : STD_LOGIC;
  SIGNAL or_3213_nl : STD_LOGIC;
  SIGNAL or_3211_nl : STD_LOGIC;
  SIGNAL mux_3625_nl : STD_LOGIC;
  SIGNAL nor_567_nl : STD_LOGIC;
  SIGNAL mux_3624_nl : STD_LOGIC;
  SIGNAL nor_568_nl : STD_LOGIC;
  SIGNAL nor_569_nl : STD_LOGIC;
  SIGNAL mux_3623_nl : STD_LOGIC;
  SIGNAL mux_3622_nl : STD_LOGIC;
  SIGNAL nor_570_nl : STD_LOGIC;
  SIGNAL mux_3621_nl : STD_LOGIC;
  SIGNAL or_3203_nl : STD_LOGIC;
  SIGNAL nor_571_nl : STD_LOGIC;
  SIGNAL mux_3620_nl : STD_LOGIC;
  SIGNAL mux_3619_nl : STD_LOGIC;
  SIGNAL nor_572_nl : STD_LOGIC;
  SIGNAL and_362_nl : STD_LOGIC;
  SIGNAL mux_3617_nl : STD_LOGIC;
  SIGNAL nor_573_nl : STD_LOGIC;
  SIGNAL nor_574_nl : STD_LOGIC;
  SIGNAL nor_575_nl : STD_LOGIC;
  SIGNAL mux_3542_nl : STD_LOGIC;
  SIGNAL nand_411_nl : STD_LOGIC;
  SIGNAL mux_3541_nl : STD_LOGIC;
  SIGNAL nor_578_nl : STD_LOGIC;
  SIGNAL mux_3540_nl : STD_LOGIC;
  SIGNAL or_3171_nl : STD_LOGIC;
  SIGNAL mux_3539_nl : STD_LOGIC;
  SIGNAL nor_579_nl : STD_LOGIC;
  SIGNAL nor_580_nl : STD_LOGIC;
  SIGNAL or_3499_nl : STD_LOGIC;
  SIGNAL mux_3538_nl : STD_LOGIC;
  SIGNAL or_3166_nl : STD_LOGIC;
  SIGNAL mux_3537_nl : STD_LOGIC;
  SIGNAL nand_139_nl : STD_LOGIC;
  SIGNAL nand_104_nl : STD_LOGIC;
  SIGNAL mux_3536_nl : STD_LOGIC;
  SIGNAL nor_582_nl : STD_LOGIC;
  SIGNAL nor_583_nl : STD_LOGIC;
  SIGNAL mux_3636_nl : STD_LOGIC;
  SIGNAL nor_562_nl : STD_LOGIC;
  SIGNAL mux_3635_nl : STD_LOGIC;
  SIGNAL or_3228_nl : STD_LOGIC;
  SIGNAL mux_3634_nl : STD_LOGIC;
  SIGNAL or_3226_nl : STD_LOGIC;
  SIGNAL or_3224_nl : STD_LOGIC;
  SIGNAL and_361_nl : STD_LOGIC;
  SIGNAL mux_3633_nl : STD_LOGIC;
  SIGNAL nor_563_nl : STD_LOGIC;
  SIGNAL nor_564_nl : STD_LOGIC;
  SIGNAL mux_3631_nl : STD_LOGIC;
  SIGNAL or_3217_nl : STD_LOGIC;
  SIGNAL or_3215_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_477_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_14_nl : STD_LOGIC;
  SIGNAL mux_3642_nl : STD_LOGIC;
  SIGNAL mux_3641_nl : STD_LOGIC;
  SIGNAL mux_3640_nl : STD_LOGIC;
  SIGNAL mux_3639_nl : STD_LOGIC;
  SIGNAL mux_3638_nl : STD_LOGIC;
  SIGNAL mux_3637_nl : STD_LOGIC;
  SIGNAL mux_3649_nl : STD_LOGIC;
  SIGNAL or_3497_nl : STD_LOGIC;
  SIGNAL mux_3648_nl : STD_LOGIC;
  SIGNAL or_3241_nl : STD_LOGIC;
  SIGNAL mux_3647_nl : STD_LOGIC;
  SIGNAL or_3240_nl : STD_LOGIC;
  SIGNAL or_3239_nl : STD_LOGIC;
  SIGNAL mux_3646_nl : STD_LOGIC;
  SIGNAL or_3236_nl : STD_LOGIC;
  SIGNAL mux_3645_nl : STD_LOGIC;
  SIGNAL or_3235_nl : STD_LOGIC;
  SIGNAL or_3234_nl : STD_LOGIC;
  SIGNAL mux_3644_nl : STD_LOGIC;
  SIGNAL or_3498_nl : STD_LOGIC;
  SIGNAL nand_410_nl : STD_LOGIC;
  SIGNAL mux_3643_nl : STD_LOGIC;
  SIGNAL nor_560_nl : STD_LOGIC;
  SIGNAL nor_561_nl : STD_LOGIC;
  SIGNAL mux_3656_nl : STD_LOGIC;
  SIGNAL mux_3655_nl : STD_LOGIC;
  SIGNAL nor_555_nl : STD_LOGIC;
  SIGNAL nor_556_nl : STD_LOGIC;
  SIGNAL mux_3654_nl : STD_LOGIC;
  SIGNAL mux_3653_nl : STD_LOGIC;
  SIGNAL or_3253_nl : STD_LOGIC;
  SIGNAL or_3251_nl : STD_LOGIC;
  SIGNAL nor_557_nl : STD_LOGIC;
  SIGNAL mux_3652_nl : STD_LOGIC;
  SIGNAL or_3249_nl : STD_LOGIC;
  SIGNAL mux_3651_nl : STD_LOGIC;
  SIGNAL nand_383_nl : STD_LOGIC;
  SIGNAL or_3246_nl : STD_LOGIC;
  SIGNAL mux_3650_nl : STD_LOGIC;
  SIGNAL or_3244_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_479_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_17_nl : STD_LOGIC;
  SIGNAL mux_3663_nl : STD_LOGIC;
  SIGNAL nand_389_nl : STD_LOGIC;
  SIGNAL mux_3662_nl : STD_LOGIC;
  SIGNAL nor_552_nl : STD_LOGIC;
  SIGNAL mux_3661_nl : STD_LOGIC;
  SIGNAL mux_3660_nl : STD_LOGIC;
  SIGNAL or_3266_nl : STD_LOGIC;
  SIGNAL nand_130_nl : STD_LOGIC;
  SIGNAL nor_553_nl : STD_LOGIC;
  SIGNAL or_3443_nl : STD_LOGIC;
  SIGNAL mux_3659_nl : STD_LOGIC;
  SIGNAL or_3353_nl : STD_LOGIC;
  SIGNAL mux_3658_nl : STD_LOGIC;
  SIGNAL or_3261_nl : STD_LOGIC;
  SIGNAL or_3260_nl : STD_LOGIC;
  SIGNAL mux_3657_nl : STD_LOGIC;
  SIGNAL mux_3670_nl : STD_LOGIC;
  SIGNAL mux_3669_nl : STD_LOGIC;
  SIGNAL nor_547_nl : STD_LOGIC;
  SIGNAL and_357_nl : STD_LOGIC;
  SIGNAL mux_3668_nl : STD_LOGIC;
  SIGNAL nor_548_nl : STD_LOGIC;
  SIGNAL mux_3667_nl : STD_LOGIC;
  SIGNAL or_3282_nl : STD_LOGIC;
  SIGNAL nand_382_nl : STD_LOGIC;
  SIGNAL and_358_nl : STD_LOGIC;
  SIGNAL mux_3666_nl : STD_LOGIC;
  SIGNAL nor_549_nl : STD_LOGIC;
  SIGNAL nor_550_nl : STD_LOGIC;
  SIGNAL nor_551_nl : STD_LOGIC;
  SIGNAL mux_3665_nl : STD_LOGIC;
  SIGNAL or_3274_nl : STD_LOGIC;
  SIGNAL mux_3664_nl : STD_LOGIC;
  SIGNAL or_3273_nl : STD_LOGIC;
  SIGNAL or_3271_nl : STD_LOGIC;
  SIGNAL or_3269_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_480_nl : STD_LOGIC;
  SIGNAL mux_3766_nl : STD_LOGIC;
  SIGNAL mux_3765_nl : STD_LOGIC;
  SIGNAL mux_3764_nl : STD_LOGIC;
  SIGNAL mux_3763_nl : STD_LOGIC;
  SIGNAL mux_3762_nl : STD_LOGIC;
  SIGNAL mux_3761_nl : STD_LOGIC;
  SIGNAL mux_3760_nl : STD_LOGIC;
  SIGNAL mux_3759_nl : STD_LOGIC;
  SIGNAL mux_3758_nl : STD_LOGIC;
  SIGNAL mux_3757_nl : STD_LOGIC;
  SIGNAL mux_3756_nl : STD_LOGIC;
  SIGNAL mux_3755_nl : STD_LOGIC;
  SIGNAL mux_3754_nl : STD_LOGIC;
  SIGNAL mux_3752_nl : STD_LOGIC;
  SIGNAL mux_3751_nl : STD_LOGIC;
  SIGNAL mux_3750_nl : STD_LOGIC;
  SIGNAL or_3302_nl : STD_LOGIC;
  SIGNAL mux_3749_nl : STD_LOGIC;
  SIGNAL mux_3748_nl : STD_LOGIC;
  SIGNAL mux_3747_nl : STD_LOGIC;
  SIGNAL mux_3746_nl : STD_LOGIC;
  SIGNAL mux_3745_nl : STD_LOGIC;
  SIGNAL mux_3744_nl : STD_LOGIC;
  SIGNAL mux_3743_nl : STD_LOGIC;
  SIGNAL nor_546_nl : STD_LOGIC;
  SIGNAL mux_3742_nl : STD_LOGIC;
  SIGNAL mux_3741_nl : STD_LOGIC;
  SIGNAL mux_3740_nl : STD_LOGIC;
  SIGNAL mux_3735_nl : STD_LOGIC;
  SIGNAL mux_3734_nl : STD_LOGIC;
  SIGNAL mux_3733_nl : STD_LOGIC;
  SIGNAL or_3298_nl : STD_LOGIC;
  SIGNAL mux_3732_nl : STD_LOGIC;
  SIGNAL mux_3731_nl : STD_LOGIC;
  SIGNAL and_349_nl : STD_LOGIC;
  SIGNAL mux_3730_nl : STD_LOGIC;
  SIGNAL mux_3729_nl : STD_LOGIC;
  SIGNAL mux_3728_nl : STD_LOGIC;
  SIGNAL mux_3727_nl : STD_LOGIC;
  SIGNAL mux_3726_nl : STD_LOGIC;
  SIGNAL mux_3725_nl : STD_LOGIC;
  SIGNAL mux_3723_nl : STD_LOGIC;
  SIGNAL mux_3722_nl : STD_LOGIC;
  SIGNAL mux_3721_nl : STD_LOGIC;
  SIGNAL mux_3719_nl : STD_LOGIC;
  SIGNAL mux_3717_nl : STD_LOGIC;
  SIGNAL mux_3716_nl : STD_LOGIC;
  SIGNAL mux_3715_nl : STD_LOGIC;
  SIGNAL mux_3714_nl : STD_LOGIC;
  SIGNAL mux_3713_nl : STD_LOGIC;
  SIGNAL mux_3711_nl : STD_LOGIC;
  SIGNAL mux_3710_nl : STD_LOGIC;
  SIGNAL mux_3709_nl : STD_LOGIC;
  SIGNAL mux_3708_nl : STD_LOGIC;
  SIGNAL mux_3707_nl : STD_LOGIC;
  SIGNAL mux_3706_nl : STD_LOGIC;
  SIGNAL or_3295_nl : STD_LOGIC;
  SIGNAL mux_3703_nl : STD_LOGIC;
  SIGNAL mux_3702_nl : STD_LOGIC;
  SIGNAL mux_3699_nl : STD_LOGIC;
  SIGNAL mux_3695_nl : STD_LOGIC;
  SIGNAL mux_3694_nl : STD_LOGIC;
  SIGNAL mux_3693_nl : STD_LOGIC;
  SIGNAL mux_3692_nl : STD_LOGIC;
  SIGNAL mux_3690_nl : STD_LOGIC;
  SIGNAL mux_3689_nl : STD_LOGIC;
  SIGNAL mux_3688_nl : STD_LOGIC;
  SIGNAL mux_3687_nl : STD_LOGIC;
  SIGNAL nand_380_nl : STD_LOGIC;
  SIGNAL mux_3686_nl : STD_LOGIC;
  SIGNAL mux_3685_nl : STD_LOGIC;
  SIGNAL mux_3684_nl : STD_LOGIC;
  SIGNAL mux_3683_nl : STD_LOGIC;
  SIGNAL mux_3682_nl : STD_LOGIC;
  SIGNAL mux_3680_nl : STD_LOGIC;
  SIGNAL mux_3678_nl : STD_LOGIC;
  SIGNAL nor_527_nl : STD_LOGIC;
  SIGNAL mux_3677_nl : STD_LOGIC;
  SIGNAL mux_3676_nl : STD_LOGIC;
  SIGNAL mux_3675_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_28_nl : STD_LOGIC;
  SIGNAL or_18_nl : STD_LOGIC;
  SIGNAL or_84_nl : STD_LOGIC;
  SIGNAL or_83_nl : STD_LOGIC;
  SIGNAL or_108_nl : STD_LOGIC;
  SIGNAL mux_1078_nl : STD_LOGIC;
  SIGNAL mux_1077_nl : STD_LOGIC;
  SIGNAL or_3394_nl : STD_LOGIC;
  SIGNAL or_510_nl : STD_LOGIC;
  SIGNAL mux_1081_nl : STD_LOGIC;
  SIGNAL or_508_nl : STD_LOGIC;
  SIGNAL or_580_nl : STD_LOGIC;
  SIGNAL or_579_nl : STD_LOGIC;
  SIGNAL or_691_nl : STD_LOGIC;
  SIGNAL or_690_nl : STD_LOGIC;
  SIGNAL or_802_nl : STD_LOGIC;
  SIGNAL or_801_nl : STD_LOGIC;
  SIGNAL or_912_nl : STD_LOGIC;
  SIGNAL or_911_nl : STD_LOGIC;
  SIGNAL or_1022_nl : STD_LOGIC;
  SIGNAL or_1021_nl : STD_LOGIC;
  SIGNAL or_1133_nl : STD_LOGIC;
  SIGNAL or_1132_nl : STD_LOGIC;
  SIGNAL or_1244_nl : STD_LOGIC;
  SIGNAL or_1243_nl : STD_LOGIC;
  SIGNAL or_1354_nl : STD_LOGIC;
  SIGNAL or_1353_nl : STD_LOGIC;
  SIGNAL or_1464_nl : STD_LOGIC;
  SIGNAL or_1463_nl : STD_LOGIC;
  SIGNAL or_1575_nl : STD_LOGIC;
  SIGNAL or_1574_nl : STD_LOGIC;
  SIGNAL or_1686_nl : STD_LOGIC;
  SIGNAL or_1685_nl : STD_LOGIC;
  SIGNAL or_1796_nl : STD_LOGIC;
  SIGNAL or_1795_nl : STD_LOGIC;
  SIGNAL or_1906_nl : STD_LOGIC;
  SIGNAL or_1905_nl : STD_LOGIC;
  SIGNAL or_2017_nl : STD_LOGIC;
  SIGNAL or_2016_nl : STD_LOGIC;
  SIGNAL or_2128_nl : STD_LOGIC;
  SIGNAL or_2127_nl : STD_LOGIC;
  SIGNAL nand_225_nl : STD_LOGIC;
  SIGNAL or_2237_nl : STD_LOGIC;
  SIGNAL mux_2175_nl : STD_LOGIC;
  SIGNAL mux_2234_nl : STD_LOGIC;
  SIGNAL mux_2239_nl : STD_LOGIC;
  SIGNAL nand_188_nl : STD_LOGIC;
  SIGNAL or_2447_nl : STD_LOGIC;
  SIGNAL mux_2352_nl : STD_LOGIC;
  SIGNAL or_2448_nl : STD_LOGIC;
  SIGNAL or_2451_nl : STD_LOGIC;
  SIGNAL or_2457_nl : STD_LOGIC;
  SIGNAL or_2459_nl : STD_LOGIC;
  SIGNAL mux_2375_nl : STD_LOGIC;
  SIGNAL or_2462_nl : STD_LOGIC;
  SIGNAL mux_2385_nl : STD_LOGIC;
  SIGNAL mux_2388_nl : STD_LOGIC;
  SIGNAL mux_2387_nl : STD_LOGIC;
  SIGNAL or_2475_nl : STD_LOGIC;
  SIGNAL or_2474_nl : STD_LOGIC;
  SIGNAL mux_2431_nl : STD_LOGIC;
  SIGNAL nor_741_nl : STD_LOGIC;
  SIGNAL mux_2430_nl : STD_LOGIC;
  SIGNAL or_2488_nl : STD_LOGIC;
  SIGNAL or_2487_nl : STD_LOGIC;
  SIGNAL mux_2429_nl : STD_LOGIC;
  SIGNAL mux_2428_nl : STD_LOGIC;
  SIGNAL nor_742_nl : STD_LOGIC;
  SIGNAL mux_2427_nl : STD_LOGIC;
  SIGNAL or_2484_nl : STD_LOGIC;
  SIGNAL nand_182_nl : STD_LOGIC;
  SIGNAL nor_743_nl : STD_LOGIC;
  SIGNAL mux_2426_nl : STD_LOGIC;
  SIGNAL nor_744_nl : STD_LOGIC;
  SIGNAL mux_2425_nl : STD_LOGIC;
  SIGNAL or_2479_nl : STD_LOGIC;
  SIGNAL or_2478_nl : STD_LOGIC;
  SIGNAL nor_745_nl : STD_LOGIC;
  SIGNAL mux_2423_nl : STD_LOGIC;
  SIGNAL mux_2422_nl : STD_LOGIC;
  SIGNAL mux_2421_nl : STD_LOGIC;
  SIGNAL nor_746_nl : STD_LOGIC;
  SIGNAL nor_747_nl : STD_LOGIC;
  SIGNAL mux_2420_nl : STD_LOGIC;
  SIGNAL nor_748_nl : STD_LOGIC;
  SIGNAL nor_749_nl : STD_LOGIC;
  SIGNAL mux_2419_nl : STD_LOGIC;
  SIGNAL nand_388_nl : STD_LOGIC;
  SIGNAL or_2465_nl : STD_LOGIC;
  SIGNAL nor_750_nl : STD_LOGIC;
  SIGNAL mux_2445_nl : STD_LOGIC;
  SIGNAL mux_2444_nl : STD_LOGIC;
  SIGNAL mux_2443_nl : STD_LOGIC;
  SIGNAL nor_729_nl : STD_LOGIC;
  SIGNAL mux_2442_nl : STD_LOGIC;
  SIGNAL or_2512_nl : STD_LOGIC;
  SIGNAL nor_730_nl : STD_LOGIC;
  SIGNAL nor_1628_nl : STD_LOGIC;
  SIGNAL mux_2441_nl : STD_LOGIC;
  SIGNAL nor_732_nl : STD_LOGIC;
  SIGNAL mux_2440_nl : STD_LOGIC;
  SIGNAL nor_733_nl : STD_LOGIC;
  SIGNAL mux_2439_nl : STD_LOGIC;
  SIGNAL nor_734_nl : STD_LOGIC;
  SIGNAL nor_735_nl : STD_LOGIC;
  SIGNAL mux_2438_nl : STD_LOGIC;
  SIGNAL mux_2437_nl : STD_LOGIC;
  SIGNAL nor_736_nl : STD_LOGIC;
  SIGNAL mux_2436_nl : STD_LOGIC;
  SIGNAL mux_2435_nl : STD_LOGIC;
  SIGNAL nor_737_nl : STD_LOGIC;
  SIGNAL nor_738_nl : STD_LOGIC;
  SIGNAL nor_739_nl : STD_LOGIC;
  SIGNAL nor_740_nl : STD_LOGIC;
  SIGNAL mux_2434_nl : STD_LOGIC;
  SIGNAL or_2495_nl : STD_LOGIC;
  SIGNAL mux_2433_nl : STD_LOGIC;
  SIGNAL or_2494_nl : STD_LOGIC;
  SIGNAL or_2490_nl : STD_LOGIC;
  SIGNAL mux_2448_nl : STD_LOGIC;
  SIGNAL mux_2447_nl : STD_LOGIC;
  SIGNAL nor_1612_nl : STD_LOGIC;
  SIGNAL mux_2453_nl : STD_LOGIC;
  SIGNAL nor_726_nl : STD_LOGIC;
  SIGNAL nor_727_nl : STD_LOGIC;
  SIGNAL mux_2681_nl : STD_LOGIC;
  SIGNAL mux_2708_nl : STD_LOGIC;
  SIGNAL nor_1575_nl : STD_LOGIC;
  SIGNAL or_2678_nl : STD_LOGIC;
  SIGNAL or_2677_nl : STD_LOGIC;
  SIGNAL mux_2756_nl : STD_LOGIC;
  SIGNAL or_2696_nl : STD_LOGIC;
  SIGNAL mux_2755_nl : STD_LOGIC;
  SIGNAL or_2695_nl : STD_LOGIC;
  SIGNAL mux_2754_nl : STD_LOGIC;
  SIGNAL or_2694_nl : STD_LOGIC;
  SIGNAL or_2693_nl : STD_LOGIC;
  SIGNAL mux_2753_nl : STD_LOGIC;
  SIGNAL mux_2752_nl : STD_LOGIC;
  SIGNAL or_2690_nl : STD_LOGIC;
  SIGNAL mux_2751_nl : STD_LOGIC;
  SIGNAL mux_2750_nl : STD_LOGIC;
  SIGNAL or_2689_nl : STD_LOGIC;
  SIGNAL or_2687_nl : STD_LOGIC;
  SIGNAL mux_2749_nl : STD_LOGIC;
  SIGNAL or_2686_nl : STD_LOGIC;
  SIGNAL or_2684_nl : STD_LOGIC;
  SIGNAL or_2682_nl : STD_LOGIC;
  SIGNAL mux_2748_nl : STD_LOGIC;
  SIGNAL mux_2747_nl : STD_LOGIC;
  SIGNAL or_2681_nl : STD_LOGIC;
  SIGNAL mux_2746_nl : STD_LOGIC;
  SIGNAL or_2676_nl : STD_LOGIC;
  SIGNAL mux_2744_nl : STD_LOGIC;
  SIGNAL or_2675_nl : STD_LOGIC;
  SIGNAL or_2674_nl : STD_LOGIC;
  SIGNAL or_2705_nl : STD_LOGIC;
  SIGNAL or_2704_nl : STD_LOGIC;
  SIGNAL mux_2839_nl : STD_LOGIC;
  SIGNAL mux_2838_nl : STD_LOGIC;
  SIGNAL mux_2837_nl : STD_LOGIC;
  SIGNAL or_2785_nl : STD_LOGIC;
  SIGNAL mux_2836_nl : STD_LOGIC;
  SIGNAL or_2784_nl : STD_LOGIC;
  SIGNAL mux_2835_nl : STD_LOGIC;
  SIGNAL mux_2834_nl : STD_LOGIC;
  SIGNAL mux_2833_nl : STD_LOGIC;
  SIGNAL mux_2832_nl : STD_LOGIC;
  SIGNAL mux_2831_nl : STD_LOGIC;
  SIGNAL mux_2830_nl : STD_LOGIC;
  SIGNAL nand_65_nl : STD_LOGIC;
  SIGNAL mux_2829_nl : STD_LOGIC;
  SIGNAL nand_394_nl : STD_LOGIC;
  SIGNAL mux_2828_nl : STD_LOGIC;
  SIGNAL mux_2827_nl : STD_LOGIC;
  SIGNAL or_2780_nl : STD_LOGIC;
  SIGNAL mux_2826_nl : STD_LOGIC;
  SIGNAL mux_2825_nl : STD_LOGIC;
  SIGNAL mux_2824_nl : STD_LOGIC;
  SIGNAL or_2778_nl : STD_LOGIC;
  SIGNAL mux_2823_nl : STD_LOGIC;
  SIGNAL mux_2822_nl : STD_LOGIC;
  SIGNAL mux_2821_nl : STD_LOGIC;
  SIGNAL mux_2820_nl : STD_LOGIC;
  SIGNAL or_2776_nl : STD_LOGIC;
  SIGNAL mux_2819_nl : STD_LOGIC;
  SIGNAL mux_2818_nl : STD_LOGIC;
  SIGNAL mux_2817_nl : STD_LOGIC;
  SIGNAL or_2775_nl : STD_LOGIC;
  SIGNAL mux_2816_nl : STD_LOGIC;
  SIGNAL or_2774_nl : STD_LOGIC;
  SIGNAL nand_64_nl : STD_LOGIC;
  SIGNAL mux_2815_nl : STD_LOGIC;
  SIGNAL mux_2814_nl : STD_LOGIC;
  SIGNAL mux_2813_nl : STD_LOGIC;
  SIGNAL or_2771_nl : STD_LOGIC;
  SIGNAL mux_2812_nl : STD_LOGIC;
  SIGNAL mux_2811_nl : STD_LOGIC;
  SIGNAL or_2770_nl : STD_LOGIC;
  SIGNAL mux_2810_nl : STD_LOGIC;
  SIGNAL mux_2809_nl : STD_LOGIC;
  SIGNAL mux_2808_nl : STD_LOGIC;
  SIGNAL mux_2807_nl : STD_LOGIC;
  SIGNAL nand_63_nl : STD_LOGIC;
  SIGNAL mux_2806_nl : STD_LOGIC;
  SIGNAL mux_2805_nl : STD_LOGIC;
  SIGNAL mux_2804_nl : STD_LOGIC;
  SIGNAL mux_2803_nl : STD_LOGIC;
  SIGNAL mux_2802_nl : STD_LOGIC;
  SIGNAL mux_2801_nl : STD_LOGIC;
  SIGNAL mux_2800_nl : STD_LOGIC;
  SIGNAL mux_2799_nl : STD_LOGIC;
  SIGNAL or_2759_nl : STD_LOGIC;
  SIGNAL mux_2798_nl : STD_LOGIC;
  SIGNAL mux_2797_nl : STD_LOGIC;
  SIGNAL mux_2795_nl : STD_LOGIC;
  SIGNAL nand_62_nl : STD_LOGIC;
  SIGNAL mux_2794_nl : STD_LOGIC;
  SIGNAL or_2754_nl : STD_LOGIC;
  SIGNAL mux_2793_nl : STD_LOGIC;
  SIGNAL mux_2792_nl : STD_LOGIC;
  SIGNAL mux_2791_nl : STD_LOGIC;
  SIGNAL or_2751_nl : STD_LOGIC;
  SIGNAL mux_2790_nl : STD_LOGIC;
  SIGNAL mux_2789_nl : STD_LOGIC;
  SIGNAL or_2747_nl : STD_LOGIC;
  SIGNAL mux_2788_nl : STD_LOGIC;
  SIGNAL or_2743_nl : STD_LOGIC;
  SIGNAL mux_2787_nl : STD_LOGIC;
  SIGNAL mux_2786_nl : STD_LOGIC;
  SIGNAL or_2740_nl : STD_LOGIC;
  SIGNAL mux_2858_nl : STD_LOGIC;
  SIGNAL mux_2875_nl : STD_LOGIC;
  SIGNAL or_2800_nl : STD_LOGIC;
  SIGNAL mux_2901_nl : STD_LOGIC;
  SIGNAL mux_2909_nl : STD_LOGIC;
  SIGNAL or_2840_nl : STD_LOGIC;
  SIGNAL mux_3002_nl : STD_LOGIC;
  SIGNAL mux_3001_nl : STD_LOGIC;
  SIGNAL nor_661_nl : STD_LOGIC;
  SIGNAL mux_3000_nl : STD_LOGIC;
  SIGNAL nor_662_nl : STD_LOGIC;
  SIGNAL mux_2999_nl : STD_LOGIC;
  SIGNAL or_2842_nl : STD_LOGIC;
  SIGNAL nor_663_nl : STD_LOGIC;
  SIGNAL nor_664_nl : STD_LOGIC;
  SIGNAL mux_2997_nl : STD_LOGIC;
  SIGNAL or_2836_nl : STD_LOGIC;
  SIGNAL or_2831_nl : STD_LOGIC;
  SIGNAL mux_2995_nl : STD_LOGIC;
  SIGNAL mux_2994_nl : STD_LOGIC;
  SIGNAL and_445_nl : STD_LOGIC;
  SIGNAL mux_2993_nl : STD_LOGIC;
  SIGNAL nor_665_nl : STD_LOGIC;
  SIGNAL mux_2992_nl : STD_LOGIC;
  SIGNAL nor_666_nl : STD_LOGIC;
  SIGNAL mux_2991_nl : STD_LOGIC;
  SIGNAL mux_2990_nl : STD_LOGIC;
  SIGNAL and_446_nl : STD_LOGIC;
  SIGNAL nor_668_nl : STD_LOGIC;
  SIGNAL nor_669_nl : STD_LOGIC;
  SIGNAL mux_3799_nl : STD_LOGIC;
  SIGNAL mux_3006_nl : STD_LOGIC;
  SIGNAL or_2848_nl : STD_LOGIC;
  SIGNAL or_2863_nl : STD_LOGIC;
  SIGNAL mux_3031_nl : STD_LOGIC;
  SIGNAL or_3367_nl : STD_LOGIC;
  SIGNAL mux_3321_nl : STD_LOGIC;
  SIGNAL or_3025_nl : STD_LOGIC;
  SIGNAL nand_149_nl : STD_LOGIC;
  SIGNAL mux_3320_nl : STD_LOGIC;
  SIGNAL mux_3319_nl : STD_LOGIC;
  SIGNAL or_3023_nl : STD_LOGIC;
  SIGNAL or_3022_nl : STD_LOGIC;
  SIGNAL mux_3342_nl : STD_LOGIC;
  SIGNAL or_3061_nl : STD_LOGIC;
  SIGNAL or_3087_nl : STD_LOGIC;
  SIGNAL or_12_nl : STD_LOGIC;
  SIGNAL mux_3416_nl : STD_LOGIC;
  SIGNAL mux_3427_nl : STD_LOGIC;
  SIGNAL mux_3426_nl : STD_LOGIC;
  SIGNAL mux_3422_nl : STD_LOGIC;
  SIGNAL mux_3431_nl : STD_LOGIC;
  SIGNAL mux_3430_nl : STD_LOGIC;
  SIGNAL mux_3433_nl : STD_LOGIC;
  SIGNAL mux_3436_nl : STD_LOGIC;
  SIGNAL mux_3452_nl : STD_LOGIC;
  SIGNAL mux_3451_nl : STD_LOGIC;
  SIGNAL mux_3450_nl : STD_LOGIC;
  SIGNAL mux_3449_nl : STD_LOGIC;
  SIGNAL mux_3448_nl : STD_LOGIC;
  SIGNAL mux_3447_nl : STD_LOGIC;
  SIGNAL mux_3446_nl : STD_LOGIC;
  SIGNAL mux_3445_nl : STD_LOGIC;
  SIGNAL mux_3444_nl : STD_LOGIC;
  SIGNAL mux_3443_nl : STD_LOGIC;
  SIGNAL mux_3442_nl : STD_LOGIC;
  SIGNAL mux_3441_nl : STD_LOGIC;
  SIGNAL mux_3440_nl : STD_LOGIC;
  SIGNAL mux_3439_nl : STD_LOGIC;
  SIGNAL mux_3438_nl : STD_LOGIC;
  SIGNAL mux_3413_nl : STD_LOGIC;
  SIGNAL mux_3412_nl : STD_LOGIC;
  SIGNAL or_3090_nl : STD_LOGIC;
  SIGNAL mux_3411_nl : STD_LOGIC;
  SIGNAL or_3088_nl : STD_LOGIC;
  SIGNAL mux_3455_nl : STD_LOGIC;
  SIGNAL mux_3454_nl : STD_LOGIC;
  SIGNAL mux_3460_nl : STD_LOGIC;
  SIGNAL mux_3462_nl : STD_LOGIC;
  SIGNAL mux_3471_nl : STD_LOGIC;
  SIGNAL mux_3470_nl : STD_LOGIC;
  SIGNAL mux_3469_nl : STD_LOGIC;
  SIGNAL mux_3468_nl : STD_LOGIC;
  SIGNAL mux_3467_nl : STD_LOGIC;
  SIGNAL mux_3466_nl : STD_LOGIC;
  SIGNAL mux_3465_nl : STD_LOGIC;
  SIGNAL or_3095_nl : STD_LOGIC;
  SIGNAL mux_3476_nl : STD_LOGIC;
  SIGNAL mux_3475_nl : STD_LOGIC;
  SIGNAL mux_3480_nl : STD_LOGIC;
  SIGNAL mux_3479_nl : STD_LOGIC;
  SIGNAL mux_3478_nl : STD_LOGIC;
  SIGNAL mux_3484_nl : STD_LOGIC;
  SIGNAL mux_3490_nl : STD_LOGIC;
  SIGNAL mux_3489_nl : STD_LOGIC;
  SIGNAL mux_3488_nl : STD_LOGIC;
  SIGNAL mux_3493_nl : STD_LOGIC;
  SIGNAL mux_3492_nl : STD_LOGIC;
  SIGNAL mux_3487_nl : STD_LOGIC;
  SIGNAL mux_3486_nl : STD_LOGIC;
  SIGNAL mux_3483_nl : STD_LOGIC;
  SIGNAL mux_3482_nl : STD_LOGIC;
  SIGNAL mux_3506_nl : STD_LOGIC;
  SIGNAL nor_603_nl : STD_LOGIC;
  SIGNAL mux_3505_nl : STD_LOGIC;
  SIGNAL or_3117_nl : STD_LOGIC;
  SIGNAL mux_3504_nl : STD_LOGIC;
  SIGNAL or_3116_nl : STD_LOGIC;
  SIGNAL or_3115_nl : STD_LOGIC;
  SIGNAL mux_3503_nl : STD_LOGIC;
  SIGNAL and_376_nl : STD_LOGIC;
  SIGNAL mux_3502_nl : STD_LOGIC;
  SIGNAL mux_3501_nl : STD_LOGIC;
  SIGNAL nor_604_nl : STD_LOGIC;
  SIGNAL nor_605_nl : STD_LOGIC;
  SIGNAL mux_3500_nl : STD_LOGIC;
  SIGNAL nor_606_nl : STD_LOGIC;
  SIGNAL nor_607_nl : STD_LOGIC;
  SIGNAL nor_608_nl : STD_LOGIC;
  SIGNAL mux_3499_nl : STD_LOGIC;
  SIGNAL mux_3498_nl : STD_LOGIC;
  SIGNAL or_3104_nl : STD_LOGIC;
  SIGNAL mux_3497_nl : STD_LOGIC;
  SIGNAL or_3099_nl : STD_LOGIC;
  SIGNAL mux_3495_nl : STD_LOGIC;
  SIGNAL or_3098_nl : STD_LOGIC;
  SIGNAL or_3097_nl : STD_LOGIC;
  SIGNAL or_3154_nl : STD_LOGIC;
  SIGNAL mux_3534_nl : STD_LOGIC;
  SIGNAL mux_3533_nl : STD_LOGIC;
  SIGNAL nor_584_nl : STD_LOGIC;
  SIGNAL nor_585_nl : STD_LOGIC;
  SIGNAL mux_3532_nl : STD_LOGIC;
  SIGNAL nand_103_nl : STD_LOGIC;
  SIGNAL or_3157_nl : STD_LOGIC;
  SIGNAL mux_3531_nl : STD_LOGIC;
  SIGNAL and_371_nl : STD_LOGIC;
  SIGNAL mux_3530_nl : STD_LOGIC;
  SIGNAL nor_586_nl : STD_LOGIC;
  SIGNAL nor_587_nl : STD_LOGIC;
  SIGNAL nor_588_nl : STD_LOGIC;
  SIGNAL mux_3528_nl : STD_LOGIC;
  SIGNAL mux_3527_nl : STD_LOGIC;
  SIGNAL and_372_nl : STD_LOGIC;
  SIGNAL mux_3526_nl : STD_LOGIC;
  SIGNAL nor_589_nl : STD_LOGIC;
  SIGNAL and_373_nl : STD_LOGIC;
  SIGNAL mux_3525_nl : STD_LOGIC;
  SIGNAL nor_590_nl : STD_LOGIC;
  SIGNAL mux_3524_nl : STD_LOGIC;
  SIGNAL nor_591_nl : STD_LOGIC;
  SIGNAL nor_593_nl : STD_LOGIC;
  SIGNAL mux_3522_nl : STD_LOGIC;
  SIGNAL or_3142_nl : STD_LOGIC;
  SIGNAL or_3141_nl : STD_LOGIC;
  SIGNAL or_3178_nl : STD_LOGIC;
  SIGNAL mux_460_nl : STD_LOGIC;
  SIGNAL or_3199_nl : STD_LOGIC;
  SIGNAL or_3222_nl : STD_LOGIC;
  SIGNAL or_3221_nl : STD_LOGIC;
  SIGNAL or_127_nl : STD_LOGIC;
  SIGNAL or_134_nl : STD_LOGIC;
  SIGNAL mux_262_nl : STD_LOGIC;
  SIGNAL mux_3738_nl : STD_LOGIC;
  SIGNAL mux_2657_nl : STD_LOGIC;
  SIGNAL mux_2656_nl : STD_LOGIC;
  SIGNAL mux_2655_nl : STD_LOGIC;
  SIGNAL mux_2654_nl : STD_LOGIC;
  SIGNAL nor_693_nl : STD_LOGIC;
  SIGNAL mux_2653_nl : STD_LOGIC;
  SIGNAL and_467_nl : STD_LOGIC;
  SIGNAL STAGE_LOOP_acc_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL and_139_nl : STD_LOGIC;
  SIGNAL mux_1093_nl : STD_LOGIC;
  SIGNAL mux_1092_nl : STD_LOGIC;
  SIGNAL mux_1091_nl : STD_LOGIC;
  SIGNAL or_522_nl : STD_LOGIC;
  SIGNAL or_520_nl : STD_LOGIC;
  SIGNAL mux_1090_nl : STD_LOGIC;
  SIGNAL mux_1089_nl : STD_LOGIC;
  SIGNAL or_518_nl : STD_LOGIC;
  SIGNAL mux_1088_nl : STD_LOGIC;
  SIGNAL or_516_nl : STD_LOGIC;
  SIGNAL mux_1087_nl : STD_LOGIC;
  SIGNAL or_515_nl : STD_LOGIC;
  SIGNAL or_513_nl : STD_LOGIC;
  SIGNAL mux_1086_nl : STD_LOGIC;
  SIGNAL mux_1085_nl : STD_LOGIC;
  SIGNAL mux_1084_nl : STD_LOGIC;
  SIGNAL or_512_nl : STD_LOGIC;
  SIGNAL or_511_nl : STD_LOGIC;
  SIGNAL mux_1083_nl : STD_LOGIC;
  SIGNAL or_506_nl : STD_LOGIC;
  SIGNAL or_504_nl : STD_LOGIC;
  SIGNAL and_144_nl : STD_LOGIC;
  SIGNAL mux_1094_nl : STD_LOGIC;
  SIGNAL nor_1513_nl : STD_LOGIC;
  SIGNAL nor_1514_nl : STD_LOGIC;
  SIGNAL and_153_nl : STD_LOGIC;
  SIGNAL mux_1095_nl : STD_LOGIC;
  SIGNAL nor_1511_nl : STD_LOGIC;
  SIGNAL nor_1512_nl : STD_LOGIC;
  SIGNAL and_162_nl : STD_LOGIC;
  SIGNAL mux_1096_nl : STD_LOGIC;
  SIGNAL nor_1509_nl : STD_LOGIC;
  SIGNAL nor_1510_nl : STD_LOGIC;
  SIGNAL and_170_nl : STD_LOGIC;
  SIGNAL mux_1097_nl : STD_LOGIC;
  SIGNAL and_758_nl : STD_LOGIC;
  SIGNAL nor_1508_nl : STD_LOGIC;
  SIGNAL and_180_nl : STD_LOGIC;
  SIGNAL mux_1098_nl : STD_LOGIC;
  SIGNAL nor_1505_nl : STD_LOGIC;
  SIGNAL nor_1506_nl : STD_LOGIC;
  SIGNAL and_187_nl : STD_LOGIC;
  SIGNAL mux_1099_nl : STD_LOGIC;
  SIGNAL nor_1503_nl : STD_LOGIC;
  SIGNAL nor_1504_nl : STD_LOGIC;
  SIGNAL and_195_nl : STD_LOGIC;
  SIGNAL mux_1100_nl : STD_LOGIC;
  SIGNAL nor_1501_nl : STD_LOGIC;
  SIGNAL nor_1502_nl : STD_LOGIC;
  SIGNAL and_201_nl : STD_LOGIC;
  SIGNAL mux_1101_nl : STD_LOGIC;
  SIGNAL nor_1499_nl : STD_LOGIC;
  SIGNAL nor_1500_nl : STD_LOGIC;
  SIGNAL nor_1625_nl : STD_LOGIC;
  SIGNAL mux_1102_nl : STD_LOGIC;
  SIGNAL or_3445_nl : STD_LOGIC;
  SIGNAL or_3446_nl : STD_LOGIC;
  SIGNAL and_213_nl : STD_LOGIC;
  SIGNAL mux_1103_nl : STD_LOGIC;
  SIGNAL nor_1495_nl : STD_LOGIC;
  SIGNAL nor_1496_nl : STD_LOGIC;
  SIGNAL and_219_nl : STD_LOGIC;
  SIGNAL mux_1104_nl : STD_LOGIC;
  SIGNAL nor_1493_nl : STD_LOGIC;
  SIGNAL nor_1494_nl : STD_LOGIC;
  SIGNAL and_225_nl : STD_LOGIC;
  SIGNAL mux_1105_nl : STD_LOGIC;
  SIGNAL and_760_nl : STD_LOGIC;
  SIGNAL nor_1492_nl : STD_LOGIC;
  SIGNAL and_235_nl : STD_LOGIC;
  SIGNAL mux_1106_nl : STD_LOGIC;
  SIGNAL nor_1489_nl : STD_LOGIC;
  SIGNAL and_748_nl : STD_LOGIC;
  SIGNAL and_241_nl : STD_LOGIC;
  SIGNAL mux_1107_nl : STD_LOGIC;
  SIGNAL and_627_nl : STD_LOGIC;
  SIGNAL nor_1488_nl : STD_LOGIC;
  SIGNAL and_249_nl : STD_LOGIC;
  SIGNAL mux_1108_nl : STD_LOGIC;
  SIGNAL nor_1486_nl : STD_LOGIC;
  SIGNAL nor_1487_nl : STD_LOGIC;
  SIGNAL mux_1138_nl : STD_LOGIC;
  SIGNAL mux_1137_nl : STD_LOGIC;
  SIGNAL mux_1136_nl : STD_LOGIC;
  SIGNAL nor_1471_nl : STD_LOGIC;
  SIGNAL mux_1135_nl : STD_LOGIC;
  SIGNAL mux_1134_nl : STD_LOGIC;
  SIGNAL or_618_nl : STD_LOGIC;
  SIGNAL or_617_nl : STD_LOGIC;
  SIGNAL or_615_nl : STD_LOGIC;
  SIGNAL nor_1472_nl : STD_LOGIC;
  SIGNAL mux_1133_nl : STD_LOGIC;
  SIGNAL nor_1473_nl : STD_LOGIC;
  SIGNAL mux_1132_nl : STD_LOGIC;
  SIGNAL nor_1474_nl : STD_LOGIC;
  SIGNAL mux_1131_nl : STD_LOGIC;
  SIGNAL nor_1475_nl : STD_LOGIC;
  SIGNAL nor_1476_nl : STD_LOGIC;
  SIGNAL mux_1130_nl : STD_LOGIC;
  SIGNAL and_626_nl : STD_LOGIC;
  SIGNAL mux_1129_nl : STD_LOGIC;
  SIGNAL or_606_nl : STD_LOGIC;
  SIGNAL mux_1128_nl : STD_LOGIC;
  SIGNAL or_605_nl : STD_LOGIC;
  SIGNAL mux_1127_nl : STD_LOGIC;
  SIGNAL nor_1477_nl : STD_LOGIC;
  SIGNAL mux_1126_nl : STD_LOGIC;
  SIGNAL or_602_nl : STD_LOGIC;
  SIGNAL mux_1125_nl : STD_LOGIC;
  SIGNAL or_600_nl : STD_LOGIC;
  SIGNAL nor_1478_nl : STD_LOGIC;
  SIGNAL mux_1124_nl : STD_LOGIC;
  SIGNAL mux_1123_nl : STD_LOGIC;
  SIGNAL mux_1122_nl : STD_LOGIC;
  SIGNAL nor_1479_nl : STD_LOGIC;
  SIGNAL mux_1121_nl : STD_LOGIC;
  SIGNAL or_596_nl : STD_LOGIC;
  SIGNAL or_594_nl : STD_LOGIC;
  SIGNAL nor_1480_nl : STD_LOGIC;
  SIGNAL mux_1120_nl : STD_LOGIC;
  SIGNAL mux_1119_nl : STD_LOGIC;
  SIGNAL or_590_nl : STD_LOGIC;
  SIGNAL nor_1481_nl : STD_LOGIC;
  SIGNAL mux_1118_nl : STD_LOGIC;
  SIGNAL mux_1117_nl : STD_LOGIC;
  SIGNAL or_583_nl : STD_LOGIC;
  SIGNAL or_581_nl : STD_LOGIC;
  SIGNAL mux_1115_nl : STD_LOGIC;
  SIGNAL nor_1482_nl : STD_LOGIC;
  SIGNAL mux_1114_nl : STD_LOGIC;
  SIGNAL mux_1113_nl : STD_LOGIC;
  SIGNAL or_576_nl : STD_LOGIC;
  SIGNAL or_574_nl : STD_LOGIC;
  SIGNAL mux_1112_nl : STD_LOGIC;
  SIGNAL or_573_nl : STD_LOGIC;
  SIGNAL or_572_nl : STD_LOGIC;
  SIGNAL mux_1111_nl : STD_LOGIC;
  SIGNAL nor_1483_nl : STD_LOGIC;
  SIGNAL mux_1110_nl : STD_LOGIC;
  SIGNAL nor_1484_nl : STD_LOGIC;
  SIGNAL nor_1485_nl : STD_LOGIC;
  SIGNAL mux_1109_nl : STD_LOGIC;
  SIGNAL or_567_nl : STD_LOGIC;
  SIGNAL or_565_nl : STD_LOGIC;
  SIGNAL mux_1171_nl : STD_LOGIC;
  SIGNAL and_623_nl : STD_LOGIC;
  SIGNAL mux_1170_nl : STD_LOGIC;
  SIGNAL nor_1440_nl : STD_LOGIC;
  SIGNAL mux_1169_nl : STD_LOGIC;
  SIGNAL or_674_nl : STD_LOGIC;
  SIGNAL or_673_nl : STD_LOGIC;
  SIGNAL mux_1168_nl : STD_LOGIC;
  SIGNAL nor_1441_nl : STD_LOGIC;
  SIGNAL mux_1167_nl : STD_LOGIC;
  SIGNAL nor_1442_nl : STD_LOGIC;
  SIGNAL nor_1443_nl : STD_LOGIC;
  SIGNAL mux_1166_nl : STD_LOGIC;
  SIGNAL mux_1165_nl : STD_LOGIC;
  SIGNAL mux_1164_nl : STD_LOGIC;
  SIGNAL nor_1444_nl : STD_LOGIC;
  SIGNAL mux_1163_nl : STD_LOGIC;
  SIGNAL mux_1162_nl : STD_LOGIC;
  SIGNAL nor_1446_nl : STD_LOGIC;
  SIGNAL nor_1447_nl : STD_LOGIC;
  SIGNAL or_660_nl : STD_LOGIC;
  SIGNAL mux_1161_nl : STD_LOGIC;
  SIGNAL nor_1448_nl : STD_LOGIC;
  SIGNAL mux_1160_nl : STD_LOGIC;
  SIGNAL nor_1449_nl : STD_LOGIC;
  SIGNAL nor_1450_nl : STD_LOGIC;
  SIGNAL mux_1159_nl : STD_LOGIC;
  SIGNAL mux_1158_nl : STD_LOGIC;
  SIGNAL nor_1451_nl : STD_LOGIC;
  SIGNAL nor_1452_nl : STD_LOGIC;
  SIGNAL nor_1453_nl : STD_LOGIC;
  SIGNAL mux_1156_nl : STD_LOGIC;
  SIGNAL mux_1155_nl : STD_LOGIC;
  SIGNAL mux_1154_nl : STD_LOGIC;
  SIGNAL mux_1153_nl : STD_LOGIC;
  SIGNAL and_624_nl : STD_LOGIC;
  SIGNAL mux_1152_nl : STD_LOGIC;
  SIGNAL nor_1454_nl : STD_LOGIC;
  SIGNAL nor_1455_nl : STD_LOGIC;
  SIGNAL and_625_nl : STD_LOGIC;
  SIGNAL mux_1151_nl : STD_LOGIC;
  SIGNAL nor_1456_nl : STD_LOGIC;
  SIGNAL nor_1457_nl : STD_LOGIC;
  SIGNAL mux_1150_nl : STD_LOGIC;
  SIGNAL nor_1458_nl : STD_LOGIC;
  SIGNAL nor_1459_nl : STD_LOGIC;
  SIGNAL mux_1148_nl : STD_LOGIC;
  SIGNAL nor_1460_nl : STD_LOGIC;
  SIGNAL mux_1147_nl : STD_LOGIC;
  SIGNAL nor_1461_nl : STD_LOGIC;
  SIGNAL nor_1462_nl : STD_LOGIC;
  SIGNAL mux_1146_nl : STD_LOGIC;
  SIGNAL mux_1145_nl : STD_LOGIC;
  SIGNAL nor_1463_nl : STD_LOGIC;
  SIGNAL nor_1464_nl : STD_LOGIC;
  SIGNAL mux_1144_nl : STD_LOGIC;
  SIGNAL mux_1143_nl : STD_LOGIC;
  SIGNAL mux_1142_nl : STD_LOGIC;
  SIGNAL nor_1465_nl : STD_LOGIC;
  SIGNAL mux_1141_nl : STD_LOGIC;
  SIGNAL nor_1466_nl : STD_LOGIC;
  SIGNAL nor_1467_nl : STD_LOGIC;
  SIGNAL nor_1468_nl : STD_LOGIC;
  SIGNAL mux_1140_nl : STD_LOGIC;
  SIGNAL nor_1469_nl : STD_LOGIC;
  SIGNAL nor_1470_nl : STD_LOGIC;
  SIGNAL mux_1202_nl : STD_LOGIC;
  SIGNAL mux_1201_nl : STD_LOGIC;
  SIGNAL mux_1200_nl : STD_LOGIC;
  SIGNAL nor_1425_nl : STD_LOGIC;
  SIGNAL mux_1199_nl : STD_LOGIC;
  SIGNAL mux_1198_nl : STD_LOGIC;
  SIGNAL or_729_nl : STD_LOGIC;
  SIGNAL or_728_nl : STD_LOGIC;
  SIGNAL or_726_nl : STD_LOGIC;
  SIGNAL nor_1426_nl : STD_LOGIC;
  SIGNAL mux_1197_nl : STD_LOGIC;
  SIGNAL nor_1427_nl : STD_LOGIC;
  SIGNAL mux_1196_nl : STD_LOGIC;
  SIGNAL nor_1428_nl : STD_LOGIC;
  SIGNAL mux_1195_nl : STD_LOGIC;
  SIGNAL nor_1429_nl : STD_LOGIC;
  SIGNAL nor_1430_nl : STD_LOGIC;
  SIGNAL mux_1194_nl : STD_LOGIC;
  SIGNAL and_622_nl : STD_LOGIC;
  SIGNAL mux_1193_nl : STD_LOGIC;
  SIGNAL or_717_nl : STD_LOGIC;
  SIGNAL mux_1192_nl : STD_LOGIC;
  SIGNAL or_716_nl : STD_LOGIC;
  SIGNAL mux_1191_nl : STD_LOGIC;
  SIGNAL nor_1431_nl : STD_LOGIC;
  SIGNAL mux_1190_nl : STD_LOGIC;
  SIGNAL or_713_nl : STD_LOGIC;
  SIGNAL mux_1189_nl : STD_LOGIC;
  SIGNAL or_711_nl : STD_LOGIC;
  SIGNAL nor_1432_nl : STD_LOGIC;
  SIGNAL mux_1188_nl : STD_LOGIC;
  SIGNAL mux_1187_nl : STD_LOGIC;
  SIGNAL mux_1186_nl : STD_LOGIC;
  SIGNAL nor_1433_nl : STD_LOGIC;
  SIGNAL mux_1185_nl : STD_LOGIC;
  SIGNAL or_707_nl : STD_LOGIC;
  SIGNAL or_705_nl : STD_LOGIC;
  SIGNAL nor_1434_nl : STD_LOGIC;
  SIGNAL mux_1184_nl : STD_LOGIC;
  SIGNAL mux_1183_nl : STD_LOGIC;
  SIGNAL or_701_nl : STD_LOGIC;
  SIGNAL nor_1435_nl : STD_LOGIC;
  SIGNAL mux_1182_nl : STD_LOGIC;
  SIGNAL mux_1181_nl : STD_LOGIC;
  SIGNAL or_694_nl : STD_LOGIC;
  SIGNAL or_692_nl : STD_LOGIC;
  SIGNAL mux_1179_nl : STD_LOGIC;
  SIGNAL nor_1436_nl : STD_LOGIC;
  SIGNAL mux_1178_nl : STD_LOGIC;
  SIGNAL mux_1177_nl : STD_LOGIC;
  SIGNAL or_687_nl : STD_LOGIC;
  SIGNAL or_685_nl : STD_LOGIC;
  SIGNAL mux_1176_nl : STD_LOGIC;
  SIGNAL or_684_nl : STD_LOGIC;
  SIGNAL or_683_nl : STD_LOGIC;
  SIGNAL mux_1175_nl : STD_LOGIC;
  SIGNAL nor_1437_nl : STD_LOGIC;
  SIGNAL mux_1174_nl : STD_LOGIC;
  SIGNAL nor_1438_nl : STD_LOGIC;
  SIGNAL nor_1439_nl : STD_LOGIC;
  SIGNAL mux_1173_nl : STD_LOGIC;
  SIGNAL or_678_nl : STD_LOGIC;
  SIGNAL or_676_nl : STD_LOGIC;
  SIGNAL mux_1235_nl : STD_LOGIC;
  SIGNAL and_619_nl : STD_LOGIC;
  SIGNAL mux_1234_nl : STD_LOGIC;
  SIGNAL nor_1394_nl : STD_LOGIC;
  SIGNAL mux_1233_nl : STD_LOGIC;
  SIGNAL or_785_nl : STD_LOGIC;
  SIGNAL or_784_nl : STD_LOGIC;
  SIGNAL mux_1232_nl : STD_LOGIC;
  SIGNAL nor_1395_nl : STD_LOGIC;
  SIGNAL mux_1231_nl : STD_LOGIC;
  SIGNAL nor_1396_nl : STD_LOGIC;
  SIGNAL nor_1397_nl : STD_LOGIC;
  SIGNAL mux_1230_nl : STD_LOGIC;
  SIGNAL mux_1229_nl : STD_LOGIC;
  SIGNAL mux_1228_nl : STD_LOGIC;
  SIGNAL nor_1398_nl : STD_LOGIC;
  SIGNAL mux_1227_nl : STD_LOGIC;
  SIGNAL mux_1226_nl : STD_LOGIC;
  SIGNAL nor_1400_nl : STD_LOGIC;
  SIGNAL nor_1401_nl : STD_LOGIC;
  SIGNAL or_771_nl : STD_LOGIC;
  SIGNAL mux_1225_nl : STD_LOGIC;
  SIGNAL nor_1402_nl : STD_LOGIC;
  SIGNAL mux_1224_nl : STD_LOGIC;
  SIGNAL nor_1403_nl : STD_LOGIC;
  SIGNAL nor_1404_nl : STD_LOGIC;
  SIGNAL mux_1223_nl : STD_LOGIC;
  SIGNAL mux_1222_nl : STD_LOGIC;
  SIGNAL nor_1405_nl : STD_LOGIC;
  SIGNAL nor_1406_nl : STD_LOGIC;
  SIGNAL nor_1407_nl : STD_LOGIC;
  SIGNAL mux_1220_nl : STD_LOGIC;
  SIGNAL mux_1219_nl : STD_LOGIC;
  SIGNAL mux_1218_nl : STD_LOGIC;
  SIGNAL mux_1217_nl : STD_LOGIC;
  SIGNAL and_620_nl : STD_LOGIC;
  SIGNAL mux_1216_nl : STD_LOGIC;
  SIGNAL nor_1408_nl : STD_LOGIC;
  SIGNAL nor_1409_nl : STD_LOGIC;
  SIGNAL and_621_nl : STD_LOGIC;
  SIGNAL mux_1215_nl : STD_LOGIC;
  SIGNAL nor_1410_nl : STD_LOGIC;
  SIGNAL nor_1411_nl : STD_LOGIC;
  SIGNAL mux_1214_nl : STD_LOGIC;
  SIGNAL nor_1412_nl : STD_LOGIC;
  SIGNAL nor_1413_nl : STD_LOGIC;
  SIGNAL mux_1212_nl : STD_LOGIC;
  SIGNAL nor_1414_nl : STD_LOGIC;
  SIGNAL mux_1211_nl : STD_LOGIC;
  SIGNAL nor_1415_nl : STD_LOGIC;
  SIGNAL nor_1416_nl : STD_LOGIC;
  SIGNAL mux_1210_nl : STD_LOGIC;
  SIGNAL mux_1209_nl : STD_LOGIC;
  SIGNAL nor_1417_nl : STD_LOGIC;
  SIGNAL nor_1418_nl : STD_LOGIC;
  SIGNAL mux_1208_nl : STD_LOGIC;
  SIGNAL mux_1207_nl : STD_LOGIC;
  SIGNAL mux_1206_nl : STD_LOGIC;
  SIGNAL nor_1419_nl : STD_LOGIC;
  SIGNAL mux_1205_nl : STD_LOGIC;
  SIGNAL nor_1420_nl : STD_LOGIC;
  SIGNAL nor_1421_nl : STD_LOGIC;
  SIGNAL nor_1422_nl : STD_LOGIC;
  SIGNAL mux_1204_nl : STD_LOGIC;
  SIGNAL nor_1423_nl : STD_LOGIC;
  SIGNAL nor_1424_nl : STD_LOGIC;
  SIGNAL mux_1266_nl : STD_LOGIC;
  SIGNAL mux_1265_nl : STD_LOGIC;
  SIGNAL mux_1264_nl : STD_LOGIC;
  SIGNAL nor_1379_nl : STD_LOGIC;
  SIGNAL mux_1263_nl : STD_LOGIC;
  SIGNAL mux_1262_nl : STD_LOGIC;
  SIGNAL or_839_nl : STD_LOGIC;
  SIGNAL or_838_nl : STD_LOGIC;
  SIGNAL or_836_nl : STD_LOGIC;
  SIGNAL nor_1380_nl : STD_LOGIC;
  SIGNAL mux_1261_nl : STD_LOGIC;
  SIGNAL nor_1381_nl : STD_LOGIC;
  SIGNAL mux_1260_nl : STD_LOGIC;
  SIGNAL nor_1382_nl : STD_LOGIC;
  SIGNAL mux_1259_nl : STD_LOGIC;
  SIGNAL nor_1383_nl : STD_LOGIC;
  SIGNAL nor_1384_nl : STD_LOGIC;
  SIGNAL mux_1258_nl : STD_LOGIC;
  SIGNAL and_618_nl : STD_LOGIC;
  SIGNAL mux_1257_nl : STD_LOGIC;
  SIGNAL or_827_nl : STD_LOGIC;
  SIGNAL mux_1256_nl : STD_LOGIC;
  SIGNAL or_826_nl : STD_LOGIC;
  SIGNAL mux_1255_nl : STD_LOGIC;
  SIGNAL nor_1385_nl : STD_LOGIC;
  SIGNAL mux_1254_nl : STD_LOGIC;
  SIGNAL or_823_nl : STD_LOGIC;
  SIGNAL mux_1253_nl : STD_LOGIC;
  SIGNAL or_821_nl : STD_LOGIC;
  SIGNAL nor_1386_nl : STD_LOGIC;
  SIGNAL mux_1252_nl : STD_LOGIC;
  SIGNAL mux_1251_nl : STD_LOGIC;
  SIGNAL mux_1250_nl : STD_LOGIC;
  SIGNAL nor_1387_nl : STD_LOGIC;
  SIGNAL mux_1249_nl : STD_LOGIC;
  SIGNAL or_817_nl : STD_LOGIC;
  SIGNAL or_815_nl : STD_LOGIC;
  SIGNAL nor_1388_nl : STD_LOGIC;
  SIGNAL mux_1248_nl : STD_LOGIC;
  SIGNAL mux_1247_nl : STD_LOGIC;
  SIGNAL or_809_nl : STD_LOGIC;
  SIGNAL nor_1389_nl : STD_LOGIC;
  SIGNAL mux_1246_nl : STD_LOGIC;
  SIGNAL mux_1245_nl : STD_LOGIC;
  SIGNAL or_805_nl : STD_LOGIC;
  SIGNAL or_803_nl : STD_LOGIC;
  SIGNAL mux_1243_nl : STD_LOGIC;
  SIGNAL nor_1390_nl : STD_LOGIC;
  SIGNAL mux_1242_nl : STD_LOGIC;
  SIGNAL mux_1241_nl : STD_LOGIC;
  SIGNAL or_798_nl : STD_LOGIC;
  SIGNAL or_796_nl : STD_LOGIC;
  SIGNAL mux_1240_nl : STD_LOGIC;
  SIGNAL or_795_nl : STD_LOGIC;
  SIGNAL or_794_nl : STD_LOGIC;
  SIGNAL mux_1239_nl : STD_LOGIC;
  SIGNAL nor_1391_nl : STD_LOGIC;
  SIGNAL mux_1238_nl : STD_LOGIC;
  SIGNAL nor_1392_nl : STD_LOGIC;
  SIGNAL nor_1393_nl : STD_LOGIC;
  SIGNAL mux_1237_nl : STD_LOGIC;
  SIGNAL or_789_nl : STD_LOGIC;
  SIGNAL or_787_nl : STD_LOGIC;
  SIGNAL mux_1299_nl : STD_LOGIC;
  SIGNAL and_615_nl : STD_LOGIC;
  SIGNAL mux_1298_nl : STD_LOGIC;
  SIGNAL nor_1348_nl : STD_LOGIC;
  SIGNAL mux_1297_nl : STD_LOGIC;
  SIGNAL or_895_nl : STD_LOGIC;
  SIGNAL or_894_nl : STD_LOGIC;
  SIGNAL mux_1296_nl : STD_LOGIC;
  SIGNAL nor_1349_nl : STD_LOGIC;
  SIGNAL mux_1295_nl : STD_LOGIC;
  SIGNAL nor_1350_nl : STD_LOGIC;
  SIGNAL nor_1351_nl : STD_LOGIC;
  SIGNAL mux_1294_nl : STD_LOGIC;
  SIGNAL mux_1293_nl : STD_LOGIC;
  SIGNAL mux_1292_nl : STD_LOGIC;
  SIGNAL nor_1352_nl : STD_LOGIC;
  SIGNAL mux_1291_nl : STD_LOGIC;
  SIGNAL mux_1290_nl : STD_LOGIC;
  SIGNAL nor_1354_nl : STD_LOGIC;
  SIGNAL nor_1355_nl : STD_LOGIC;
  SIGNAL or_881_nl : STD_LOGIC;
  SIGNAL mux_1289_nl : STD_LOGIC;
  SIGNAL nor_1356_nl : STD_LOGIC;
  SIGNAL mux_1288_nl : STD_LOGIC;
  SIGNAL nor_1357_nl : STD_LOGIC;
  SIGNAL nor_1358_nl : STD_LOGIC;
  SIGNAL mux_1287_nl : STD_LOGIC;
  SIGNAL mux_1286_nl : STD_LOGIC;
  SIGNAL nor_1359_nl : STD_LOGIC;
  SIGNAL nor_1360_nl : STD_LOGIC;
  SIGNAL nor_1361_nl : STD_LOGIC;
  SIGNAL mux_1284_nl : STD_LOGIC;
  SIGNAL mux_1283_nl : STD_LOGIC;
  SIGNAL mux_1282_nl : STD_LOGIC;
  SIGNAL mux_1281_nl : STD_LOGIC;
  SIGNAL and_616_nl : STD_LOGIC;
  SIGNAL mux_1280_nl : STD_LOGIC;
  SIGNAL nor_1362_nl : STD_LOGIC;
  SIGNAL nor_1363_nl : STD_LOGIC;
  SIGNAL and_617_nl : STD_LOGIC;
  SIGNAL mux_1279_nl : STD_LOGIC;
  SIGNAL nor_1364_nl : STD_LOGIC;
  SIGNAL nor_1365_nl : STD_LOGIC;
  SIGNAL mux_1278_nl : STD_LOGIC;
  SIGNAL nor_1366_nl : STD_LOGIC;
  SIGNAL nor_1367_nl : STD_LOGIC;
  SIGNAL mux_1276_nl : STD_LOGIC;
  SIGNAL nor_1368_nl : STD_LOGIC;
  SIGNAL mux_1275_nl : STD_LOGIC;
  SIGNAL nor_1369_nl : STD_LOGIC;
  SIGNAL nor_1370_nl : STD_LOGIC;
  SIGNAL mux_1274_nl : STD_LOGIC;
  SIGNAL mux_1273_nl : STD_LOGIC;
  SIGNAL nor_1371_nl : STD_LOGIC;
  SIGNAL nor_1372_nl : STD_LOGIC;
  SIGNAL mux_1272_nl : STD_LOGIC;
  SIGNAL mux_1271_nl : STD_LOGIC;
  SIGNAL mux_1270_nl : STD_LOGIC;
  SIGNAL nor_1373_nl : STD_LOGIC;
  SIGNAL mux_1269_nl : STD_LOGIC;
  SIGNAL nor_1374_nl : STD_LOGIC;
  SIGNAL nor_1375_nl : STD_LOGIC;
  SIGNAL nor_1376_nl : STD_LOGIC;
  SIGNAL mux_1268_nl : STD_LOGIC;
  SIGNAL nor_1377_nl : STD_LOGIC;
  SIGNAL nor_1378_nl : STD_LOGIC;
  SIGNAL mux_1330_nl : STD_LOGIC;
  SIGNAL mux_1329_nl : STD_LOGIC;
  SIGNAL mux_1328_nl : STD_LOGIC;
  SIGNAL nor_1333_nl : STD_LOGIC;
  SIGNAL mux_1327_nl : STD_LOGIC;
  SIGNAL mux_1326_nl : STD_LOGIC;
  SIGNAL or_949_nl : STD_LOGIC;
  SIGNAL nand_404_nl : STD_LOGIC;
  SIGNAL or_946_nl : STD_LOGIC;
  SIGNAL nor_1334_nl : STD_LOGIC;
  SIGNAL mux_1325_nl : STD_LOGIC;
  SIGNAL nor_1335_nl : STD_LOGIC;
  SIGNAL mux_1324_nl : STD_LOGIC;
  SIGNAL nor_1336_nl : STD_LOGIC;
  SIGNAL mux_1323_nl : STD_LOGIC;
  SIGNAL nor_1337_nl : STD_LOGIC;
  SIGNAL nor_1338_nl : STD_LOGIC;
  SIGNAL mux_1322_nl : STD_LOGIC;
  SIGNAL and_614_nl : STD_LOGIC;
  SIGNAL mux_1321_nl : STD_LOGIC;
  SIGNAL nand_327_nl : STD_LOGIC;
  SIGNAL mux_1320_nl : STD_LOGIC;
  SIGNAL or_936_nl : STD_LOGIC;
  SIGNAL mux_1319_nl : STD_LOGIC;
  SIGNAL nor_1339_nl : STD_LOGIC;
  SIGNAL mux_1318_nl : STD_LOGIC;
  SIGNAL or_933_nl : STD_LOGIC;
  SIGNAL mux_1317_nl : STD_LOGIC;
  SIGNAL or_931_nl : STD_LOGIC;
  SIGNAL nor_1340_nl : STD_LOGIC;
  SIGNAL mux_1316_nl : STD_LOGIC;
  SIGNAL mux_1315_nl : STD_LOGIC;
  SIGNAL mux_1314_nl : STD_LOGIC;
  SIGNAL nor_1341_nl : STD_LOGIC;
  SIGNAL mux_1313_nl : STD_LOGIC;
  SIGNAL or_927_nl : STD_LOGIC;
  SIGNAL or_925_nl : STD_LOGIC;
  SIGNAL nor_1342_nl : STD_LOGIC;
  SIGNAL mux_1312_nl : STD_LOGIC;
  SIGNAL mux_1311_nl : STD_LOGIC;
  SIGNAL or_919_nl : STD_LOGIC;
  SIGNAL nor_1343_nl : STD_LOGIC;
  SIGNAL mux_1310_nl : STD_LOGIC;
  SIGNAL mux_1309_nl : STD_LOGIC;
  SIGNAL or_915_nl : STD_LOGIC;
  SIGNAL or_913_nl : STD_LOGIC;
  SIGNAL mux_1307_nl : STD_LOGIC;
  SIGNAL nor_1344_nl : STD_LOGIC;
  SIGNAL mux_1306_nl : STD_LOGIC;
  SIGNAL mux_1305_nl : STD_LOGIC;
  SIGNAL or_908_nl : STD_LOGIC;
  SIGNAL or_906_nl : STD_LOGIC;
  SIGNAL mux_1304_nl : STD_LOGIC;
  SIGNAL or_905_nl : STD_LOGIC;
  SIGNAL or_904_nl : STD_LOGIC;
  SIGNAL mux_1303_nl : STD_LOGIC;
  SIGNAL nor_1345_nl : STD_LOGIC;
  SIGNAL mux_1302_nl : STD_LOGIC;
  SIGNAL nor_1346_nl : STD_LOGIC;
  SIGNAL nor_1347_nl : STD_LOGIC;
  SIGNAL mux_1301_nl : STD_LOGIC;
  SIGNAL or_899_nl : STD_LOGIC;
  SIGNAL or_897_nl : STD_LOGIC;
  SIGNAL mux_1363_nl : STD_LOGIC;
  SIGNAL and_611_nl : STD_LOGIC;
  SIGNAL mux_1362_nl : STD_LOGIC;
  SIGNAL nor_1302_nl : STD_LOGIC;
  SIGNAL mux_1361_nl : STD_LOGIC;
  SIGNAL or_1005_nl : STD_LOGIC;
  SIGNAL or_1004_nl : STD_LOGIC;
  SIGNAL mux_1360_nl : STD_LOGIC;
  SIGNAL nor_1303_nl : STD_LOGIC;
  SIGNAL mux_1359_nl : STD_LOGIC;
  SIGNAL nor_1304_nl : STD_LOGIC;
  SIGNAL nor_1305_nl : STD_LOGIC;
  SIGNAL mux_1358_nl : STD_LOGIC;
  SIGNAL mux_1357_nl : STD_LOGIC;
  SIGNAL mux_1356_nl : STD_LOGIC;
  SIGNAL nor_1306_nl : STD_LOGIC;
  SIGNAL mux_1355_nl : STD_LOGIC;
  SIGNAL mux_1354_nl : STD_LOGIC;
  SIGNAL nor_1308_nl : STD_LOGIC;
  SIGNAL nor_1309_nl : STD_LOGIC;
  SIGNAL or_991_nl : STD_LOGIC;
  SIGNAL mux_1353_nl : STD_LOGIC;
  SIGNAL nor_1310_nl : STD_LOGIC;
  SIGNAL mux_1352_nl : STD_LOGIC;
  SIGNAL nor_1311_nl : STD_LOGIC;
  SIGNAL nor_1312_nl : STD_LOGIC;
  SIGNAL mux_1351_nl : STD_LOGIC;
  SIGNAL mux_1350_nl : STD_LOGIC;
  SIGNAL nor_1313_nl : STD_LOGIC;
  SIGNAL nor_1314_nl : STD_LOGIC;
  SIGNAL nor_1315_nl : STD_LOGIC;
  SIGNAL mux_1348_nl : STD_LOGIC;
  SIGNAL mux_1347_nl : STD_LOGIC;
  SIGNAL mux_1346_nl : STD_LOGIC;
  SIGNAL mux_1345_nl : STD_LOGIC;
  SIGNAL and_612_nl : STD_LOGIC;
  SIGNAL mux_1344_nl : STD_LOGIC;
  SIGNAL nor_1316_nl : STD_LOGIC;
  SIGNAL nor_1317_nl : STD_LOGIC;
  SIGNAL and_613_nl : STD_LOGIC;
  SIGNAL mux_1343_nl : STD_LOGIC;
  SIGNAL nor_1318_nl : STD_LOGIC;
  SIGNAL nor_1319_nl : STD_LOGIC;
  SIGNAL mux_1342_nl : STD_LOGIC;
  SIGNAL nor_1320_nl : STD_LOGIC;
  SIGNAL nor_1321_nl : STD_LOGIC;
  SIGNAL mux_1340_nl : STD_LOGIC;
  SIGNAL nor_1322_nl : STD_LOGIC;
  SIGNAL mux_1339_nl : STD_LOGIC;
  SIGNAL nor_1323_nl : STD_LOGIC;
  SIGNAL nor_1324_nl : STD_LOGIC;
  SIGNAL mux_1338_nl : STD_LOGIC;
  SIGNAL mux_1337_nl : STD_LOGIC;
  SIGNAL nor_1325_nl : STD_LOGIC;
  SIGNAL nor_1326_nl : STD_LOGIC;
  SIGNAL mux_1336_nl : STD_LOGIC;
  SIGNAL mux_1335_nl : STD_LOGIC;
  SIGNAL mux_1334_nl : STD_LOGIC;
  SIGNAL nor_1327_nl : STD_LOGIC;
  SIGNAL mux_1333_nl : STD_LOGIC;
  SIGNAL nor_1328_nl : STD_LOGIC;
  SIGNAL nor_1329_nl : STD_LOGIC;
  SIGNAL nor_1330_nl : STD_LOGIC;
  SIGNAL mux_1332_nl : STD_LOGIC;
  SIGNAL nor_1331_nl : STD_LOGIC;
  SIGNAL nor_1332_nl : STD_LOGIC;
  SIGNAL mux_1394_nl : STD_LOGIC;
  SIGNAL mux_1393_nl : STD_LOGIC;
  SIGNAL mux_1392_nl : STD_LOGIC;
  SIGNAL nor_1287_nl : STD_LOGIC;
  SIGNAL mux_1391_nl : STD_LOGIC;
  SIGNAL mux_1390_nl : STD_LOGIC;
  SIGNAL or_1060_nl : STD_LOGIC;
  SIGNAL or_1059_nl : STD_LOGIC;
  SIGNAL or_1057_nl : STD_LOGIC;
  SIGNAL nor_1288_nl : STD_LOGIC;
  SIGNAL mux_1389_nl : STD_LOGIC;
  SIGNAL nor_1289_nl : STD_LOGIC;
  SIGNAL mux_1388_nl : STD_LOGIC;
  SIGNAL nor_1290_nl : STD_LOGIC;
  SIGNAL mux_1387_nl : STD_LOGIC;
  SIGNAL nor_1291_nl : STD_LOGIC;
  SIGNAL nor_1292_nl : STD_LOGIC;
  SIGNAL mux_1386_nl : STD_LOGIC;
  SIGNAL and_610_nl : STD_LOGIC;
  SIGNAL mux_1385_nl : STD_LOGIC;
  SIGNAL or_1048_nl : STD_LOGIC;
  SIGNAL mux_1384_nl : STD_LOGIC;
  SIGNAL or_1047_nl : STD_LOGIC;
  SIGNAL mux_1383_nl : STD_LOGIC;
  SIGNAL nor_1293_nl : STD_LOGIC;
  SIGNAL mux_1382_nl : STD_LOGIC;
  SIGNAL or_1044_nl : STD_LOGIC;
  SIGNAL mux_1381_nl : STD_LOGIC;
  SIGNAL or_1042_nl : STD_LOGIC;
  SIGNAL nor_1294_nl : STD_LOGIC;
  SIGNAL mux_1380_nl : STD_LOGIC;
  SIGNAL mux_1379_nl : STD_LOGIC;
  SIGNAL mux_1378_nl : STD_LOGIC;
  SIGNAL nor_1295_nl : STD_LOGIC;
  SIGNAL mux_1377_nl : STD_LOGIC;
  SIGNAL or_1038_nl : STD_LOGIC;
  SIGNAL or_1036_nl : STD_LOGIC;
  SIGNAL nor_1296_nl : STD_LOGIC;
  SIGNAL mux_1376_nl : STD_LOGIC;
  SIGNAL mux_1375_nl : STD_LOGIC;
  SIGNAL or_1032_nl : STD_LOGIC;
  SIGNAL nor_1297_nl : STD_LOGIC;
  SIGNAL mux_1374_nl : STD_LOGIC;
  SIGNAL mux_1373_nl : STD_LOGIC;
  SIGNAL or_1025_nl : STD_LOGIC;
  SIGNAL or_1023_nl : STD_LOGIC;
  SIGNAL mux_1371_nl : STD_LOGIC;
  SIGNAL nor_1298_nl : STD_LOGIC;
  SIGNAL mux_1370_nl : STD_LOGIC;
  SIGNAL mux_1369_nl : STD_LOGIC;
  SIGNAL or_1018_nl : STD_LOGIC;
  SIGNAL or_1016_nl : STD_LOGIC;
  SIGNAL mux_1368_nl : STD_LOGIC;
  SIGNAL or_1015_nl : STD_LOGIC;
  SIGNAL or_1014_nl : STD_LOGIC;
  SIGNAL mux_1367_nl : STD_LOGIC;
  SIGNAL nor_1299_nl : STD_LOGIC;
  SIGNAL mux_1366_nl : STD_LOGIC;
  SIGNAL nor_1300_nl : STD_LOGIC;
  SIGNAL nor_1301_nl : STD_LOGIC;
  SIGNAL mux_1365_nl : STD_LOGIC;
  SIGNAL or_1009_nl : STD_LOGIC;
  SIGNAL or_1007_nl : STD_LOGIC;
  SIGNAL mux_1427_nl : STD_LOGIC;
  SIGNAL and_607_nl : STD_LOGIC;
  SIGNAL mux_1426_nl : STD_LOGIC;
  SIGNAL nor_1256_nl : STD_LOGIC;
  SIGNAL mux_1425_nl : STD_LOGIC;
  SIGNAL or_1116_nl : STD_LOGIC;
  SIGNAL or_1115_nl : STD_LOGIC;
  SIGNAL mux_1424_nl : STD_LOGIC;
  SIGNAL nor_1257_nl : STD_LOGIC;
  SIGNAL mux_1423_nl : STD_LOGIC;
  SIGNAL nor_1258_nl : STD_LOGIC;
  SIGNAL nor_1259_nl : STD_LOGIC;
  SIGNAL mux_1422_nl : STD_LOGIC;
  SIGNAL mux_1421_nl : STD_LOGIC;
  SIGNAL mux_1420_nl : STD_LOGIC;
  SIGNAL nor_1260_nl : STD_LOGIC;
  SIGNAL mux_1419_nl : STD_LOGIC;
  SIGNAL mux_1418_nl : STD_LOGIC;
  SIGNAL nor_1262_nl : STD_LOGIC;
  SIGNAL nor_1263_nl : STD_LOGIC;
  SIGNAL or_1102_nl : STD_LOGIC;
  SIGNAL mux_1417_nl : STD_LOGIC;
  SIGNAL nor_1264_nl : STD_LOGIC;
  SIGNAL mux_1416_nl : STD_LOGIC;
  SIGNAL nor_1265_nl : STD_LOGIC;
  SIGNAL nor_1266_nl : STD_LOGIC;
  SIGNAL mux_1415_nl : STD_LOGIC;
  SIGNAL mux_1414_nl : STD_LOGIC;
  SIGNAL nor_1267_nl : STD_LOGIC;
  SIGNAL nor_1268_nl : STD_LOGIC;
  SIGNAL nor_1269_nl : STD_LOGIC;
  SIGNAL mux_1412_nl : STD_LOGIC;
  SIGNAL mux_1411_nl : STD_LOGIC;
  SIGNAL mux_1410_nl : STD_LOGIC;
  SIGNAL mux_1409_nl : STD_LOGIC;
  SIGNAL and_608_nl : STD_LOGIC;
  SIGNAL mux_1408_nl : STD_LOGIC;
  SIGNAL nor_1270_nl : STD_LOGIC;
  SIGNAL nor_1271_nl : STD_LOGIC;
  SIGNAL and_609_nl : STD_LOGIC;
  SIGNAL mux_1407_nl : STD_LOGIC;
  SIGNAL nor_1272_nl : STD_LOGIC;
  SIGNAL nor_1273_nl : STD_LOGIC;
  SIGNAL mux_1406_nl : STD_LOGIC;
  SIGNAL nor_1274_nl : STD_LOGIC;
  SIGNAL nor_1275_nl : STD_LOGIC;
  SIGNAL mux_1404_nl : STD_LOGIC;
  SIGNAL nor_1276_nl : STD_LOGIC;
  SIGNAL mux_1403_nl : STD_LOGIC;
  SIGNAL nor_1277_nl : STD_LOGIC;
  SIGNAL nor_1278_nl : STD_LOGIC;
  SIGNAL mux_1402_nl : STD_LOGIC;
  SIGNAL mux_1401_nl : STD_LOGIC;
  SIGNAL nor_1279_nl : STD_LOGIC;
  SIGNAL nor_1280_nl : STD_LOGIC;
  SIGNAL mux_1400_nl : STD_LOGIC;
  SIGNAL mux_1399_nl : STD_LOGIC;
  SIGNAL mux_1398_nl : STD_LOGIC;
  SIGNAL nor_1281_nl : STD_LOGIC;
  SIGNAL mux_1397_nl : STD_LOGIC;
  SIGNAL nor_1282_nl : STD_LOGIC;
  SIGNAL nor_1283_nl : STD_LOGIC;
  SIGNAL nor_1284_nl : STD_LOGIC;
  SIGNAL mux_1396_nl : STD_LOGIC;
  SIGNAL nor_1285_nl : STD_LOGIC;
  SIGNAL nor_1286_nl : STD_LOGIC;
  SIGNAL mux_1458_nl : STD_LOGIC;
  SIGNAL mux_1457_nl : STD_LOGIC;
  SIGNAL mux_1456_nl : STD_LOGIC;
  SIGNAL nor_1241_nl : STD_LOGIC;
  SIGNAL mux_1455_nl : STD_LOGIC;
  SIGNAL mux_1454_nl : STD_LOGIC;
  SIGNAL or_1171_nl : STD_LOGIC;
  SIGNAL nand_403_nl : STD_LOGIC;
  SIGNAL or_1168_nl : STD_LOGIC;
  SIGNAL nor_1242_nl : STD_LOGIC;
  SIGNAL mux_1453_nl : STD_LOGIC;
  SIGNAL nor_1243_nl : STD_LOGIC;
  SIGNAL mux_1452_nl : STD_LOGIC;
  SIGNAL nor_1244_nl : STD_LOGIC;
  SIGNAL mux_1451_nl : STD_LOGIC;
  SIGNAL nor_1245_nl : STD_LOGIC;
  SIGNAL nor_1246_nl : STD_LOGIC;
  SIGNAL mux_1450_nl : STD_LOGIC;
  SIGNAL and_606_nl : STD_LOGIC;
  SIGNAL mux_1449_nl : STD_LOGIC;
  SIGNAL nand_318_nl : STD_LOGIC;
  SIGNAL mux_1448_nl : STD_LOGIC;
  SIGNAL or_1158_nl : STD_LOGIC;
  SIGNAL mux_1447_nl : STD_LOGIC;
  SIGNAL nor_1247_nl : STD_LOGIC;
  SIGNAL mux_1446_nl : STD_LOGIC;
  SIGNAL or_1155_nl : STD_LOGIC;
  SIGNAL mux_1445_nl : STD_LOGIC;
  SIGNAL or_1153_nl : STD_LOGIC;
  SIGNAL nor_1248_nl : STD_LOGIC;
  SIGNAL mux_1444_nl : STD_LOGIC;
  SIGNAL mux_1443_nl : STD_LOGIC;
  SIGNAL mux_1442_nl : STD_LOGIC;
  SIGNAL nor_1249_nl : STD_LOGIC;
  SIGNAL mux_1441_nl : STD_LOGIC;
  SIGNAL or_1149_nl : STD_LOGIC;
  SIGNAL or_1147_nl : STD_LOGIC;
  SIGNAL nor_1250_nl : STD_LOGIC;
  SIGNAL mux_1440_nl : STD_LOGIC;
  SIGNAL mux_1439_nl : STD_LOGIC;
  SIGNAL or_1143_nl : STD_LOGIC;
  SIGNAL nor_1251_nl : STD_LOGIC;
  SIGNAL mux_1438_nl : STD_LOGIC;
  SIGNAL mux_1437_nl : STD_LOGIC;
  SIGNAL or_1136_nl : STD_LOGIC;
  SIGNAL or_1134_nl : STD_LOGIC;
  SIGNAL mux_1435_nl : STD_LOGIC;
  SIGNAL nor_1252_nl : STD_LOGIC;
  SIGNAL mux_1434_nl : STD_LOGIC;
  SIGNAL mux_1433_nl : STD_LOGIC;
  SIGNAL or_1129_nl : STD_LOGIC;
  SIGNAL or_1127_nl : STD_LOGIC;
  SIGNAL mux_1432_nl : STD_LOGIC;
  SIGNAL or_1126_nl : STD_LOGIC;
  SIGNAL or_1125_nl : STD_LOGIC;
  SIGNAL mux_1431_nl : STD_LOGIC;
  SIGNAL nor_1253_nl : STD_LOGIC;
  SIGNAL mux_1430_nl : STD_LOGIC;
  SIGNAL nor_1254_nl : STD_LOGIC;
  SIGNAL nor_1255_nl : STD_LOGIC;
  SIGNAL mux_1429_nl : STD_LOGIC;
  SIGNAL or_1120_nl : STD_LOGIC;
  SIGNAL or_1118_nl : STD_LOGIC;
  SIGNAL mux_1491_nl : STD_LOGIC;
  SIGNAL and_603_nl : STD_LOGIC;
  SIGNAL mux_1490_nl : STD_LOGIC;
  SIGNAL nor_1210_nl : STD_LOGIC;
  SIGNAL mux_1489_nl : STD_LOGIC;
  SIGNAL or_1227_nl : STD_LOGIC;
  SIGNAL or_1226_nl : STD_LOGIC;
  SIGNAL mux_1488_nl : STD_LOGIC;
  SIGNAL nor_1211_nl : STD_LOGIC;
  SIGNAL mux_1487_nl : STD_LOGIC;
  SIGNAL nor_1212_nl : STD_LOGIC;
  SIGNAL nor_1213_nl : STD_LOGIC;
  SIGNAL mux_1486_nl : STD_LOGIC;
  SIGNAL mux_1485_nl : STD_LOGIC;
  SIGNAL mux_1484_nl : STD_LOGIC;
  SIGNAL nor_1214_nl : STD_LOGIC;
  SIGNAL mux_1483_nl : STD_LOGIC;
  SIGNAL mux_1482_nl : STD_LOGIC;
  SIGNAL nor_1216_nl : STD_LOGIC;
  SIGNAL nor_1217_nl : STD_LOGIC;
  SIGNAL or_1213_nl : STD_LOGIC;
  SIGNAL mux_1481_nl : STD_LOGIC;
  SIGNAL nor_1218_nl : STD_LOGIC;
  SIGNAL mux_1480_nl : STD_LOGIC;
  SIGNAL nor_1219_nl : STD_LOGIC;
  SIGNAL nor_1220_nl : STD_LOGIC;
  SIGNAL mux_1479_nl : STD_LOGIC;
  SIGNAL mux_1478_nl : STD_LOGIC;
  SIGNAL nor_1221_nl : STD_LOGIC;
  SIGNAL nor_1222_nl : STD_LOGIC;
  SIGNAL nor_1223_nl : STD_LOGIC;
  SIGNAL mux_1476_nl : STD_LOGIC;
  SIGNAL mux_1475_nl : STD_LOGIC;
  SIGNAL mux_1474_nl : STD_LOGIC;
  SIGNAL mux_1473_nl : STD_LOGIC;
  SIGNAL and_604_nl : STD_LOGIC;
  SIGNAL mux_1472_nl : STD_LOGIC;
  SIGNAL nor_1224_nl : STD_LOGIC;
  SIGNAL nor_1225_nl : STD_LOGIC;
  SIGNAL and_605_nl : STD_LOGIC;
  SIGNAL mux_1471_nl : STD_LOGIC;
  SIGNAL nor_1226_nl : STD_LOGIC;
  SIGNAL nor_1227_nl : STD_LOGIC;
  SIGNAL mux_1470_nl : STD_LOGIC;
  SIGNAL nor_1228_nl : STD_LOGIC;
  SIGNAL nor_1229_nl : STD_LOGIC;
  SIGNAL mux_1468_nl : STD_LOGIC;
  SIGNAL nor_1230_nl : STD_LOGIC;
  SIGNAL mux_1467_nl : STD_LOGIC;
  SIGNAL nor_1231_nl : STD_LOGIC;
  SIGNAL nor_1232_nl : STD_LOGIC;
  SIGNAL mux_1466_nl : STD_LOGIC;
  SIGNAL mux_1465_nl : STD_LOGIC;
  SIGNAL nor_1233_nl : STD_LOGIC;
  SIGNAL nor_1234_nl : STD_LOGIC;
  SIGNAL mux_1464_nl : STD_LOGIC;
  SIGNAL mux_1463_nl : STD_LOGIC;
  SIGNAL mux_1462_nl : STD_LOGIC;
  SIGNAL nor_1235_nl : STD_LOGIC;
  SIGNAL mux_1461_nl : STD_LOGIC;
  SIGNAL nor_1236_nl : STD_LOGIC;
  SIGNAL nor_1237_nl : STD_LOGIC;
  SIGNAL nor_1238_nl : STD_LOGIC;
  SIGNAL mux_1460_nl : STD_LOGIC;
  SIGNAL nor_1239_nl : STD_LOGIC;
  SIGNAL nor_1240_nl : STD_LOGIC;
  SIGNAL mux_1522_nl : STD_LOGIC;
  SIGNAL mux_1521_nl : STD_LOGIC;
  SIGNAL mux_1520_nl : STD_LOGIC;
  SIGNAL nor_1195_nl : STD_LOGIC;
  SIGNAL mux_1519_nl : STD_LOGIC;
  SIGNAL mux_1518_nl : STD_LOGIC;
  SIGNAL or_1281_nl : STD_LOGIC;
  SIGNAL nand_402_nl : STD_LOGIC;
  SIGNAL or_1278_nl : STD_LOGIC;
  SIGNAL nor_1196_nl : STD_LOGIC;
  SIGNAL mux_1517_nl : STD_LOGIC;
  SIGNAL nor_1197_nl : STD_LOGIC;
  SIGNAL mux_1516_nl : STD_LOGIC;
  SIGNAL nor_1198_nl : STD_LOGIC;
  SIGNAL mux_1515_nl : STD_LOGIC;
  SIGNAL nor_1199_nl : STD_LOGIC;
  SIGNAL nor_1200_nl : STD_LOGIC;
  SIGNAL mux_1514_nl : STD_LOGIC;
  SIGNAL and_602_nl : STD_LOGIC;
  SIGNAL mux_1513_nl : STD_LOGIC;
  SIGNAL nand_313_nl : STD_LOGIC;
  SIGNAL mux_1512_nl : STD_LOGIC;
  SIGNAL or_1268_nl : STD_LOGIC;
  SIGNAL mux_1511_nl : STD_LOGIC;
  SIGNAL nor_1201_nl : STD_LOGIC;
  SIGNAL mux_1510_nl : STD_LOGIC;
  SIGNAL or_1265_nl : STD_LOGIC;
  SIGNAL mux_1509_nl : STD_LOGIC;
  SIGNAL or_1263_nl : STD_LOGIC;
  SIGNAL nor_1202_nl : STD_LOGIC;
  SIGNAL mux_1508_nl : STD_LOGIC;
  SIGNAL mux_1507_nl : STD_LOGIC;
  SIGNAL mux_1506_nl : STD_LOGIC;
  SIGNAL nor_1203_nl : STD_LOGIC;
  SIGNAL mux_1505_nl : STD_LOGIC;
  SIGNAL or_1259_nl : STD_LOGIC;
  SIGNAL or_1257_nl : STD_LOGIC;
  SIGNAL nor_1204_nl : STD_LOGIC;
  SIGNAL mux_1504_nl : STD_LOGIC;
  SIGNAL mux_1503_nl : STD_LOGIC;
  SIGNAL or_1251_nl : STD_LOGIC;
  SIGNAL nor_1205_nl : STD_LOGIC;
  SIGNAL mux_1502_nl : STD_LOGIC;
  SIGNAL mux_1501_nl : STD_LOGIC;
  SIGNAL or_1247_nl : STD_LOGIC;
  SIGNAL or_1245_nl : STD_LOGIC;
  SIGNAL mux_1499_nl : STD_LOGIC;
  SIGNAL nor_1206_nl : STD_LOGIC;
  SIGNAL mux_1498_nl : STD_LOGIC;
  SIGNAL mux_1497_nl : STD_LOGIC;
  SIGNAL or_1240_nl : STD_LOGIC;
  SIGNAL or_1238_nl : STD_LOGIC;
  SIGNAL mux_1496_nl : STD_LOGIC;
  SIGNAL or_1237_nl : STD_LOGIC;
  SIGNAL or_1236_nl : STD_LOGIC;
  SIGNAL mux_1495_nl : STD_LOGIC;
  SIGNAL nor_1207_nl : STD_LOGIC;
  SIGNAL mux_1494_nl : STD_LOGIC;
  SIGNAL nor_1208_nl : STD_LOGIC;
  SIGNAL nor_1209_nl : STD_LOGIC;
  SIGNAL mux_1493_nl : STD_LOGIC;
  SIGNAL or_1231_nl : STD_LOGIC;
  SIGNAL or_1229_nl : STD_LOGIC;
  SIGNAL mux_1555_nl : STD_LOGIC;
  SIGNAL and_599_nl : STD_LOGIC;
  SIGNAL mux_1554_nl : STD_LOGIC;
  SIGNAL nor_1164_nl : STD_LOGIC;
  SIGNAL mux_1553_nl : STD_LOGIC;
  SIGNAL or_1337_nl : STD_LOGIC;
  SIGNAL or_1336_nl : STD_LOGIC;
  SIGNAL mux_1552_nl : STD_LOGIC;
  SIGNAL nor_1165_nl : STD_LOGIC;
  SIGNAL mux_1551_nl : STD_LOGIC;
  SIGNAL nor_1166_nl : STD_LOGIC;
  SIGNAL nor_1167_nl : STD_LOGIC;
  SIGNAL mux_1550_nl : STD_LOGIC;
  SIGNAL mux_1549_nl : STD_LOGIC;
  SIGNAL mux_1548_nl : STD_LOGIC;
  SIGNAL nor_1168_nl : STD_LOGIC;
  SIGNAL mux_1547_nl : STD_LOGIC;
  SIGNAL mux_1546_nl : STD_LOGIC;
  SIGNAL nor_1170_nl : STD_LOGIC;
  SIGNAL nor_1171_nl : STD_LOGIC;
  SIGNAL or_1323_nl : STD_LOGIC;
  SIGNAL mux_1545_nl : STD_LOGIC;
  SIGNAL nor_1172_nl : STD_LOGIC;
  SIGNAL mux_1544_nl : STD_LOGIC;
  SIGNAL nor_1173_nl : STD_LOGIC;
  SIGNAL nor_1174_nl : STD_LOGIC;
  SIGNAL mux_1543_nl : STD_LOGIC;
  SIGNAL mux_1542_nl : STD_LOGIC;
  SIGNAL nor_1175_nl : STD_LOGIC;
  SIGNAL nor_1176_nl : STD_LOGIC;
  SIGNAL nor_1177_nl : STD_LOGIC;
  SIGNAL mux_1540_nl : STD_LOGIC;
  SIGNAL mux_1539_nl : STD_LOGIC;
  SIGNAL mux_1538_nl : STD_LOGIC;
  SIGNAL mux_1537_nl : STD_LOGIC;
  SIGNAL and_600_nl : STD_LOGIC;
  SIGNAL mux_1536_nl : STD_LOGIC;
  SIGNAL nor_1178_nl : STD_LOGIC;
  SIGNAL nor_1179_nl : STD_LOGIC;
  SIGNAL and_601_nl : STD_LOGIC;
  SIGNAL mux_1535_nl : STD_LOGIC;
  SIGNAL nor_1180_nl : STD_LOGIC;
  SIGNAL nor_1181_nl : STD_LOGIC;
  SIGNAL mux_1534_nl : STD_LOGIC;
  SIGNAL nor_1182_nl : STD_LOGIC;
  SIGNAL nor_1183_nl : STD_LOGIC;
  SIGNAL mux_1532_nl : STD_LOGIC;
  SIGNAL nor_1184_nl : STD_LOGIC;
  SIGNAL mux_1531_nl : STD_LOGIC;
  SIGNAL nor_1185_nl : STD_LOGIC;
  SIGNAL nor_1186_nl : STD_LOGIC;
  SIGNAL mux_1530_nl : STD_LOGIC;
  SIGNAL mux_1529_nl : STD_LOGIC;
  SIGNAL nor_1187_nl : STD_LOGIC;
  SIGNAL nor_1188_nl : STD_LOGIC;
  SIGNAL mux_1528_nl : STD_LOGIC;
  SIGNAL mux_1527_nl : STD_LOGIC;
  SIGNAL mux_1526_nl : STD_LOGIC;
  SIGNAL nor_1189_nl : STD_LOGIC;
  SIGNAL mux_1525_nl : STD_LOGIC;
  SIGNAL nor_1190_nl : STD_LOGIC;
  SIGNAL nor_1191_nl : STD_LOGIC;
  SIGNAL nor_1192_nl : STD_LOGIC;
  SIGNAL mux_1524_nl : STD_LOGIC;
  SIGNAL nor_1193_nl : STD_LOGIC;
  SIGNAL nor_1194_nl : STD_LOGIC;
  SIGNAL mux_1586_nl : STD_LOGIC;
  SIGNAL mux_1585_nl : STD_LOGIC;
  SIGNAL mux_1584_nl : STD_LOGIC;
  SIGNAL nor_1149_nl : STD_LOGIC;
  SIGNAL mux_1583_nl : STD_LOGIC;
  SIGNAL mux_1582_nl : STD_LOGIC;
  SIGNAL nand_302_nl : STD_LOGIC;
  SIGNAL nand_401_nl : STD_LOGIC;
  SIGNAL or_1388_nl : STD_LOGIC;
  SIGNAL nor_1150_nl : STD_LOGIC;
  SIGNAL mux_1581_nl : STD_LOGIC;
  SIGNAL and_762_nl : STD_LOGIC;
  SIGNAL mux_1580_nl : STD_LOGIC;
  SIGNAL nor_1152_nl : STD_LOGIC;
  SIGNAL mux_1579_nl : STD_LOGIC;
  SIGNAL nor_1153_nl : STD_LOGIC;
  SIGNAL nor_1154_nl : STD_LOGIC;
  SIGNAL mux_1578_nl : STD_LOGIC;
  SIGNAL and_598_nl : STD_LOGIC;
  SIGNAL mux_1577_nl : STD_LOGIC;
  SIGNAL nand_305_nl : STD_LOGIC;
  SIGNAL mux_1576_nl : STD_LOGIC;
  SIGNAL or_1378_nl : STD_LOGIC;
  SIGNAL mux_1575_nl : STD_LOGIC;
  SIGNAL nor_1155_nl : STD_LOGIC;
  SIGNAL mux_1574_nl : STD_LOGIC;
  SIGNAL or_1375_nl : STD_LOGIC;
  SIGNAL mux_1573_nl : STD_LOGIC;
  SIGNAL nand_400_nl : STD_LOGIC;
  SIGNAL nor_1156_nl : STD_LOGIC;
  SIGNAL mux_1572_nl : STD_LOGIC;
  SIGNAL mux_1571_nl : STD_LOGIC;
  SIGNAL mux_1570_nl : STD_LOGIC;
  SIGNAL nor_1157_nl : STD_LOGIC;
  SIGNAL mux_1569_nl : STD_LOGIC;
  SIGNAL or_1369_nl : STD_LOGIC;
  SIGNAL or_1367_nl : STD_LOGIC;
  SIGNAL nor_1158_nl : STD_LOGIC;
  SIGNAL mux_1568_nl : STD_LOGIC;
  SIGNAL mux_1567_nl : STD_LOGIC;
  SIGNAL or_1361_nl : STD_LOGIC;
  SIGNAL nor_1159_nl : STD_LOGIC;
  SIGNAL mux_1566_nl : STD_LOGIC;
  SIGNAL mux_1565_nl : STD_LOGIC;
  SIGNAL or_1357_nl : STD_LOGIC;
  SIGNAL or_1355_nl : STD_LOGIC;
  SIGNAL mux_1563_nl : STD_LOGIC;
  SIGNAL nor_1160_nl : STD_LOGIC;
  SIGNAL mux_1562_nl : STD_LOGIC;
  SIGNAL mux_1561_nl : STD_LOGIC;
  SIGNAL or_1350_nl : STD_LOGIC;
  SIGNAL or_1348_nl : STD_LOGIC;
  SIGNAL mux_1560_nl : STD_LOGIC;
  SIGNAL nand_310_nl : STD_LOGIC;
  SIGNAL or_1346_nl : STD_LOGIC;
  SIGNAL mux_1559_nl : STD_LOGIC;
  SIGNAL nor_1161_nl : STD_LOGIC;
  SIGNAL mux_1558_nl : STD_LOGIC;
  SIGNAL and_763_nl : STD_LOGIC;
  SIGNAL nor_1163_nl : STD_LOGIC;
  SIGNAL mux_1557_nl : STD_LOGIC;
  SIGNAL or_1341_nl : STD_LOGIC;
  SIGNAL or_1339_nl : STD_LOGIC;
  SIGNAL mux_1619_nl : STD_LOGIC;
  SIGNAL and_593_nl : STD_LOGIC;
  SIGNAL mux_1618_nl : STD_LOGIC;
  SIGNAL nor_1120_nl : STD_LOGIC;
  SIGNAL mux_1617_nl : STD_LOGIC;
  SIGNAL or_1447_nl : STD_LOGIC;
  SIGNAL or_1446_nl : STD_LOGIC;
  SIGNAL mux_1616_nl : STD_LOGIC;
  SIGNAL nor_1121_nl : STD_LOGIC;
  SIGNAL mux_1615_nl : STD_LOGIC;
  SIGNAL nor_1122_nl : STD_LOGIC;
  SIGNAL nor_1123_nl : STD_LOGIC;
  SIGNAL mux_1614_nl : STD_LOGIC;
  SIGNAL mux_1613_nl : STD_LOGIC;
  SIGNAL mux_1612_nl : STD_LOGIC;
  SIGNAL nor_1124_nl : STD_LOGIC;
  SIGNAL mux_1611_nl : STD_LOGIC;
  SIGNAL mux_1610_nl : STD_LOGIC;
  SIGNAL nor_1126_nl : STD_LOGIC;
  SIGNAL nor_1127_nl : STD_LOGIC;
  SIGNAL nand_295_nl : STD_LOGIC;
  SIGNAL mux_1609_nl : STD_LOGIC;
  SIGNAL nor_1128_nl : STD_LOGIC;
  SIGNAL mux_1608_nl : STD_LOGIC;
  SIGNAL nor_1129_nl : STD_LOGIC;
  SIGNAL nor_1130_nl : STD_LOGIC;
  SIGNAL mux_1607_nl : STD_LOGIC;
  SIGNAL mux_1606_nl : STD_LOGIC;
  SIGNAL nor_1131_nl : STD_LOGIC;
  SIGNAL nor_1132_nl : STD_LOGIC;
  SIGNAL nor_1133_nl : STD_LOGIC;
  SIGNAL mux_1604_nl : STD_LOGIC;
  SIGNAL mux_1603_nl : STD_LOGIC;
  SIGNAL mux_1602_nl : STD_LOGIC;
  SIGNAL mux_1601_nl : STD_LOGIC;
  SIGNAL and_594_nl : STD_LOGIC;
  SIGNAL mux_1600_nl : STD_LOGIC;
  SIGNAL nor_1134_nl : STD_LOGIC;
  SIGNAL nor_1135_nl : STD_LOGIC;
  SIGNAL and_595_nl : STD_LOGIC;
  SIGNAL mux_1599_nl : STD_LOGIC;
  SIGNAL nor_1136_nl : STD_LOGIC;
  SIGNAL nor_1137_nl : STD_LOGIC;
  SIGNAL mux_1598_nl : STD_LOGIC;
  SIGNAL nor_1138_nl : STD_LOGIC;
  SIGNAL nor_1139_nl : STD_LOGIC;
  SIGNAL mux_1596_nl : STD_LOGIC;
  SIGNAL nor_1140_nl : STD_LOGIC;
  SIGNAL mux_1595_nl : STD_LOGIC;
  SIGNAL nor_1141_nl : STD_LOGIC;
  SIGNAL and_596_nl : STD_LOGIC;
  SIGNAL mux_1594_nl : STD_LOGIC;
  SIGNAL mux_1593_nl : STD_LOGIC;
  SIGNAL nor_1142_nl : STD_LOGIC;
  SIGNAL nor_1143_nl : STD_LOGIC;
  SIGNAL mux_1592_nl : STD_LOGIC;
  SIGNAL mux_1591_nl : STD_LOGIC;
  SIGNAL mux_1590_nl : STD_LOGIC;
  SIGNAL nor_1144_nl : STD_LOGIC;
  SIGNAL mux_1589_nl : STD_LOGIC;
  SIGNAL nor_1145_nl : STD_LOGIC;
  SIGNAL nor_1146_nl : STD_LOGIC;
  SIGNAL nor_1147_nl : STD_LOGIC;
  SIGNAL mux_1588_nl : STD_LOGIC;
  SIGNAL and_597_nl : STD_LOGIC;
  SIGNAL nor_1148_nl : STD_LOGIC;
  SIGNAL mux_1650_nl : STD_LOGIC;
  SIGNAL mux_1649_nl : STD_LOGIC;
  SIGNAL mux_1648_nl : STD_LOGIC;
  SIGNAL nor_1105_nl : STD_LOGIC;
  SIGNAL mux_1647_nl : STD_LOGIC;
  SIGNAL mux_1646_nl : STD_LOGIC;
  SIGNAL or_1502_nl : STD_LOGIC;
  SIGNAL or_1501_nl : STD_LOGIC;
  SIGNAL or_1499_nl : STD_LOGIC;
  SIGNAL nor_1106_nl : STD_LOGIC;
  SIGNAL mux_1645_nl : STD_LOGIC;
  SIGNAL nor_1107_nl : STD_LOGIC;
  SIGNAL mux_1644_nl : STD_LOGIC;
  SIGNAL nor_1108_nl : STD_LOGIC;
  SIGNAL mux_1643_nl : STD_LOGIC;
  SIGNAL nor_1109_nl : STD_LOGIC;
  SIGNAL nor_1110_nl : STD_LOGIC;
  SIGNAL mux_1642_nl : STD_LOGIC;
  SIGNAL and_592_nl : STD_LOGIC;
  SIGNAL mux_1641_nl : STD_LOGIC;
  SIGNAL or_1490_nl : STD_LOGIC;
  SIGNAL mux_1640_nl : STD_LOGIC;
  SIGNAL or_1489_nl : STD_LOGIC;
  SIGNAL mux_1639_nl : STD_LOGIC;
  SIGNAL nor_1111_nl : STD_LOGIC;
  SIGNAL mux_1638_nl : STD_LOGIC;
  SIGNAL or_1486_nl : STD_LOGIC;
  SIGNAL mux_1637_nl : STD_LOGIC;
  SIGNAL or_1484_nl : STD_LOGIC;
  SIGNAL nor_1112_nl : STD_LOGIC;
  SIGNAL mux_1636_nl : STD_LOGIC;
  SIGNAL mux_1635_nl : STD_LOGIC;
  SIGNAL mux_1634_nl : STD_LOGIC;
  SIGNAL nor_1113_nl : STD_LOGIC;
  SIGNAL mux_1633_nl : STD_LOGIC;
  SIGNAL or_1480_nl : STD_LOGIC;
  SIGNAL or_1478_nl : STD_LOGIC;
  SIGNAL nor_1114_nl : STD_LOGIC;
  SIGNAL mux_1632_nl : STD_LOGIC;
  SIGNAL mux_1631_nl : STD_LOGIC;
  SIGNAL or_1474_nl : STD_LOGIC;
  SIGNAL nor_1115_nl : STD_LOGIC;
  SIGNAL mux_1630_nl : STD_LOGIC;
  SIGNAL mux_1629_nl : STD_LOGIC;
  SIGNAL or_1467_nl : STD_LOGIC;
  SIGNAL or_1465_nl : STD_LOGIC;
  SIGNAL mux_1627_nl : STD_LOGIC;
  SIGNAL nor_1116_nl : STD_LOGIC;
  SIGNAL mux_1626_nl : STD_LOGIC;
  SIGNAL mux_1625_nl : STD_LOGIC;
  SIGNAL or_1460_nl : STD_LOGIC;
  SIGNAL or_1458_nl : STD_LOGIC;
  SIGNAL mux_1624_nl : STD_LOGIC;
  SIGNAL or_1457_nl : STD_LOGIC;
  SIGNAL or_1456_nl : STD_LOGIC;
  SIGNAL mux_1623_nl : STD_LOGIC;
  SIGNAL nor_1117_nl : STD_LOGIC;
  SIGNAL mux_1622_nl : STD_LOGIC;
  SIGNAL nor_1118_nl : STD_LOGIC;
  SIGNAL nor_1119_nl : STD_LOGIC;
  SIGNAL mux_1621_nl : STD_LOGIC;
  SIGNAL or_1451_nl : STD_LOGIC;
  SIGNAL or_1449_nl : STD_LOGIC;
  SIGNAL mux_1683_nl : STD_LOGIC;
  SIGNAL and_589_nl : STD_LOGIC;
  SIGNAL mux_1682_nl : STD_LOGIC;
  SIGNAL nor_1074_nl : STD_LOGIC;
  SIGNAL mux_1681_nl : STD_LOGIC;
  SIGNAL or_1558_nl : STD_LOGIC;
  SIGNAL or_1557_nl : STD_LOGIC;
  SIGNAL mux_1680_nl : STD_LOGIC;
  SIGNAL nor_1075_nl : STD_LOGIC;
  SIGNAL mux_1679_nl : STD_LOGIC;
  SIGNAL nor_1076_nl : STD_LOGIC;
  SIGNAL nor_1077_nl : STD_LOGIC;
  SIGNAL mux_1678_nl : STD_LOGIC;
  SIGNAL mux_1677_nl : STD_LOGIC;
  SIGNAL mux_1676_nl : STD_LOGIC;
  SIGNAL nor_1078_nl : STD_LOGIC;
  SIGNAL mux_1675_nl : STD_LOGIC;
  SIGNAL mux_1674_nl : STD_LOGIC;
  SIGNAL nor_1080_nl : STD_LOGIC;
  SIGNAL nor_1081_nl : STD_LOGIC;
  SIGNAL or_1544_nl : STD_LOGIC;
  SIGNAL mux_1673_nl : STD_LOGIC;
  SIGNAL nor_1082_nl : STD_LOGIC;
  SIGNAL mux_1672_nl : STD_LOGIC;
  SIGNAL nor_1083_nl : STD_LOGIC;
  SIGNAL nor_1084_nl : STD_LOGIC;
  SIGNAL mux_1671_nl : STD_LOGIC;
  SIGNAL mux_1670_nl : STD_LOGIC;
  SIGNAL nor_1085_nl : STD_LOGIC;
  SIGNAL nor_1086_nl : STD_LOGIC;
  SIGNAL nor_1087_nl : STD_LOGIC;
  SIGNAL mux_1668_nl : STD_LOGIC;
  SIGNAL mux_1667_nl : STD_LOGIC;
  SIGNAL mux_1666_nl : STD_LOGIC;
  SIGNAL mux_1665_nl : STD_LOGIC;
  SIGNAL and_590_nl : STD_LOGIC;
  SIGNAL mux_1664_nl : STD_LOGIC;
  SIGNAL nor_1088_nl : STD_LOGIC;
  SIGNAL nor_1089_nl : STD_LOGIC;
  SIGNAL and_591_nl : STD_LOGIC;
  SIGNAL mux_1663_nl : STD_LOGIC;
  SIGNAL nor_1090_nl : STD_LOGIC;
  SIGNAL nor_1091_nl : STD_LOGIC;
  SIGNAL mux_1662_nl : STD_LOGIC;
  SIGNAL nor_1092_nl : STD_LOGIC;
  SIGNAL nor_1093_nl : STD_LOGIC;
  SIGNAL mux_1660_nl : STD_LOGIC;
  SIGNAL nor_1094_nl : STD_LOGIC;
  SIGNAL mux_1659_nl : STD_LOGIC;
  SIGNAL nor_1095_nl : STD_LOGIC;
  SIGNAL nor_1096_nl : STD_LOGIC;
  SIGNAL mux_1658_nl : STD_LOGIC;
  SIGNAL mux_1657_nl : STD_LOGIC;
  SIGNAL nor_1097_nl : STD_LOGIC;
  SIGNAL nor_1098_nl : STD_LOGIC;
  SIGNAL mux_1656_nl : STD_LOGIC;
  SIGNAL mux_1655_nl : STD_LOGIC;
  SIGNAL mux_1654_nl : STD_LOGIC;
  SIGNAL nor_1099_nl : STD_LOGIC;
  SIGNAL mux_1653_nl : STD_LOGIC;
  SIGNAL nor_1100_nl : STD_LOGIC;
  SIGNAL nor_1101_nl : STD_LOGIC;
  SIGNAL nor_1102_nl : STD_LOGIC;
  SIGNAL mux_1652_nl : STD_LOGIC;
  SIGNAL nor_1103_nl : STD_LOGIC;
  SIGNAL nor_1104_nl : STD_LOGIC;
  SIGNAL mux_1714_nl : STD_LOGIC;
  SIGNAL mux_1713_nl : STD_LOGIC;
  SIGNAL mux_1712_nl : STD_LOGIC;
  SIGNAL nor_1059_nl : STD_LOGIC;
  SIGNAL mux_1711_nl : STD_LOGIC;
  SIGNAL mux_1710_nl : STD_LOGIC;
  SIGNAL or_1613_nl : STD_LOGIC;
  SIGNAL or_1612_nl : STD_LOGIC;
  SIGNAL or_1610_nl : STD_LOGIC;
  SIGNAL nor_1060_nl : STD_LOGIC;
  SIGNAL mux_1709_nl : STD_LOGIC;
  SIGNAL nor_1061_nl : STD_LOGIC;
  SIGNAL mux_1708_nl : STD_LOGIC;
  SIGNAL nor_1062_nl : STD_LOGIC;
  SIGNAL mux_1707_nl : STD_LOGIC;
  SIGNAL nor_1063_nl : STD_LOGIC;
  SIGNAL nor_1064_nl : STD_LOGIC;
  SIGNAL mux_1706_nl : STD_LOGIC;
  SIGNAL and_588_nl : STD_LOGIC;
  SIGNAL mux_1705_nl : STD_LOGIC;
  SIGNAL nand_287_nl : STD_LOGIC;
  SIGNAL mux_1704_nl : STD_LOGIC;
  SIGNAL or_1600_nl : STD_LOGIC;
  SIGNAL mux_1703_nl : STD_LOGIC;
  SIGNAL nor_1065_nl : STD_LOGIC;
  SIGNAL mux_1702_nl : STD_LOGIC;
  SIGNAL or_1597_nl : STD_LOGIC;
  SIGNAL mux_1701_nl : STD_LOGIC;
  SIGNAL or_1595_nl : STD_LOGIC;
  SIGNAL nor_1066_nl : STD_LOGIC;
  SIGNAL mux_1700_nl : STD_LOGIC;
  SIGNAL mux_1699_nl : STD_LOGIC;
  SIGNAL mux_1698_nl : STD_LOGIC;
  SIGNAL nor_1067_nl : STD_LOGIC;
  SIGNAL mux_1697_nl : STD_LOGIC;
  SIGNAL or_1591_nl : STD_LOGIC;
  SIGNAL or_1589_nl : STD_LOGIC;
  SIGNAL nor_1068_nl : STD_LOGIC;
  SIGNAL mux_1696_nl : STD_LOGIC;
  SIGNAL mux_1695_nl : STD_LOGIC;
  SIGNAL or_1585_nl : STD_LOGIC;
  SIGNAL nor_1069_nl : STD_LOGIC;
  SIGNAL mux_1694_nl : STD_LOGIC;
  SIGNAL mux_1693_nl : STD_LOGIC;
  SIGNAL or_1578_nl : STD_LOGIC;
  SIGNAL or_1576_nl : STD_LOGIC;
  SIGNAL mux_1691_nl : STD_LOGIC;
  SIGNAL nor_1070_nl : STD_LOGIC;
  SIGNAL mux_1690_nl : STD_LOGIC;
  SIGNAL mux_1689_nl : STD_LOGIC;
  SIGNAL or_1571_nl : STD_LOGIC;
  SIGNAL or_1569_nl : STD_LOGIC;
  SIGNAL mux_1688_nl : STD_LOGIC;
  SIGNAL or_1568_nl : STD_LOGIC;
  SIGNAL or_1567_nl : STD_LOGIC;
  SIGNAL mux_1687_nl : STD_LOGIC;
  SIGNAL nor_1071_nl : STD_LOGIC;
  SIGNAL mux_1686_nl : STD_LOGIC;
  SIGNAL nor_1072_nl : STD_LOGIC;
  SIGNAL nor_1073_nl : STD_LOGIC;
  SIGNAL mux_1685_nl : STD_LOGIC;
  SIGNAL or_1562_nl : STD_LOGIC;
  SIGNAL or_1560_nl : STD_LOGIC;
  SIGNAL mux_1747_nl : STD_LOGIC;
  SIGNAL and_585_nl : STD_LOGIC;
  SIGNAL mux_1746_nl : STD_LOGIC;
  SIGNAL nor_1028_nl : STD_LOGIC;
  SIGNAL mux_1745_nl : STD_LOGIC;
  SIGNAL or_1669_nl : STD_LOGIC;
  SIGNAL or_1668_nl : STD_LOGIC;
  SIGNAL mux_1744_nl : STD_LOGIC;
  SIGNAL nor_1029_nl : STD_LOGIC;
  SIGNAL mux_1743_nl : STD_LOGIC;
  SIGNAL nor_1030_nl : STD_LOGIC;
  SIGNAL nor_1031_nl : STD_LOGIC;
  SIGNAL mux_1742_nl : STD_LOGIC;
  SIGNAL mux_1741_nl : STD_LOGIC;
  SIGNAL mux_1740_nl : STD_LOGIC;
  SIGNAL nor_1032_nl : STD_LOGIC;
  SIGNAL mux_1739_nl : STD_LOGIC;
  SIGNAL mux_1738_nl : STD_LOGIC;
  SIGNAL nor_1034_nl : STD_LOGIC;
  SIGNAL nor_1035_nl : STD_LOGIC;
  SIGNAL or_1655_nl : STD_LOGIC;
  SIGNAL mux_1737_nl : STD_LOGIC;
  SIGNAL nor_1036_nl : STD_LOGIC;
  SIGNAL mux_1736_nl : STD_LOGIC;
  SIGNAL nor_1037_nl : STD_LOGIC;
  SIGNAL nor_1038_nl : STD_LOGIC;
  SIGNAL mux_1735_nl : STD_LOGIC;
  SIGNAL mux_1734_nl : STD_LOGIC;
  SIGNAL nor_1039_nl : STD_LOGIC;
  SIGNAL nor_1040_nl : STD_LOGIC;
  SIGNAL nor_1041_nl : STD_LOGIC;
  SIGNAL mux_1732_nl : STD_LOGIC;
  SIGNAL mux_1731_nl : STD_LOGIC;
  SIGNAL mux_1730_nl : STD_LOGIC;
  SIGNAL mux_1729_nl : STD_LOGIC;
  SIGNAL and_586_nl : STD_LOGIC;
  SIGNAL mux_1728_nl : STD_LOGIC;
  SIGNAL nor_1042_nl : STD_LOGIC;
  SIGNAL nor_1043_nl : STD_LOGIC;
  SIGNAL and_587_nl : STD_LOGIC;
  SIGNAL mux_1727_nl : STD_LOGIC;
  SIGNAL nor_1044_nl : STD_LOGIC;
  SIGNAL nor_1045_nl : STD_LOGIC;
  SIGNAL mux_1726_nl : STD_LOGIC;
  SIGNAL nor_1046_nl : STD_LOGIC;
  SIGNAL nor_1047_nl : STD_LOGIC;
  SIGNAL mux_1724_nl : STD_LOGIC;
  SIGNAL nor_1048_nl : STD_LOGIC;
  SIGNAL mux_1723_nl : STD_LOGIC;
  SIGNAL nor_1049_nl : STD_LOGIC;
  SIGNAL nor_1050_nl : STD_LOGIC;
  SIGNAL mux_1722_nl : STD_LOGIC;
  SIGNAL mux_1721_nl : STD_LOGIC;
  SIGNAL nor_1051_nl : STD_LOGIC;
  SIGNAL nor_1052_nl : STD_LOGIC;
  SIGNAL mux_1720_nl : STD_LOGIC;
  SIGNAL mux_1719_nl : STD_LOGIC;
  SIGNAL mux_1718_nl : STD_LOGIC;
  SIGNAL nor_1053_nl : STD_LOGIC;
  SIGNAL mux_1717_nl : STD_LOGIC;
  SIGNAL nor_1054_nl : STD_LOGIC;
  SIGNAL nor_1055_nl : STD_LOGIC;
  SIGNAL nor_1056_nl : STD_LOGIC;
  SIGNAL mux_1716_nl : STD_LOGIC;
  SIGNAL nor_1057_nl : STD_LOGIC;
  SIGNAL nor_1058_nl : STD_LOGIC;
  SIGNAL mux_1778_nl : STD_LOGIC;
  SIGNAL mux_1777_nl : STD_LOGIC;
  SIGNAL mux_1776_nl : STD_LOGIC;
  SIGNAL nor_1013_nl : STD_LOGIC;
  SIGNAL mux_1775_nl : STD_LOGIC;
  SIGNAL mux_1774_nl : STD_LOGIC;
  SIGNAL or_1723_nl : STD_LOGIC;
  SIGNAL or_1722_nl : STD_LOGIC;
  SIGNAL or_1720_nl : STD_LOGIC;
  SIGNAL nor_1014_nl : STD_LOGIC;
  SIGNAL mux_1773_nl : STD_LOGIC;
  SIGNAL nor_1015_nl : STD_LOGIC;
  SIGNAL mux_1772_nl : STD_LOGIC;
  SIGNAL nor_1016_nl : STD_LOGIC;
  SIGNAL mux_1771_nl : STD_LOGIC;
  SIGNAL nor_1017_nl : STD_LOGIC;
  SIGNAL nor_1018_nl : STD_LOGIC;
  SIGNAL mux_1770_nl : STD_LOGIC;
  SIGNAL and_584_nl : STD_LOGIC;
  SIGNAL mux_1769_nl : STD_LOGIC;
  SIGNAL nand_282_nl : STD_LOGIC;
  SIGNAL mux_1768_nl : STD_LOGIC;
  SIGNAL or_1710_nl : STD_LOGIC;
  SIGNAL mux_1767_nl : STD_LOGIC;
  SIGNAL nor_1019_nl : STD_LOGIC;
  SIGNAL mux_1766_nl : STD_LOGIC;
  SIGNAL or_1707_nl : STD_LOGIC;
  SIGNAL mux_1765_nl : STD_LOGIC;
  SIGNAL or_1705_nl : STD_LOGIC;
  SIGNAL nor_1020_nl : STD_LOGIC;
  SIGNAL mux_1764_nl : STD_LOGIC;
  SIGNAL mux_1763_nl : STD_LOGIC;
  SIGNAL mux_1762_nl : STD_LOGIC;
  SIGNAL nor_1021_nl : STD_LOGIC;
  SIGNAL mux_1761_nl : STD_LOGIC;
  SIGNAL or_1701_nl : STD_LOGIC;
  SIGNAL or_1699_nl : STD_LOGIC;
  SIGNAL nor_1022_nl : STD_LOGIC;
  SIGNAL mux_1760_nl : STD_LOGIC;
  SIGNAL mux_1759_nl : STD_LOGIC;
  SIGNAL or_1693_nl : STD_LOGIC;
  SIGNAL nor_1023_nl : STD_LOGIC;
  SIGNAL mux_1758_nl : STD_LOGIC;
  SIGNAL mux_1757_nl : STD_LOGIC;
  SIGNAL or_1689_nl : STD_LOGIC;
  SIGNAL or_1687_nl : STD_LOGIC;
  SIGNAL mux_1755_nl : STD_LOGIC;
  SIGNAL nor_1024_nl : STD_LOGIC;
  SIGNAL mux_1754_nl : STD_LOGIC;
  SIGNAL mux_1753_nl : STD_LOGIC;
  SIGNAL or_1682_nl : STD_LOGIC;
  SIGNAL or_1680_nl : STD_LOGIC;
  SIGNAL mux_1752_nl : STD_LOGIC;
  SIGNAL or_1679_nl : STD_LOGIC;
  SIGNAL or_1678_nl : STD_LOGIC;
  SIGNAL mux_1751_nl : STD_LOGIC;
  SIGNAL nor_1025_nl : STD_LOGIC;
  SIGNAL mux_1750_nl : STD_LOGIC;
  SIGNAL and_761_nl : STD_LOGIC;
  SIGNAL nor_1027_nl : STD_LOGIC;
  SIGNAL mux_1749_nl : STD_LOGIC;
  SIGNAL or_1673_nl : STD_LOGIC;
  SIGNAL or_1671_nl : STD_LOGIC;
  SIGNAL mux_1811_nl : STD_LOGIC;
  SIGNAL and_581_nl : STD_LOGIC;
  SIGNAL mux_1810_nl : STD_LOGIC;
  SIGNAL nor_982_nl : STD_LOGIC;
  SIGNAL mux_1809_nl : STD_LOGIC;
  SIGNAL or_1779_nl : STD_LOGIC;
  SIGNAL or_1778_nl : STD_LOGIC;
  SIGNAL mux_1808_nl : STD_LOGIC;
  SIGNAL nor_983_nl : STD_LOGIC;
  SIGNAL mux_1807_nl : STD_LOGIC;
  SIGNAL nor_984_nl : STD_LOGIC;
  SIGNAL nor_985_nl : STD_LOGIC;
  SIGNAL mux_1806_nl : STD_LOGIC;
  SIGNAL mux_1805_nl : STD_LOGIC;
  SIGNAL mux_1804_nl : STD_LOGIC;
  SIGNAL nor_986_nl : STD_LOGIC;
  SIGNAL mux_1803_nl : STD_LOGIC;
  SIGNAL mux_1802_nl : STD_LOGIC;
  SIGNAL nor_988_nl : STD_LOGIC;
  SIGNAL nor_989_nl : STD_LOGIC;
  SIGNAL or_1765_nl : STD_LOGIC;
  SIGNAL mux_1801_nl : STD_LOGIC;
  SIGNAL nor_990_nl : STD_LOGIC;
  SIGNAL mux_1800_nl : STD_LOGIC;
  SIGNAL nor_991_nl : STD_LOGIC;
  SIGNAL nor_992_nl : STD_LOGIC;
  SIGNAL mux_1799_nl : STD_LOGIC;
  SIGNAL mux_1798_nl : STD_LOGIC;
  SIGNAL nor_993_nl : STD_LOGIC;
  SIGNAL nor_994_nl : STD_LOGIC;
  SIGNAL nor_995_nl : STD_LOGIC;
  SIGNAL mux_1796_nl : STD_LOGIC;
  SIGNAL mux_1795_nl : STD_LOGIC;
  SIGNAL mux_1794_nl : STD_LOGIC;
  SIGNAL mux_1793_nl : STD_LOGIC;
  SIGNAL and_582_nl : STD_LOGIC;
  SIGNAL mux_1792_nl : STD_LOGIC;
  SIGNAL nor_996_nl : STD_LOGIC;
  SIGNAL nor_997_nl : STD_LOGIC;
  SIGNAL and_583_nl : STD_LOGIC;
  SIGNAL mux_1791_nl : STD_LOGIC;
  SIGNAL nor_998_nl : STD_LOGIC;
  SIGNAL nor_999_nl : STD_LOGIC;
  SIGNAL mux_1790_nl : STD_LOGIC;
  SIGNAL nor_1000_nl : STD_LOGIC;
  SIGNAL nor_1001_nl : STD_LOGIC;
  SIGNAL mux_1788_nl : STD_LOGIC;
  SIGNAL nor_1002_nl : STD_LOGIC;
  SIGNAL mux_1787_nl : STD_LOGIC;
  SIGNAL nor_1003_nl : STD_LOGIC;
  SIGNAL nor_1004_nl : STD_LOGIC;
  SIGNAL mux_1786_nl : STD_LOGIC;
  SIGNAL mux_1785_nl : STD_LOGIC;
  SIGNAL nor_1005_nl : STD_LOGIC;
  SIGNAL nor_1006_nl : STD_LOGIC;
  SIGNAL mux_1784_nl : STD_LOGIC;
  SIGNAL mux_1783_nl : STD_LOGIC;
  SIGNAL mux_1782_nl : STD_LOGIC;
  SIGNAL nor_1007_nl : STD_LOGIC;
  SIGNAL mux_1781_nl : STD_LOGIC;
  SIGNAL nor_1008_nl : STD_LOGIC;
  SIGNAL nor_1009_nl : STD_LOGIC;
  SIGNAL nor_1010_nl : STD_LOGIC;
  SIGNAL mux_1780_nl : STD_LOGIC;
  SIGNAL nor_1011_nl : STD_LOGIC;
  SIGNAL nor_1012_nl : STD_LOGIC;
  SIGNAL mux_1842_nl : STD_LOGIC;
  SIGNAL mux_1841_nl : STD_LOGIC;
  SIGNAL mux_1840_nl : STD_LOGIC;
  SIGNAL nor_967_nl : STD_LOGIC;
  SIGNAL mux_1839_nl : STD_LOGIC;
  SIGNAL mux_1838_nl : STD_LOGIC;
  SIGNAL nand_272_nl : STD_LOGIC;
  SIGNAL or_1832_nl : STD_LOGIC;
  SIGNAL or_1830_nl : STD_LOGIC;
  SIGNAL nor_968_nl : STD_LOGIC;
  SIGNAL mux_1837_nl : STD_LOGIC;
  SIGNAL nor_969_nl : STD_LOGIC;
  SIGNAL mux_1836_nl : STD_LOGIC;
  SIGNAL nor_970_nl : STD_LOGIC;
  SIGNAL mux_1835_nl : STD_LOGIC;
  SIGNAL nor_971_nl : STD_LOGIC;
  SIGNAL nor_972_nl : STD_LOGIC;
  SIGNAL mux_1834_nl : STD_LOGIC;
  SIGNAL and_580_nl : STD_LOGIC;
  SIGNAL mux_1833_nl : STD_LOGIC;
  SIGNAL nand_274_nl : STD_LOGIC;
  SIGNAL mux_1832_nl : STD_LOGIC;
  SIGNAL or_1820_nl : STD_LOGIC;
  SIGNAL mux_1831_nl : STD_LOGIC;
  SIGNAL nor_973_nl : STD_LOGIC;
  SIGNAL mux_1830_nl : STD_LOGIC;
  SIGNAL nand_398_nl : STD_LOGIC;
  SIGNAL mux_1829_nl : STD_LOGIC;
  SIGNAL or_1815_nl : STD_LOGIC;
  SIGNAL nor_974_nl : STD_LOGIC;
  SIGNAL mux_1828_nl : STD_LOGIC;
  SIGNAL mux_1827_nl : STD_LOGIC;
  SIGNAL mux_1826_nl : STD_LOGIC;
  SIGNAL nor_975_nl : STD_LOGIC;
  SIGNAL mux_1825_nl : STD_LOGIC;
  SIGNAL or_1811_nl : STD_LOGIC;
  SIGNAL or_1809_nl : STD_LOGIC;
  SIGNAL nor_976_nl : STD_LOGIC;
  SIGNAL mux_1824_nl : STD_LOGIC;
  SIGNAL mux_1823_nl : STD_LOGIC;
  SIGNAL or_1803_nl : STD_LOGIC;
  SIGNAL nor_977_nl : STD_LOGIC;
  SIGNAL mux_1822_nl : STD_LOGIC;
  SIGNAL mux_1821_nl : STD_LOGIC;
  SIGNAL or_1799_nl : STD_LOGIC;
  SIGNAL or_1797_nl : STD_LOGIC;
  SIGNAL mux_1819_nl : STD_LOGIC;
  SIGNAL nor_978_nl : STD_LOGIC;
  SIGNAL mux_1818_nl : STD_LOGIC;
  SIGNAL mux_1817_nl : STD_LOGIC;
  SIGNAL or_1792_nl : STD_LOGIC;
  SIGNAL or_1790_nl : STD_LOGIC;
  SIGNAL mux_1816_nl : STD_LOGIC;
  SIGNAL nand_277_nl : STD_LOGIC;
  SIGNAL or_1788_nl : STD_LOGIC;
  SIGNAL mux_1815_nl : STD_LOGIC;
  SIGNAL nor_979_nl : STD_LOGIC;
  SIGNAL mux_1814_nl : STD_LOGIC;
  SIGNAL nor_980_nl : STD_LOGIC;
  SIGNAL nor_981_nl : STD_LOGIC;
  SIGNAL mux_1813_nl : STD_LOGIC;
  SIGNAL or_1783_nl : STD_LOGIC;
  SIGNAL or_1781_nl : STD_LOGIC;
  SIGNAL mux_1875_nl : STD_LOGIC;
  SIGNAL and_575_nl : STD_LOGIC;
  SIGNAL mux_1874_nl : STD_LOGIC;
  SIGNAL nor_938_nl : STD_LOGIC;
  SIGNAL mux_1873_nl : STD_LOGIC;
  SIGNAL or_1889_nl : STD_LOGIC;
  SIGNAL or_1888_nl : STD_LOGIC;
  SIGNAL mux_1872_nl : STD_LOGIC;
  SIGNAL nor_939_nl : STD_LOGIC;
  SIGNAL mux_1871_nl : STD_LOGIC;
  SIGNAL nor_940_nl : STD_LOGIC;
  SIGNAL nor_941_nl : STD_LOGIC;
  SIGNAL mux_1870_nl : STD_LOGIC;
  SIGNAL mux_1869_nl : STD_LOGIC;
  SIGNAL mux_1868_nl : STD_LOGIC;
  SIGNAL nor_942_nl : STD_LOGIC;
  SIGNAL mux_1867_nl : STD_LOGIC;
  SIGNAL mux_1866_nl : STD_LOGIC;
  SIGNAL nor_944_nl : STD_LOGIC;
  SIGNAL nor_945_nl : STD_LOGIC;
  SIGNAL nand_265_nl : STD_LOGIC;
  SIGNAL mux_1865_nl : STD_LOGIC;
  SIGNAL nor_946_nl : STD_LOGIC;
  SIGNAL mux_1864_nl : STD_LOGIC;
  SIGNAL nor_947_nl : STD_LOGIC;
  SIGNAL nor_948_nl : STD_LOGIC;
  SIGNAL mux_1863_nl : STD_LOGIC;
  SIGNAL mux_1862_nl : STD_LOGIC;
  SIGNAL nor_949_nl : STD_LOGIC;
  SIGNAL nor_950_nl : STD_LOGIC;
  SIGNAL nor_951_nl : STD_LOGIC;
  SIGNAL mux_1860_nl : STD_LOGIC;
  SIGNAL mux_1859_nl : STD_LOGIC;
  SIGNAL mux_1858_nl : STD_LOGIC;
  SIGNAL mux_1857_nl : STD_LOGIC;
  SIGNAL and_576_nl : STD_LOGIC;
  SIGNAL mux_1856_nl : STD_LOGIC;
  SIGNAL nor_952_nl : STD_LOGIC;
  SIGNAL nor_953_nl : STD_LOGIC;
  SIGNAL and_577_nl : STD_LOGIC;
  SIGNAL mux_1855_nl : STD_LOGIC;
  SIGNAL nor_954_nl : STD_LOGIC;
  SIGNAL nor_955_nl : STD_LOGIC;
  SIGNAL mux_1854_nl : STD_LOGIC;
  SIGNAL nor_956_nl : STD_LOGIC;
  SIGNAL nor_957_nl : STD_LOGIC;
  SIGNAL mux_1852_nl : STD_LOGIC;
  SIGNAL nor_958_nl : STD_LOGIC;
  SIGNAL mux_1851_nl : STD_LOGIC;
  SIGNAL nor_959_nl : STD_LOGIC;
  SIGNAL and_578_nl : STD_LOGIC;
  SIGNAL mux_1850_nl : STD_LOGIC;
  SIGNAL mux_1849_nl : STD_LOGIC;
  SIGNAL nor_960_nl : STD_LOGIC;
  SIGNAL nor_961_nl : STD_LOGIC;
  SIGNAL mux_1848_nl : STD_LOGIC;
  SIGNAL mux_1847_nl : STD_LOGIC;
  SIGNAL mux_1846_nl : STD_LOGIC;
  SIGNAL nor_962_nl : STD_LOGIC;
  SIGNAL mux_1845_nl : STD_LOGIC;
  SIGNAL nor_963_nl : STD_LOGIC;
  SIGNAL nor_964_nl : STD_LOGIC;
  SIGNAL nor_965_nl : STD_LOGIC;
  SIGNAL mux_1844_nl : STD_LOGIC;
  SIGNAL and_579_nl : STD_LOGIC;
  SIGNAL nor_966_nl : STD_LOGIC;
  SIGNAL mux_1906_nl : STD_LOGIC;
  SIGNAL mux_1905_nl : STD_LOGIC;
  SIGNAL mux_1904_nl : STD_LOGIC;
  SIGNAL nor_923_nl : STD_LOGIC;
  SIGNAL mux_1903_nl : STD_LOGIC;
  SIGNAL mux_1902_nl : STD_LOGIC;
  SIGNAL or_1944_nl : STD_LOGIC;
  SIGNAL or_1943_nl : STD_LOGIC;
  SIGNAL or_1941_nl : STD_LOGIC;
  SIGNAL nor_924_nl : STD_LOGIC;
  SIGNAL mux_1901_nl : STD_LOGIC;
  SIGNAL nor_925_nl : STD_LOGIC;
  SIGNAL mux_1900_nl : STD_LOGIC;
  SIGNAL nor_926_nl : STD_LOGIC;
  SIGNAL mux_1899_nl : STD_LOGIC;
  SIGNAL nor_927_nl : STD_LOGIC;
  SIGNAL nor_928_nl : STD_LOGIC;
  SIGNAL mux_1898_nl : STD_LOGIC;
  SIGNAL and_574_nl : STD_LOGIC;
  SIGNAL mux_1897_nl : STD_LOGIC;
  SIGNAL nand_261_nl : STD_LOGIC;
  SIGNAL mux_1896_nl : STD_LOGIC;
  SIGNAL or_1931_nl : STD_LOGIC;
  SIGNAL mux_1895_nl : STD_LOGIC;
  SIGNAL nor_929_nl : STD_LOGIC;
  SIGNAL mux_1894_nl : STD_LOGIC;
  SIGNAL or_1928_nl : STD_LOGIC;
  SIGNAL mux_1893_nl : STD_LOGIC;
  SIGNAL or_1926_nl : STD_LOGIC;
  SIGNAL nor_930_nl : STD_LOGIC;
  SIGNAL mux_1892_nl : STD_LOGIC;
  SIGNAL mux_1891_nl : STD_LOGIC;
  SIGNAL mux_1890_nl : STD_LOGIC;
  SIGNAL nor_931_nl : STD_LOGIC;
  SIGNAL mux_1889_nl : STD_LOGIC;
  SIGNAL or_1922_nl : STD_LOGIC;
  SIGNAL or_1920_nl : STD_LOGIC;
  SIGNAL nor_932_nl : STD_LOGIC;
  SIGNAL mux_1888_nl : STD_LOGIC;
  SIGNAL mux_1887_nl : STD_LOGIC;
  SIGNAL or_1916_nl : STD_LOGIC;
  SIGNAL nor_933_nl : STD_LOGIC;
  SIGNAL mux_1886_nl : STD_LOGIC;
  SIGNAL mux_1885_nl : STD_LOGIC;
  SIGNAL or_1909_nl : STD_LOGIC;
  SIGNAL or_1907_nl : STD_LOGIC;
  SIGNAL mux_1883_nl : STD_LOGIC;
  SIGNAL nor_934_nl : STD_LOGIC;
  SIGNAL mux_1882_nl : STD_LOGIC;
  SIGNAL mux_1881_nl : STD_LOGIC;
  SIGNAL or_1902_nl : STD_LOGIC;
  SIGNAL or_1900_nl : STD_LOGIC;
  SIGNAL mux_1880_nl : STD_LOGIC;
  SIGNAL or_1899_nl : STD_LOGIC;
  SIGNAL or_1898_nl : STD_LOGIC;
  SIGNAL mux_1879_nl : STD_LOGIC;
  SIGNAL nor_935_nl : STD_LOGIC;
  SIGNAL mux_1878_nl : STD_LOGIC;
  SIGNAL nor_936_nl : STD_LOGIC;
  SIGNAL nor_937_nl : STD_LOGIC;
  SIGNAL mux_1877_nl : STD_LOGIC;
  SIGNAL or_1893_nl : STD_LOGIC;
  SIGNAL or_1891_nl : STD_LOGIC;
  SIGNAL mux_1939_nl : STD_LOGIC;
  SIGNAL and_571_nl : STD_LOGIC;
  SIGNAL mux_1938_nl : STD_LOGIC;
  SIGNAL nor_892_nl : STD_LOGIC;
  SIGNAL mux_1937_nl : STD_LOGIC;
  SIGNAL or_2000_nl : STD_LOGIC;
  SIGNAL or_1999_nl : STD_LOGIC;
  SIGNAL mux_1936_nl : STD_LOGIC;
  SIGNAL nor_893_nl : STD_LOGIC;
  SIGNAL mux_1935_nl : STD_LOGIC;
  SIGNAL nor_894_nl : STD_LOGIC;
  SIGNAL nor_895_nl : STD_LOGIC;
  SIGNAL mux_1934_nl : STD_LOGIC;
  SIGNAL mux_1933_nl : STD_LOGIC;
  SIGNAL mux_1932_nl : STD_LOGIC;
  SIGNAL nor_896_nl : STD_LOGIC;
  SIGNAL mux_1931_nl : STD_LOGIC;
  SIGNAL mux_1930_nl : STD_LOGIC;
  SIGNAL nor_898_nl : STD_LOGIC;
  SIGNAL nor_899_nl : STD_LOGIC;
  SIGNAL or_1986_nl : STD_LOGIC;
  SIGNAL mux_1929_nl : STD_LOGIC;
  SIGNAL nor_900_nl : STD_LOGIC;
  SIGNAL mux_1928_nl : STD_LOGIC;
  SIGNAL nor_901_nl : STD_LOGIC;
  SIGNAL nor_902_nl : STD_LOGIC;
  SIGNAL mux_1927_nl : STD_LOGIC;
  SIGNAL mux_1926_nl : STD_LOGIC;
  SIGNAL nor_903_nl : STD_LOGIC;
  SIGNAL nor_904_nl : STD_LOGIC;
  SIGNAL nor_905_nl : STD_LOGIC;
  SIGNAL mux_1924_nl : STD_LOGIC;
  SIGNAL mux_1923_nl : STD_LOGIC;
  SIGNAL mux_1922_nl : STD_LOGIC;
  SIGNAL mux_1921_nl : STD_LOGIC;
  SIGNAL and_572_nl : STD_LOGIC;
  SIGNAL mux_1920_nl : STD_LOGIC;
  SIGNAL nor_906_nl : STD_LOGIC;
  SIGNAL nor_907_nl : STD_LOGIC;
  SIGNAL and_573_nl : STD_LOGIC;
  SIGNAL mux_1919_nl : STD_LOGIC;
  SIGNAL nor_908_nl : STD_LOGIC;
  SIGNAL nor_909_nl : STD_LOGIC;
  SIGNAL mux_1918_nl : STD_LOGIC;
  SIGNAL nor_910_nl : STD_LOGIC;
  SIGNAL nor_911_nl : STD_LOGIC;
  SIGNAL mux_1916_nl : STD_LOGIC;
  SIGNAL nor_912_nl : STD_LOGIC;
  SIGNAL mux_1915_nl : STD_LOGIC;
  SIGNAL nor_913_nl : STD_LOGIC;
  SIGNAL nor_914_nl : STD_LOGIC;
  SIGNAL mux_1914_nl : STD_LOGIC;
  SIGNAL mux_1913_nl : STD_LOGIC;
  SIGNAL nor_915_nl : STD_LOGIC;
  SIGNAL nor_916_nl : STD_LOGIC;
  SIGNAL mux_1912_nl : STD_LOGIC;
  SIGNAL mux_1911_nl : STD_LOGIC;
  SIGNAL mux_1910_nl : STD_LOGIC;
  SIGNAL nor_917_nl : STD_LOGIC;
  SIGNAL mux_1909_nl : STD_LOGIC;
  SIGNAL nor_918_nl : STD_LOGIC;
  SIGNAL nor_919_nl : STD_LOGIC;
  SIGNAL nor_920_nl : STD_LOGIC;
  SIGNAL mux_1908_nl : STD_LOGIC;
  SIGNAL nor_921_nl : STD_LOGIC;
  SIGNAL nor_922_nl : STD_LOGIC;
  SIGNAL mux_1970_nl : STD_LOGIC;
  SIGNAL mux_1969_nl : STD_LOGIC;
  SIGNAL mux_1968_nl : STD_LOGIC;
  SIGNAL nor_877_nl : STD_LOGIC;
  SIGNAL mux_1967_nl : STD_LOGIC;
  SIGNAL mux_1966_nl : STD_LOGIC;
  SIGNAL nand_250_nl : STD_LOGIC;
  SIGNAL or_2054_nl : STD_LOGIC;
  SIGNAL or_2052_nl : STD_LOGIC;
  SIGNAL nor_878_nl : STD_LOGIC;
  SIGNAL mux_1965_nl : STD_LOGIC;
  SIGNAL nor_879_nl : STD_LOGIC;
  SIGNAL mux_1964_nl : STD_LOGIC;
  SIGNAL nor_880_nl : STD_LOGIC;
  SIGNAL mux_1963_nl : STD_LOGIC;
  SIGNAL nor_881_nl : STD_LOGIC;
  SIGNAL nor_882_nl : STD_LOGIC;
  SIGNAL mux_1962_nl : STD_LOGIC;
  SIGNAL and_570_nl : STD_LOGIC;
  SIGNAL mux_1961_nl : STD_LOGIC;
  SIGNAL nand_252_nl : STD_LOGIC;
  SIGNAL mux_1960_nl : STD_LOGIC;
  SIGNAL or_2042_nl : STD_LOGIC;
  SIGNAL mux_1959_nl : STD_LOGIC;
  SIGNAL nor_883_nl : STD_LOGIC;
  SIGNAL mux_1958_nl : STD_LOGIC;
  SIGNAL nand_397_nl : STD_LOGIC;
  SIGNAL mux_1957_nl : STD_LOGIC;
  SIGNAL or_2037_nl : STD_LOGIC;
  SIGNAL nor_884_nl : STD_LOGIC;
  SIGNAL mux_1956_nl : STD_LOGIC;
  SIGNAL mux_1955_nl : STD_LOGIC;
  SIGNAL mux_1954_nl : STD_LOGIC;
  SIGNAL nor_885_nl : STD_LOGIC;
  SIGNAL mux_1953_nl : STD_LOGIC;
  SIGNAL or_2033_nl : STD_LOGIC;
  SIGNAL or_2031_nl : STD_LOGIC;
  SIGNAL nor_886_nl : STD_LOGIC;
  SIGNAL mux_1952_nl : STD_LOGIC;
  SIGNAL mux_1951_nl : STD_LOGIC;
  SIGNAL or_2027_nl : STD_LOGIC;
  SIGNAL nor_887_nl : STD_LOGIC;
  SIGNAL mux_1950_nl : STD_LOGIC;
  SIGNAL mux_1949_nl : STD_LOGIC;
  SIGNAL or_2020_nl : STD_LOGIC;
  SIGNAL or_2018_nl : STD_LOGIC;
  SIGNAL mux_1947_nl : STD_LOGIC;
  SIGNAL nor_888_nl : STD_LOGIC;
  SIGNAL mux_1946_nl : STD_LOGIC;
  SIGNAL mux_1945_nl : STD_LOGIC;
  SIGNAL or_2013_nl : STD_LOGIC;
  SIGNAL or_2011_nl : STD_LOGIC;
  SIGNAL mux_1944_nl : STD_LOGIC;
  SIGNAL nand_255_nl : STD_LOGIC;
  SIGNAL or_2009_nl : STD_LOGIC;
  SIGNAL mux_1943_nl : STD_LOGIC;
  SIGNAL nor_889_nl : STD_LOGIC;
  SIGNAL mux_1942_nl : STD_LOGIC;
  SIGNAL nor_890_nl : STD_LOGIC;
  SIGNAL nor_891_nl : STD_LOGIC;
  SIGNAL mux_1941_nl : STD_LOGIC;
  SIGNAL or_2004_nl : STD_LOGIC;
  SIGNAL or_2002_nl : STD_LOGIC;
  SIGNAL mux_2003_nl : STD_LOGIC;
  SIGNAL and_565_nl : STD_LOGIC;
  SIGNAL mux_2002_nl : STD_LOGIC;
  SIGNAL nor_848_nl : STD_LOGIC;
  SIGNAL mux_2001_nl : STD_LOGIC;
  SIGNAL or_2111_nl : STD_LOGIC;
  SIGNAL or_2110_nl : STD_LOGIC;
  SIGNAL mux_2000_nl : STD_LOGIC;
  SIGNAL nor_849_nl : STD_LOGIC;
  SIGNAL mux_1999_nl : STD_LOGIC;
  SIGNAL nor_850_nl : STD_LOGIC;
  SIGNAL nor_851_nl : STD_LOGIC;
  SIGNAL mux_1998_nl : STD_LOGIC;
  SIGNAL mux_1997_nl : STD_LOGIC;
  SIGNAL mux_1996_nl : STD_LOGIC;
  SIGNAL nor_852_nl : STD_LOGIC;
  SIGNAL mux_1995_nl : STD_LOGIC;
  SIGNAL mux_1994_nl : STD_LOGIC;
  SIGNAL nor_854_nl : STD_LOGIC;
  SIGNAL nor_855_nl : STD_LOGIC;
  SIGNAL nand_243_nl : STD_LOGIC;
  SIGNAL mux_1993_nl : STD_LOGIC;
  SIGNAL nor_856_nl : STD_LOGIC;
  SIGNAL mux_1992_nl : STD_LOGIC;
  SIGNAL nor_857_nl : STD_LOGIC;
  SIGNAL nor_858_nl : STD_LOGIC;
  SIGNAL mux_1991_nl : STD_LOGIC;
  SIGNAL mux_1990_nl : STD_LOGIC;
  SIGNAL nor_859_nl : STD_LOGIC;
  SIGNAL nor_860_nl : STD_LOGIC;
  SIGNAL nor_861_nl : STD_LOGIC;
  SIGNAL mux_1988_nl : STD_LOGIC;
  SIGNAL mux_1987_nl : STD_LOGIC;
  SIGNAL mux_1986_nl : STD_LOGIC;
  SIGNAL mux_1985_nl : STD_LOGIC;
  SIGNAL and_566_nl : STD_LOGIC;
  SIGNAL mux_1984_nl : STD_LOGIC;
  SIGNAL nor_862_nl : STD_LOGIC;
  SIGNAL nor_863_nl : STD_LOGIC;
  SIGNAL and_567_nl : STD_LOGIC;
  SIGNAL mux_1983_nl : STD_LOGIC;
  SIGNAL nor_864_nl : STD_LOGIC;
  SIGNAL nor_865_nl : STD_LOGIC;
  SIGNAL mux_1982_nl : STD_LOGIC;
  SIGNAL nor_866_nl : STD_LOGIC;
  SIGNAL nor_867_nl : STD_LOGIC;
  SIGNAL mux_1980_nl : STD_LOGIC;
  SIGNAL nor_868_nl : STD_LOGIC;
  SIGNAL mux_1979_nl : STD_LOGIC;
  SIGNAL nor_869_nl : STD_LOGIC;
  SIGNAL and_568_nl : STD_LOGIC;
  SIGNAL mux_1978_nl : STD_LOGIC;
  SIGNAL mux_1977_nl : STD_LOGIC;
  SIGNAL nor_870_nl : STD_LOGIC;
  SIGNAL nor_871_nl : STD_LOGIC;
  SIGNAL mux_1976_nl : STD_LOGIC;
  SIGNAL mux_1975_nl : STD_LOGIC;
  SIGNAL mux_1974_nl : STD_LOGIC;
  SIGNAL nor_872_nl : STD_LOGIC;
  SIGNAL mux_1973_nl : STD_LOGIC;
  SIGNAL nor_873_nl : STD_LOGIC;
  SIGNAL nor_874_nl : STD_LOGIC;
  SIGNAL nor_875_nl : STD_LOGIC;
  SIGNAL mux_1972_nl : STD_LOGIC;
  SIGNAL and_569_nl : STD_LOGIC;
  SIGNAL nor_876_nl : STD_LOGIC;
  SIGNAL mux_2034_nl : STD_LOGIC;
  SIGNAL mux_2033_nl : STD_LOGIC;
  SIGNAL mux_2032_nl : STD_LOGIC;
  SIGNAL nor_833_nl : STD_LOGIC;
  SIGNAL mux_2031_nl : STD_LOGIC;
  SIGNAL mux_2030_nl : STD_LOGIC;
  SIGNAL nand_235_nl : STD_LOGIC;
  SIGNAL or_2164_nl : STD_LOGIC;
  SIGNAL or_2162_nl : STD_LOGIC;
  SIGNAL nor_834_nl : STD_LOGIC;
  SIGNAL mux_2029_nl : STD_LOGIC;
  SIGNAL nor_835_nl : STD_LOGIC;
  SIGNAL mux_2028_nl : STD_LOGIC;
  SIGNAL nor_836_nl : STD_LOGIC;
  SIGNAL mux_2027_nl : STD_LOGIC;
  SIGNAL nor_837_nl : STD_LOGIC;
  SIGNAL nor_838_nl : STD_LOGIC;
  SIGNAL mux_2026_nl : STD_LOGIC;
  SIGNAL and_563_nl : STD_LOGIC;
  SIGNAL mux_2025_nl : STD_LOGIC;
  SIGNAL nand_236_nl : STD_LOGIC;
  SIGNAL mux_2024_nl : STD_LOGIC;
  SIGNAL or_2152_nl : STD_LOGIC;
  SIGNAL mux_2023_nl : STD_LOGIC;
  SIGNAL nor_839_nl : STD_LOGIC;
  SIGNAL mux_2022_nl : STD_LOGIC;
  SIGNAL nand_396_nl : STD_LOGIC;
  SIGNAL mux_2021_nl : STD_LOGIC;
  SIGNAL or_2147_nl : STD_LOGIC;
  SIGNAL nor_840_nl : STD_LOGIC;
  SIGNAL mux_2020_nl : STD_LOGIC;
  SIGNAL mux_2019_nl : STD_LOGIC;
  SIGNAL mux_2018_nl : STD_LOGIC;
  SIGNAL nor_841_nl : STD_LOGIC;
  SIGNAL mux_2017_nl : STD_LOGIC;
  SIGNAL or_2143_nl : STD_LOGIC;
  SIGNAL or_2141_nl : STD_LOGIC;
  SIGNAL nor_842_nl : STD_LOGIC;
  SIGNAL mux_2016_nl : STD_LOGIC;
  SIGNAL mux_2015_nl : STD_LOGIC;
  SIGNAL or_2135_nl : STD_LOGIC;
  SIGNAL nor_843_nl : STD_LOGIC;
  SIGNAL mux_2014_nl : STD_LOGIC;
  SIGNAL mux_2013_nl : STD_LOGIC;
  SIGNAL or_2131_nl : STD_LOGIC;
  SIGNAL or_2129_nl : STD_LOGIC;
  SIGNAL mux_2011_nl : STD_LOGIC;
  SIGNAL nor_844_nl : STD_LOGIC;
  SIGNAL mux_2010_nl : STD_LOGIC;
  SIGNAL mux_2009_nl : STD_LOGIC;
  SIGNAL or_2124_nl : STD_LOGIC;
  SIGNAL or_2122_nl : STD_LOGIC;
  SIGNAL mux_2008_nl : STD_LOGIC;
  SIGNAL nand_239_nl : STD_LOGIC;
  SIGNAL or_2120_nl : STD_LOGIC;
  SIGNAL mux_2007_nl : STD_LOGIC;
  SIGNAL nor_845_nl : STD_LOGIC;
  SIGNAL mux_2006_nl : STD_LOGIC;
  SIGNAL nor_846_nl : STD_LOGIC;
  SIGNAL nor_847_nl : STD_LOGIC;
  SIGNAL mux_2005_nl : STD_LOGIC;
  SIGNAL or_2115_nl : STD_LOGIC;
  SIGNAL or_2113_nl : STD_LOGIC;
  SIGNAL mux_2067_nl : STD_LOGIC;
  SIGNAL and_558_nl : STD_LOGIC;
  SIGNAL mux_2066_nl : STD_LOGIC;
  SIGNAL nor_804_nl : STD_LOGIC;
  SIGNAL mux_2065_nl : STD_LOGIC;
  SIGNAL or_2221_nl : STD_LOGIC;
  SIGNAL or_2220_nl : STD_LOGIC;
  SIGNAL mux_2064_nl : STD_LOGIC;
  SIGNAL nor_805_nl : STD_LOGIC;
  SIGNAL mux_2063_nl : STD_LOGIC;
  SIGNAL nor_806_nl : STD_LOGIC;
  SIGNAL nor_807_nl : STD_LOGIC;
  SIGNAL mux_2062_nl : STD_LOGIC;
  SIGNAL mux_2061_nl : STD_LOGIC;
  SIGNAL mux_2060_nl : STD_LOGIC;
  SIGNAL nor_808_nl : STD_LOGIC;
  SIGNAL mux_2059_nl : STD_LOGIC;
  SIGNAL mux_2058_nl : STD_LOGIC;
  SIGNAL nor_810_nl : STD_LOGIC;
  SIGNAL nor_811_nl : STD_LOGIC;
  SIGNAL nand_228_nl : STD_LOGIC;
  SIGNAL mux_2057_nl : STD_LOGIC;
  SIGNAL nor_812_nl : STD_LOGIC;
  SIGNAL mux_2056_nl : STD_LOGIC;
  SIGNAL nor_813_nl : STD_LOGIC;
  SIGNAL nor_814_nl : STD_LOGIC;
  SIGNAL mux_2055_nl : STD_LOGIC;
  SIGNAL mux_2054_nl : STD_LOGIC;
  SIGNAL nor_815_nl : STD_LOGIC;
  SIGNAL nor_816_nl : STD_LOGIC;
  SIGNAL nor_817_nl : STD_LOGIC;
  SIGNAL mux_2052_nl : STD_LOGIC;
  SIGNAL mux_2051_nl : STD_LOGIC;
  SIGNAL mux_2050_nl : STD_LOGIC;
  SIGNAL mux_2049_nl : STD_LOGIC;
  SIGNAL and_559_nl : STD_LOGIC;
  SIGNAL mux_2048_nl : STD_LOGIC;
  SIGNAL nor_818_nl : STD_LOGIC;
  SIGNAL nor_819_nl : STD_LOGIC;
  SIGNAL and_560_nl : STD_LOGIC;
  SIGNAL mux_2047_nl : STD_LOGIC;
  SIGNAL nor_820_nl : STD_LOGIC;
  SIGNAL nor_821_nl : STD_LOGIC;
  SIGNAL mux_2046_nl : STD_LOGIC;
  SIGNAL nor_822_nl : STD_LOGIC;
  SIGNAL nor_823_nl : STD_LOGIC;
  SIGNAL mux_2044_nl : STD_LOGIC;
  SIGNAL nor_824_nl : STD_LOGIC;
  SIGNAL mux_2043_nl : STD_LOGIC;
  SIGNAL nor_825_nl : STD_LOGIC;
  SIGNAL and_561_nl : STD_LOGIC;
  SIGNAL mux_2042_nl : STD_LOGIC;
  SIGNAL mux_2041_nl : STD_LOGIC;
  SIGNAL nor_826_nl : STD_LOGIC;
  SIGNAL nor_827_nl : STD_LOGIC;
  SIGNAL mux_2040_nl : STD_LOGIC;
  SIGNAL mux_2039_nl : STD_LOGIC;
  SIGNAL mux_2038_nl : STD_LOGIC;
  SIGNAL nor_828_nl : STD_LOGIC;
  SIGNAL mux_2037_nl : STD_LOGIC;
  SIGNAL nor_829_nl : STD_LOGIC;
  SIGNAL nor_830_nl : STD_LOGIC;
  SIGNAL nor_831_nl : STD_LOGIC;
  SIGNAL mux_2036_nl : STD_LOGIC;
  SIGNAL and_562_nl : STD_LOGIC;
  SIGNAL nor_832_nl : STD_LOGIC;
  SIGNAL mux_2098_nl : STD_LOGIC;
  SIGNAL mux_2097_nl : STD_LOGIC;
  SIGNAL mux_2096_nl : STD_LOGIC;
  SIGNAL nor_789_nl : STD_LOGIC;
  SIGNAL mux_2095_nl : STD_LOGIC;
  SIGNAL mux_2094_nl : STD_LOGIC;
  SIGNAL and_554_nl : STD_LOGIC;
  SIGNAL or_2271_nl : STD_LOGIC;
  SIGNAL nor_790_nl : STD_LOGIC;
  SIGNAL mux_2093_nl : STD_LOGIC;
  SIGNAL nor_791_nl : STD_LOGIC;
  SIGNAL mux_2092_nl : STD_LOGIC;
  SIGNAL nor_792_nl : STD_LOGIC;
  SIGNAL mux_2091_nl : STD_LOGIC;
  SIGNAL nor_793_nl : STD_LOGIC;
  SIGNAL nor_794_nl : STD_LOGIC;
  SIGNAL mux_2090_nl : STD_LOGIC;
  SIGNAL and_555_nl : STD_LOGIC;
  SIGNAL mux_2089_nl : STD_LOGIC;
  SIGNAL nand_215_nl : STD_LOGIC;
  SIGNAL mux_2088_nl : STD_LOGIC;
  SIGNAL or_2261_nl : STD_LOGIC;
  SIGNAL mux_2087_nl : STD_LOGIC;
  SIGNAL nor_795_nl : STD_LOGIC;
  SIGNAL mux_2086_nl : STD_LOGIC;
  SIGNAL nand_395_nl : STD_LOGIC;
  SIGNAL mux_2085_nl : STD_LOGIC;
  SIGNAL or_2256_nl : STD_LOGIC;
  SIGNAL nor_796_nl : STD_LOGIC;
  SIGNAL mux_2084_nl : STD_LOGIC;
  SIGNAL mux_2083_nl : STD_LOGIC;
  SIGNAL mux_2082_nl : STD_LOGIC;
  SIGNAL nor_797_nl : STD_LOGIC;
  SIGNAL mux_2081_nl : STD_LOGIC;
  SIGNAL or_2253_nl : STD_LOGIC;
  SIGNAL or_2251_nl : STD_LOGIC;
  SIGNAL nor_798_nl : STD_LOGIC;
  SIGNAL mux_2080_nl : STD_LOGIC;
  SIGNAL mux_2079_nl : STD_LOGIC;
  SIGNAL or_2245_nl : STD_LOGIC;
  SIGNAL nor_799_nl : STD_LOGIC;
  SIGNAL mux_2078_nl : STD_LOGIC;
  SIGNAL mux_2077_nl : STD_LOGIC;
  SIGNAL or_2241_nl : STD_LOGIC;
  SIGNAL nand_219_nl : STD_LOGIC;
  SIGNAL mux_2075_nl : STD_LOGIC;
  SIGNAL nor_800_nl : STD_LOGIC;
  SIGNAL mux_2074_nl : STD_LOGIC;
  SIGNAL mux_2073_nl : STD_LOGIC;
  SIGNAL or_2234_nl : STD_LOGIC;
  SIGNAL or_2232_nl : STD_LOGIC;
  SIGNAL mux_2072_nl : STD_LOGIC;
  SIGNAL nand_220_nl : STD_LOGIC;
  SIGNAL nand_221_nl : STD_LOGIC;
  SIGNAL mux_2071_nl : STD_LOGIC;
  SIGNAL nor_801_nl : STD_LOGIC;
  SIGNAL mux_2070_nl : STD_LOGIC;
  SIGNAL nor_802_nl : STD_LOGIC;
  SIGNAL nor_803_nl : STD_LOGIC;
  SIGNAL mux_2069_nl : STD_LOGIC;
  SIGNAL or_2225_nl : STD_LOGIC;
  SIGNAL nand_223_nl : STD_LOGIC;
  SIGNAL mux_2131_nl : STD_LOGIC;
  SIGNAL and_546_nl : STD_LOGIC;
  SIGNAL mux_2130_nl : STD_LOGIC;
  SIGNAL nor_763_nl : STD_LOGIC;
  SIGNAL mux_2129_nl : STD_LOGIC;
  SIGNAL nand_199_nl : STD_LOGIC;
  SIGNAL or_2327_nl : STD_LOGIC;
  SIGNAL mux_2128_nl : STD_LOGIC;
  SIGNAL nor_764_nl : STD_LOGIC;
  SIGNAL mux_2127_nl : STD_LOGIC;
  SIGNAL nor_765_nl : STD_LOGIC;
  SIGNAL nor_766_nl : STD_LOGIC;
  SIGNAL mux_2126_nl : STD_LOGIC;
  SIGNAL mux_2125_nl : STD_LOGIC;
  SIGNAL mux_2124_nl : STD_LOGIC;
  SIGNAL nor_767_nl : STD_LOGIC;
  SIGNAL mux_2123_nl : STD_LOGIC;
  SIGNAL mux_2122_nl : STD_LOGIC;
  SIGNAL nor_769_nl : STD_LOGIC;
  SIGNAL nor_770_nl : STD_LOGIC;
  SIGNAL nand_203_nl : STD_LOGIC;
  SIGNAL mux_2121_nl : STD_LOGIC;
  SIGNAL nor_771_nl : STD_LOGIC;
  SIGNAL mux_2120_nl : STD_LOGIC;
  SIGNAL and_547_nl : STD_LOGIC;
  SIGNAL nor_772_nl : STD_LOGIC;
  SIGNAL mux_2119_nl : STD_LOGIC;
  SIGNAL mux_2118_nl : STD_LOGIC;
  SIGNAL nor_773_nl : STD_LOGIC;
  SIGNAL nor_774_nl : STD_LOGIC;
  SIGNAL nor_775_nl : STD_LOGIC;
  SIGNAL mux_2116_nl : STD_LOGIC;
  SIGNAL mux_2115_nl : STD_LOGIC;
  SIGNAL mux_2114_nl : STD_LOGIC;
  SIGNAL mux_2113_nl : STD_LOGIC;
  SIGNAL and_548_nl : STD_LOGIC;
  SIGNAL mux_2112_nl : STD_LOGIC;
  SIGNAL nor_776_nl : STD_LOGIC;
  SIGNAL nor_777_nl : STD_LOGIC;
  SIGNAL and_549_nl : STD_LOGIC;
  SIGNAL mux_2111_nl : STD_LOGIC;
  SIGNAL nor_778_nl : STD_LOGIC;
  SIGNAL and_759_nl : STD_LOGIC;
  SIGNAL mux_2110_nl : STD_LOGIC;
  SIGNAL nor_780_nl : STD_LOGIC;
  SIGNAL nor_781_nl : STD_LOGIC;
  SIGNAL mux_2108_nl : STD_LOGIC;
  SIGNAL nor_782_nl : STD_LOGIC;
  SIGNAL mux_2107_nl : STD_LOGIC;
  SIGNAL and_550_nl : STD_LOGIC;
  SIGNAL and_551_nl : STD_LOGIC;
  SIGNAL mux_2106_nl : STD_LOGIC;
  SIGNAL mux_2105_nl : STD_LOGIC;
  SIGNAL nor_783_nl : STD_LOGIC;
  SIGNAL nor_784_nl : STD_LOGIC;
  SIGNAL mux_2104_nl : STD_LOGIC;
  SIGNAL mux_2103_nl : STD_LOGIC;
  SIGNAL mux_2102_nl : STD_LOGIC;
  SIGNAL nor_785_nl : STD_LOGIC;
  SIGNAL mux_2101_nl : STD_LOGIC;
  SIGNAL nor_786_nl : STD_LOGIC;
  SIGNAL nor_787_nl : STD_LOGIC;
  SIGNAL and_552_nl : STD_LOGIC;
  SIGNAL mux_2100_nl : STD_LOGIC;
  SIGNAL and_553_nl : STD_LOGIC;
  SIGNAL nor_788_nl : STD_LOGIC;
  SIGNAL mux_3811_nl : STD_LOGIC;
  SIGNAL nor_1648_nl : STD_LOGIC;
  SIGNAL mux_3810_nl : STD_LOGIC;
  SIGNAL mux_3809_nl : STD_LOGIC;
  SIGNAL or_3467_nl : STD_LOGIC;
  SIGNAL or_3466_nl : STD_LOGIC;
  SIGNAL or_3465_nl : STD_LOGIC;
  SIGNAL mux_3808_nl : STD_LOGIC;
  SIGNAL nor_1649_nl : STD_LOGIC;
  SIGNAL mux_3807_nl : STD_LOGIC;
  SIGNAL mux_3806_nl : STD_LOGIC;
  SIGNAL mux_3805_nl : STD_LOGIC;
  SIGNAL nor_1650_nl : STD_LOGIC;
  SIGNAL nor_1651_nl : STD_LOGIC;
  SIGNAL nor_1652_nl : STD_LOGIC;
  SIGNAL and_nl : STD_LOGIC;
  SIGNAL mux_3804_nl : STD_LOGIC;
  SIGNAL or_3456_nl : STD_LOGIC;
  SIGNAL mux_3803_nl : STD_LOGIC;
  SIGNAL mux_3802_nl : STD_LOGIC;
  SIGNAL and_1158_nl : STD_LOGIC;
  SIGNAL mux_3801_nl : STD_LOGIC;
  SIGNAL nor_1653_nl : STD_LOGIC;
  SIGNAL nor_1654_nl : STD_LOGIC;
  SIGNAL mux_3800_nl : STD_LOGIC;
  SIGNAL nor_1655_nl : STD_LOGIC;
  SIGNAL nor_1656_nl : STD_LOGIC;
  SIGNAL mux_3828_nl : STD_LOGIC;
  SIGNAL or_3448_nl : STD_LOGIC;
  SIGNAL mux_3821_nl : STD_LOGIC;
  SIGNAL mux_3829_nl : STD_LOGIC;
  SIGNAL or_3510_nl : STD_LOGIC;
  SIGNAL mux_3842_nl : STD_LOGIC;
  SIGNAL or_3520_nl : STD_LOGIC;
  SIGNAL or_3527_nl : STD_LOGIC;
  SIGNAL mux_3849_nl : STD_LOGIC;
  SIGNAL mux_3893_nl : STD_LOGIC;
  SIGNAL or_3564_nl : STD_LOGIC;
  SIGNAL mux_3904_nl : STD_LOGIC;
  SIGNAL or_3586_nl : STD_LOGIC;
  SIGNAL or_3585_nl : STD_LOGIC;
  SIGNAL mux_3907_nl : STD_LOGIC;
  SIGNAL or_3584_nl : STD_LOGIC;
  SIGNAL or_3583_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_mux_2_nl : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL operator_64_false_1_mux_3_nl : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_COMP_LOOP_or_72_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_73_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_575_nl : STD_LOGIC_VECTOR (62 DOWNTO 0);
  SIGNAL COMP_LOOP_COMP_LOOP_and_938_nl : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL COMP_LOOP_nor_695_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_acc_105_nl : STD_LOGIC_VECTOR (12 DOWNTO 0);
  SIGNAL COMP_LOOP_mux1h_576_nl : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL COMP_LOOP_mux1h_577_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL COMP_LOOP_or_69_nl : STD_LOGIC;
  SIGNAL acc_3_nl : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL COMP_LOOP_COMP_LOOP_or_74_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_mux_18_nl : STD_LOGIC_VECTOR (8 DOWNTO 0);
  SIGNAL COMP_LOOP_or_70_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_mux_19_nl : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL COMP_LOOP_COMP_LOOP_or_75_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_76_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_77_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_78_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux_82_nl : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_COMP_LOOP_mux_20_nl : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL COMP_LOOP_COMP_LOOP_or_79_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_80_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_81_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_82_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_71_nl : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL COMP_LOOP_mux1h_578_nl : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL and_1178_nl : STD_LOGIC;
  SIGNAL and_1179_nl : STD_LOGIC;
  SIGNAL and_1180_nl : STD_LOGIC;
  SIGNAL and_1181_nl : STD_LOGIC;
  SIGNAL and_1182_nl : STD_LOGIC;
  SIGNAL and_1183_nl : STD_LOGIC;
  SIGNAL and_1184_nl : STD_LOGIC;
  SIGNAL and_1185_nl : STD_LOGIC;
  SIGNAL acc_6_nl : STD_LOGIC_VECTOR (65 DOWNTO 0);
  SIGNAL COMP_LOOP_COMP_LOOP_or_83_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_84_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_85_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_86_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_87_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_88_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_89_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_90_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_91_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_92_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_93_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_94_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_95_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_96_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_97_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_98_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_99_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_100_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_101_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_102_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_103_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_104_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_105_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_106_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_107_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_108_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_109_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_110_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_111_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_112_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_113_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_114_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_115_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_116_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_117_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_118_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_119_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_120_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_121_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_122_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_123_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_124_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_125_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_126_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_127_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_128_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_129_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_130_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_131_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_132_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_133_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_134_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_135_nl : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL COMP_LOOP_and_398_nl : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL COMP_LOOP_mux_83_nl : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL COMP_LOOP_or_72_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_73_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_579_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_580_nl : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL COMP_LOOP_or_74_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_136_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_137_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_138_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_75_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL COMP_LOOP_and_401_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL COMP_LOOP_COMP_LOOP_mux_21_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL COMP_LOOP_nor_706_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_139_nl : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL COMP_LOOP_and_402_nl : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL COMP_LOOP_nor_707_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_140_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_141_nl : STD_LOGIC;
  SIGNAL acc_7_nl : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL COMP_LOOP_COMP_LOOP_or_142_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_581_nl : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL COMP_LOOP_or_76_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_mux_22_nl : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL COMP_LOOP_or_77_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_143_nl : STD_LOGIC;
  SIGNAL modExp_while_if_mux_1_nl : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mux_3947_nl : STD_LOGIC;
  SIGNAL mux_3948_nl : STD_LOGIC;
  SIGNAL nor_1711_nl : STD_LOGIC;
  SIGNAL mux_3949_nl : STD_LOGIC;
  SIGNAL or_3639_nl : STD_LOGIC;
  SIGNAL mux_3950_nl : STD_LOGIC;
  SIGNAL or_3640_nl : STD_LOGIC;
  SIGNAL mux_3951_nl : STD_LOGIC;
  SIGNAL and_1186_nl : STD_LOGIC;
  SIGNAL mux_3952_nl : STD_LOGIC;
  SIGNAL mux_3953_nl : STD_LOGIC;
  SIGNAL nor_1712_nl : STD_LOGIC;
  SIGNAL mux_3954_nl : STD_LOGIC;
  SIGNAL or_3641_nl : STD_LOGIC;
  SIGNAL or_3642_nl : STD_LOGIC;
  SIGNAL nor_1713_nl : STD_LOGIC;
  SIGNAL mux_3955_nl : STD_LOGIC;
  SIGNAL nand_428_nl : STD_LOGIC;
  SIGNAL or_3643_nl : STD_LOGIC;
  SIGNAL mux_3956_nl : STD_LOGIC;
  SIGNAL mux_3957_nl : STD_LOGIC;
  SIGNAL and_1187_nl : STD_LOGIC;
  SIGNAL mux_3958_nl : STD_LOGIC;
  SIGNAL and_1188_nl : STD_LOGIC;
  SIGNAL mux_3959_nl : STD_LOGIC;
  SIGNAL or_3644_nl : STD_LOGIC;
  SIGNAL nor_1714_nl : STD_LOGIC;
  SIGNAL mux_3960_nl : STD_LOGIC;
  SIGNAL or_3645_nl : STD_LOGIC;
  SIGNAL p_rsci_dat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL p_rsci_idat_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL r_rsci_dat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL r_rsci_idat_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL modulo_result_rem_cmp_a_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL modulo_result_rem_cmp_b_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL modulo_result_rem_cmp_z_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL operator_66_true_div_cmp_a_1 : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL operator_66_true_div_cmp_b : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL operator_66_true_div_cmp_z_1 : STD_LOGIC_VECTOR (64 DOWNTO 0);

  SIGNAL STAGE_LOOP_lshift_rg_a : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL STAGE_LOOP_lshift_rg_s : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL STAGE_LOOP_lshift_rg_z : STD_LOGIC_VECTOR (9 DOWNTO 0);

  COMPONENT inPlaceNTT_DIT_core_core_fsm
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      fsm_output : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
      STAGE_LOOP_C_8_tr0 : IN STD_LOGIC;
      modExp_while_C_38_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_1_tr0 : IN STD_LOGIC;
      COMP_LOOP_1_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_64_tr0 : IN STD_LOGIC;
      COMP_LOOP_2_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_128_tr0 : IN STD_LOGIC;
      COMP_LOOP_3_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_192_tr0 : IN STD_LOGIC;
      COMP_LOOP_4_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_256_tr0 : IN STD_LOGIC;
      COMP_LOOP_5_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_320_tr0 : IN STD_LOGIC;
      COMP_LOOP_6_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_384_tr0 : IN STD_LOGIC;
      COMP_LOOP_7_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_448_tr0 : IN STD_LOGIC;
      COMP_LOOP_8_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_512_tr0 : IN STD_LOGIC;
      COMP_LOOP_9_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_576_tr0 : IN STD_LOGIC;
      COMP_LOOP_10_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_640_tr0 : IN STD_LOGIC;
      COMP_LOOP_11_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_704_tr0 : IN STD_LOGIC;
      COMP_LOOP_12_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_768_tr0 : IN STD_LOGIC;
      COMP_LOOP_13_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_832_tr0 : IN STD_LOGIC;
      COMP_LOOP_14_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_896_tr0 : IN STD_LOGIC;
      COMP_LOOP_15_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_960_tr0 : IN STD_LOGIC;
      COMP_LOOP_16_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_1024_tr0 : IN STD_LOGIC;
      VEC_LOOP_C_0_tr0 : IN STD_LOGIC;
      STAGE_LOOP_C_9_tr0 : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_fsm_output : STD_LOGIC_VECTOR (10 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_8_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_1_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_64_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_2_modExp_1_while_C_38_tr0 :
      STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_128_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_3_modExp_1_while_C_38_tr0 :
      STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_192_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_4_modExp_1_while_C_38_tr0 :
      STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_256_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_5_modExp_1_while_C_38_tr0 :
      STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_320_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_6_modExp_1_while_C_38_tr0 :
      STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_384_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_7_modExp_1_while_C_38_tr0 :
      STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_448_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_8_modExp_1_while_C_38_tr0 :
      STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_512_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_9_modExp_1_while_C_38_tr0 :
      STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_576_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_10_modExp_1_while_C_38_tr0 :
      STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_640_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_11_modExp_1_while_C_38_tr0 :
      STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_704_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_12_modExp_1_while_C_38_tr0 :
      STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_768_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_13_modExp_1_while_C_38_tr0 :
      STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_832_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_14_modExp_1_while_C_38_tr0 :
      STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_896_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_15_modExp_1_while_C_38_tr0 :
      STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_960_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_16_modExp_1_while_C_38_tr0 :
      STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_C_0_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_9_tr0 : STD_LOGIC;

  FUNCTION CONV_SL_1_1(input_val:BOOLEAN)
  RETURN STD_LOGIC IS
  BEGIN
    IF input_val THEN RETURN '1';ELSE RETURN '0';END IF;
  END;

  FUNCTION MUX1HOT_s_1_3_2(input_2 : STD_LOGIC;
  input_1 : STD_LOGIC;
  input_0 : STD_LOGIC;
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;
    VARIABLE tmp : STD_LOGIC;

    BEGIN
      tmp := sel(0);
      result := input_0 and tmp;
      tmp := sel(1);
      result := result or ( input_1 and tmp);
      tmp := sel(2);
      result := result or ( input_2 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_s_1_4_2(input_3 : STD_LOGIC;
  input_2 : STD_LOGIC;
  input_1 : STD_LOGIC;
  input_0 : STD_LOGIC;
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;
    VARIABLE tmp : STD_LOGIC;

    BEGIN
      tmp := sel(0);
      result := input_0 and tmp;
      tmp := sel(1);
      result := result or ( input_1 and tmp);
      tmp := sel(2);
      result := result or ( input_2 and tmp);
      tmp := sel(3);
      result := result or ( input_3 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_s_1_6_2(input_5 : STD_LOGIC;
  input_4 : STD_LOGIC;
  input_3 : STD_LOGIC;
  input_2 : STD_LOGIC;
  input_1 : STD_LOGIC;
  input_0 : STD_LOGIC;
  sel : STD_LOGIC_VECTOR(5 DOWNTO 0))
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;
    VARIABLE tmp : STD_LOGIC;

    BEGIN
      tmp := sel(0);
      result := input_0 and tmp;
      tmp := sel(1);
      result := result or ( input_1 and tmp);
      tmp := sel(2);
      result := result or ( input_2 and tmp);
      tmp := sel(3);
      result := result or ( input_3 and tmp);
      tmp := sel(4);
      result := result or ( input_4 and tmp);
      tmp := sel(5);
      result := result or ( input_5 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_3_3_2(input_2 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(2 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(2 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_4_7_2(input_6 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(6 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(3 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(3 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_63_4_2(input_3 : STD_LOGIC_VECTOR(62 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(62 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(62 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(62 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(62 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(62 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_64_17_2(input_16 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_15 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_14 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_13 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_12 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_11 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_10 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(16 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(63 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(63 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
      tmp := (OTHERS=>sel( 9));
      result := result or ( input_9 and tmp);
      tmp := (OTHERS=>sel( 10));
      result := result or ( input_10 and tmp);
      tmp := (OTHERS=>sel( 11));
      result := result or ( input_11 and tmp);
      tmp := (OTHERS=>sel( 12));
      result := result or ( input_12 and tmp);
      tmp := (OTHERS=>sel( 13));
      result := result or ( input_13 and tmp);
      tmp := (OTHERS=>sel( 14));
      result := result or ( input_14 and tmp);
      tmp := (OTHERS=>sel( 15));
      result := result or ( input_15 and tmp);
      tmp := (OTHERS=>sel( 16));
      result := result or ( input_16 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_64_21_2(input_20 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_19 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_18 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_17 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_16 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_15 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_14 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_13 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_12 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_11 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_10 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(20 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(63 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(63 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
      tmp := (OTHERS=>sel( 9));
      result := result or ( input_9 and tmp);
      tmp := (OTHERS=>sel( 10));
      result := result or ( input_10 and tmp);
      tmp := (OTHERS=>sel( 11));
      result := result or ( input_11 and tmp);
      tmp := (OTHERS=>sel( 12));
      result := result or ( input_12 and tmp);
      tmp := (OTHERS=>sel( 13));
      result := result or ( input_13 and tmp);
      tmp := (OTHERS=>sel( 14));
      result := result or ( input_14 and tmp);
      tmp := (OTHERS=>sel( 15));
      result := result or ( input_15 and tmp);
      tmp := (OTHERS=>sel( 16));
      result := result or ( input_16 and tmp);
      tmp := (OTHERS=>sel( 17));
      result := result or ( input_17 and tmp);
      tmp := (OTHERS=>sel( 18));
      result := result or ( input_18 and tmp);
      tmp := (OTHERS=>sel( 19));
      result := result or ( input_19 and tmp);
      tmp := (OTHERS=>sel( 20));
      result := result or ( input_20 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_64_3_2(input_2 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(63 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(63 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_64_6_2(input_5 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(5 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(63 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(63 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_65_3_2(input_2 : STD_LOGIC_VECTOR(64 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(64 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(64 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(64 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(64 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_6_4_2(input_3 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(5 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(5 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_7_4_2(input_3 : STD_LOGIC_VECTOR(6 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(6 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(6 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(6 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(6 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(6 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_7_5_2(input_4 : STD_LOGIC_VECTOR(6 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(6 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(6 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(6 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(6 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(4 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(6 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(6 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_8_19_2(input_18 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_17 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_16 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_15 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_14 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_13 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_12 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_11 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_10 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(18 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(7 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(7 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
      tmp := (OTHERS=>sel( 9));
      result := result or ( input_9 and tmp);
      tmp := (OTHERS=>sel( 10));
      result := result or ( input_10 and tmp);
      tmp := (OTHERS=>sel( 11));
      result := result or ( input_11 and tmp);
      tmp := (OTHERS=>sel( 12));
      result := result or ( input_12 and tmp);
      tmp := (OTHERS=>sel( 13));
      result := result or ( input_13 and tmp);
      tmp := (OTHERS=>sel( 14));
      result := result or ( input_14 and tmp);
      tmp := (OTHERS=>sel( 15));
      result := result or ( input_15 and tmp);
      tmp := (OTHERS=>sel( 16));
      result := result or ( input_16 and tmp);
      tmp := (OTHERS=>sel( 17));
      result := result or ( input_17 and tmp);
      tmp := (OTHERS=>sel( 18));
      result := result or ( input_18 and tmp);
    RETURN result;
  END;

  FUNCTION MUX_s_1_2_2(input_0 : STD_LOGIC;
  input_1 : STD_LOGIC;
  sel : STD_LOGIC)
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_10_2_2(input_0 : STD_LOGIC_VECTOR(9 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(9 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(9 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_12_2_2(input_0 : STD_LOGIC_VECTOR(11 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(11 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(11 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_2_2_2(input_0 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(1 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_3_2_2(input_0 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(2 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_4_2_2(input_0 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(3 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_63_2_2(input_0 : STD_LOGIC_VECTOR(62 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(62 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(62 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_64_2_2(input_0 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(63 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_65_2_2(input_0 : STD_LOGIC_VECTOR(64 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(64 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(64 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_9_2_2(input_0 : STD_LOGIC_VECTOR(8 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(8 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(8 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  p_rsci : work.ccs_in_pkg_v1.ccs_in_v1
    GENERIC MAP(
      rscid => 2,
      width => 64
      )
    PORT MAP(
      dat => p_rsci_dat,
      idat => p_rsci_idat_1
    );
  p_rsci_dat <= p_rsc_dat;
  p_rsci_idat <= p_rsci_idat_1;

  r_rsci : work.ccs_in_pkg_v1.ccs_in_v1
    GENERIC MAP(
      rscid => 3,
      width => 64
      )
    PORT MAP(
      dat => r_rsci_dat,
      idat => r_rsci_idat_1
    );
  r_rsci_dat <= r_rsc_dat;
  r_rsci_idat <= r_rsci_idat_1;

  vec_rsc_triosy_0_15_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_15_lz
    );
  vec_rsc_triosy_0_14_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_14_lz
    );
  vec_rsc_triosy_0_13_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_13_lz
    );
  vec_rsc_triosy_0_12_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_12_lz
    );
  vec_rsc_triosy_0_11_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_11_lz
    );
  vec_rsc_triosy_0_10_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_10_lz
    );
  vec_rsc_triosy_0_9_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_9_lz
    );
  vec_rsc_triosy_0_8_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_8_lz
    );
  vec_rsc_triosy_0_7_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_7_lz
    );
  vec_rsc_triosy_0_6_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_6_lz
    );
  vec_rsc_triosy_0_5_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_5_lz
    );
  vec_rsc_triosy_0_4_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_4_lz
    );
  vec_rsc_triosy_0_3_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_3_lz
    );
  vec_rsc_triosy_0_2_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_2_lz
    );
  vec_rsc_triosy_0_1_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_1_lz
    );
  vec_rsc_triosy_0_0_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_0_lz
    );
  p_rsc_triosy_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => p_rsc_triosy_lz
    );
  r_rsc_triosy_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => r_rsc_triosy_lz
    );
  modulo_result_rem_cmp : work.mgc_comps.mgc_rem
    GENERIC MAP(
      width_a => 64,
      width_b => 64,
      signd => 1
      )
    PORT MAP(
      a => modulo_result_rem_cmp_a_1,
      b => modulo_result_rem_cmp_b_1,
      z => modulo_result_rem_cmp_z_1
    );
  modulo_result_rem_cmp_a_1 <= modulo_result_rem_cmp_a;
  modulo_result_rem_cmp_b_1 <= modulo_result_rem_cmp_b;
  modulo_result_rem_cmp_z <= modulo_result_rem_cmp_z_1;

  operator_66_true_div_cmp : work.mgc_comps.mgc_div
    GENERIC MAP(
      width_a => 65,
      width_b => 11,
      signd => 1
      )
    PORT MAP(
      a => operator_66_true_div_cmp_a_1,
      b => operator_66_true_div_cmp_b,
      z => operator_66_true_div_cmp_z_1
    );
  operator_66_true_div_cmp_a_1 <= operator_66_true_div_cmp_a;
  operator_66_true_div_cmp_b <= STD_LOGIC_VECTOR(UNSIGNED'( "0") & UNSIGNED(operator_66_true_div_cmp_b_9_0));
  operator_66_true_div_cmp_z <= operator_66_true_div_cmp_z_1;

  STAGE_LOOP_lshift_rg : work.mgc_shift_comps_v5.mgc_shift_l_v5
    GENERIC MAP(
      width_a => 1,
      signd_a => 0,
      width_s => 4,
      width_z => 10
      )
    PORT MAP(
      a => STAGE_LOOP_lshift_rg_a,
      s => STAGE_LOOP_lshift_rg_s,
      z => STAGE_LOOP_lshift_rg_z
    );
  STAGE_LOOP_lshift_rg_a(0) <= '1';
  STAGE_LOOP_lshift_rg_s <= STAGE_LOOP_i_3_0_sva;
  STAGE_LOOP_lshift_psp_sva_mx0w0 <= STAGE_LOOP_lshift_rg_z;

  inPlaceNTT_DIT_core_core_fsm_inst : inPlaceNTT_DIT_core_core_fsm
    PORT MAP(
      clk => clk,
      rst => rst,
      fsm_output => inPlaceNTT_DIT_core_core_fsm_inst_fsm_output,
      STAGE_LOOP_C_8_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_8_tr0,
      modExp_while_C_38_tr0 => COMP_LOOP_COMP_LOOP_and_137_itm,
      COMP_LOOP_C_1_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_1_tr0,
      COMP_LOOP_1_modExp_1_while_C_38_tr0 => COMP_LOOP_COMP_LOOP_and_137_itm,
      COMP_LOOP_C_64_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_64_tr0,
      COMP_LOOP_2_modExp_1_while_C_38_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_2_modExp_1_while_C_38_tr0,
      COMP_LOOP_C_128_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_128_tr0,
      COMP_LOOP_3_modExp_1_while_C_38_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_3_modExp_1_while_C_38_tr0,
      COMP_LOOP_C_192_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_192_tr0,
      COMP_LOOP_4_modExp_1_while_C_38_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_4_modExp_1_while_C_38_tr0,
      COMP_LOOP_C_256_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_256_tr0,
      COMP_LOOP_5_modExp_1_while_C_38_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_5_modExp_1_while_C_38_tr0,
      COMP_LOOP_C_320_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_320_tr0,
      COMP_LOOP_6_modExp_1_while_C_38_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_6_modExp_1_while_C_38_tr0,
      COMP_LOOP_C_384_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_384_tr0,
      COMP_LOOP_7_modExp_1_while_C_38_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_7_modExp_1_while_C_38_tr0,
      COMP_LOOP_C_448_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_448_tr0,
      COMP_LOOP_8_modExp_1_while_C_38_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_8_modExp_1_while_C_38_tr0,
      COMP_LOOP_C_512_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_512_tr0,
      COMP_LOOP_9_modExp_1_while_C_38_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_9_modExp_1_while_C_38_tr0,
      COMP_LOOP_C_576_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_576_tr0,
      COMP_LOOP_10_modExp_1_while_C_38_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_10_modExp_1_while_C_38_tr0,
      COMP_LOOP_C_640_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_640_tr0,
      COMP_LOOP_11_modExp_1_while_C_38_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_11_modExp_1_while_C_38_tr0,
      COMP_LOOP_C_704_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_704_tr0,
      COMP_LOOP_12_modExp_1_while_C_38_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_12_modExp_1_while_C_38_tr0,
      COMP_LOOP_C_768_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_768_tr0,
      COMP_LOOP_13_modExp_1_while_C_38_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_13_modExp_1_while_C_38_tr0,
      COMP_LOOP_C_832_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_832_tr0,
      COMP_LOOP_14_modExp_1_while_C_38_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_14_modExp_1_while_C_38_tr0,
      COMP_LOOP_C_896_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_896_tr0,
      COMP_LOOP_15_modExp_1_while_C_38_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_15_modExp_1_while_C_38_tr0,
      COMP_LOOP_C_960_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_960_tr0,
      COMP_LOOP_16_modExp_1_while_C_38_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_16_modExp_1_while_C_38_tr0,
      COMP_LOOP_C_1024_tr0 => COMP_LOOP_COMP_LOOP_and_10_itm,
      VEC_LOOP_C_0_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_C_0_tr0,
      STAGE_LOOP_C_9_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_9_tr0
    );
  fsm_output <= inPlaceNTT_DIT_core_core_fsm_inst_fsm_output;
  inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_8_tr0 <= NOT (z_out_1(64));
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_1_tr0 <= NOT COMP_LOOP_nor_11_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_64_tr0 <= NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_2_modExp_1_while_C_38_tr0 <= NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_128_tr0 <= NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_3_modExp_1_while_C_38_tr0 <= NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_192_tr0 <= NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_4_modExp_1_while_C_38_tr0 <= NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_256_tr0 <= NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_5_modExp_1_while_C_38_tr0 <= NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_320_tr0 <= NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_6_modExp_1_while_C_38_tr0 <= NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_384_tr0 <= NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_7_modExp_1_while_C_38_tr0 <= NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_448_tr0 <= NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_8_modExp_1_while_C_38_tr0 <= NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_512_tr0 <= NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_9_modExp_1_while_C_38_tr0 <= NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_576_tr0 <= NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_10_modExp_1_while_C_38_tr0 <= NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_640_tr0 <= NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_11_modExp_1_while_C_38_tr0 <= NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_704_tr0 <= NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_12_modExp_1_while_C_38_tr0 <= NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_768_tr0 <= NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_13_modExp_1_while_C_38_tr0 <= NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_832_tr0 <= NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_14_modExp_1_while_C_38_tr0 <= NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_896_tr0 <= NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_15_modExp_1_while_C_38_tr0 <= NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_960_tr0 <= NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_16_modExp_1_while_C_38_tr0 <= NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_C_0_tr0 <= z_out(12);
  inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_9_tr0 <= NOT STAGE_LOOP_acc_itm_2_1;

  nor_1445_cse <= NOT((fsm_output(7)) OR (fsm_output(3)) OR (NOT (fsm_output(9)))
      OR (fsm_output(2)) OR (fsm_output(10)));
  or_651_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (NOT
      (fsm_output(2))) OR (fsm_output(10));
  or_650_nl <= (COMP_LOOP_acc_16_psp_sva(0)) OR (VEC_LOOP_j_sva_11_0(2)) OR (fsm_output(7))
      OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9))) OR (fsm_output(2)) OR (fsm_output(10));
  mux_1157_cse <= MUX_s_1_2_2(or_651_nl, or_650_nl, fsm_output(5));
  or_638_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9)))
      OR (fsm_output(2)) OR (fsm_output(10));
  or_637_nl <= (fsm_output(7)) OR CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_253;
  mux_1149_cse <= MUX_s_1_2_2(or_638_nl, or_637_nl, fsm_output(5));
  nand_332_cse <= NOT((VEC_LOOP_j_sva_11_0(0)) AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm);
  or_859_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9)))
      OR (fsm_output(2)) OR (fsm_output(10));
  or_858_nl <= (fsm_output(7)) OR CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_253;
  mux_1277_cse <= MUX_s_1_2_2(or_859_nl, or_858_nl, fsm_output(5));
  nand_324_cse <= NOT((NOT (fsm_output(1))) AND CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1
      DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm);
  or_1093_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (NOT
      (fsm_output(2))) OR (fsm_output(10));
  or_1092_nl <= (COMP_LOOP_acc_16_psp_sva(0)) OR (NOT (VEC_LOOP_j_sva_11_0(2))) OR
      (fsm_output(7)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9))) OR (fsm_output(2))
      OR (fsm_output(10));
  mux_1413_cse <= MUX_s_1_2_2(or_1093_nl, or_1092_nl, fsm_output(5));
  or_1080_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9)))
      OR (fsm_output(2)) OR (fsm_output(10));
  or_1079_nl <= (fsm_output(7)) OR CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO
      0)/=STD_LOGIC_VECTOR'("010")) OR (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_253;
  mux_1405_cse <= MUX_s_1_2_2(or_1080_nl, or_1079_nl, fsm_output(5));
  or_1301_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9)))
      OR (fsm_output(2)) OR (fsm_output(10));
  or_1300_nl <= (fsm_output(7)) OR CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO
      0)/=STD_LOGIC_VECTOR'("011")) OR (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_253;
  mux_1533_cse <= MUX_s_1_2_2(or_1301_nl, or_1300_nl, fsm_output(5));
  or_1535_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (NOT
      (fsm_output(2))) OR (fsm_output(10));
  or_1534_nl <= (NOT (COMP_LOOP_acc_16_psp_sva(0))) OR (VEC_LOOP_j_sva_11_0(2)) OR
      (fsm_output(7)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9))) OR (fsm_output(2))
      OR (fsm_output(10));
  mux_1669_cse <= MUX_s_1_2_2(or_1535_nl, or_1534_nl, fsm_output(5));
  or_1522_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9)))
      OR (fsm_output(2)) OR (fsm_output(10));
  or_1521_nl <= (fsm_output(7)) OR CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO
      0)/=STD_LOGIC_VECTOR'("100")) OR (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_253;
  mux_1661_cse <= MUX_s_1_2_2(or_1522_nl, or_1521_nl, fsm_output(5));
  or_1743_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9)))
      OR (fsm_output(2)) OR (fsm_output(10));
  or_1742_nl <= (fsm_output(7)) OR CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO
      0)/=STD_LOGIC_VECTOR'("101")) OR (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_253;
  mux_1789_cse <= MUX_s_1_2_2(or_1743_nl, or_1742_nl, fsm_output(5));
  nand_259_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND (fsm_output(7)) AND (fsm_output(3)) AND (NOT (fsm_output(9))) AND (fsm_output(2))
      AND (NOT (fsm_output(10))));
  or_1976_nl <= (NOT (COMP_LOOP_acc_16_psp_sva(0))) OR (NOT (VEC_LOOP_j_sva_11_0(2)))
      OR (fsm_output(7)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9))) OR (fsm_output(2))
      OR (fsm_output(10));
  mux_1925_cse <= MUX_s_1_2_2(nand_259_nl, or_1976_nl, fsm_output(5));
  or_1964_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9)))
      OR (fsm_output(2)) OR (fsm_output(10));
  or_1963_nl <= (fsm_output(7)) OR CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO
      0)/=STD_LOGIC_VECTOR'("110")) OR (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_253;
  mux_1917_cse <= MUX_s_1_2_2(or_1964_nl, or_1963_nl, fsm_output(5));
  nand_231_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"))
      AND (fsm_output(7)) AND (fsm_output(3)) AND (fsm_output(9)) AND (NOT (fsm_output(2)))
      AND (NOT (fsm_output(10))));
  or_2184_nl <= (fsm_output(7)) OR CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO
      0)/=STD_LOGIC_VECTOR'("111")) OR (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_253;
  mux_2045_cse <= MUX_s_1_2_2(nand_231_nl, or_2184_nl, fsm_output(5));
  or_3388_cse <= CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"));
  and_527_cse <= or_3388_cse AND (fsm_output(2));
  and_526_cse <= CONV_SL_1_1(fsm_output(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"));
  or_2377_cse <= and_526_cse OR (fsm_output(2));
  or_2368_cse <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("00"));
  and_529_cse <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)=STD_LOGIC_VECTOR'("11"));
  nor_758_cse <= NOT(CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("00")));
  nand_196_cse <= NOT(CONV_SL_1_1(fsm_output(2 DOWNTO 1)=STD_LOGIC_VECTOR'("11")));
  or_2419_cse <= (NOT (fsm_output(1))) OR (fsm_output(9));
  nor_297_cse <= NOT((fsm_output(0)) OR (fsm_output(1)) OR (NOT (fsm_output(9))));
  nor_303_cse <= NOT((fsm_output(1)) OR (NOT (fsm_output(9))));
  nor_1584_nl <= NOT((fsm_output(3)) OR (NOT (fsm_output(8))) OR (fsm_output(6))
      OR (NOT (fsm_output(10))));
  and_739_nl <= (fsm_output(3)) AND (fsm_output(8)) AND (fsm_output(6)) AND (NOT
      (fsm_output(10)));
  mux_125_cse <= MUX_s_1_2_2(nor_1584_nl, and_739_nl, fsm_output(7));
  and_536_cse <= CONV_SL_1_1(fsm_output(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"));
  nor_753_cse <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")));
  or_2387_cse <= CONV_SL_1_1(fsm_output(10 DOWNTO 8)/=STD_LOGIC_VECTOR'("110"));
  or_2414_cse <= CONV_SL_1_1(fsm_output(10 DOWNTO 9)/=STD_LOGIC_VECTOR'("00"));
  or_2407_cse <= CONV_SL_1_1(fsm_output(10 DOWNTO 8)/=STD_LOGIC_VECTOR'("010"));
  mux_2171_cse <= MUX_s_1_2_2((fsm_output(7)), or_tmp_2276, fsm_output(9));
  mux_2203_cse <= MUX_s_1_2_2(or_tmp_2281, (fsm_output(7)), fsm_output(9));
  or_2400_cse <= (NOT (fsm_output(0))) OR (NOT (fsm_output(1))) OR (fsm_output(9));
  and_521_cse <= (NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))))
      AND (fsm_output(9));
  or_2421_cse <= nor_753_cse OR (fsm_output(9));
  nand_356_cse <= NOT((fsm_output(5)) AND (fsm_output(7)) AND (fsm_output(9)) AND
      (fsm_output(10)));
  or_491_cse <= CONV_SL_1_1(fsm_output(4 DOWNTO 2)/=STD_LOGIC_VECTOR'("000"));
  nand_357_cse <= NOT((fsm_output(7)) AND (fsm_output(9)) AND (fsm_output(10)));
  nand_358_cse <= NOT(CONV_SL_1_1(fsm_output(10 DOWNTO 9)=STD_LOGIC_VECTOR'("11")));
  or_2921_cse <= (fsm_output(1)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(2)))
      OR (fsm_output(6)) OR (fsm_output(10));
  or_2918_cse <= (fsm_output(1)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(2)))
      OR (NOT (fsm_output(6))) OR (fsm_output(10));
  or_2912_cse <= (fsm_output(1)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(2)))
      OR (fsm_output(6)) OR (NOT (fsm_output(10)));
  or_2905_cse <= (NOT (fsm_output(1))) OR (NOT (fsm_output(9))) OR (fsm_output(2))
      OR (NOT (fsm_output(6))) OR (fsm_output(10));
  nor_697_cse <= NOT(and_526_cse OR (fsm_output(2)));
  mux_3254_cse <= MUX_s_1_2_2(or_2947_cse, or_2921_cse, fsm_output(0));
  mux_3245_cse <= MUX_s_1_2_2(mux_3281_cse, or_2905_cse, fsm_output(0));
  or_2914_cse <= (NOT (fsm_output(1))) OR (fsm_output(9)) OR (fsm_output(2)) OR (fsm_output(6))
      OR (NOT (fsm_output(10)));
  or_2920_nl <= (fsm_output(0)) OR (fsm_output(1)) OR (fsm_output(9)) OR (fsm_output(2))
      OR (fsm_output(6)) OR (NOT (fsm_output(10)));
  mux_3255_nl <= MUX_s_1_2_2(mux_3254_cse, or_2920_nl, fsm_output(3));
  nor_640_nl <= NOT((fsm_output(4)) OR (NOT (fsm_output(8))) OR mux_3255_nl);
  mux_3252_nl <= MUX_s_1_2_2(or_2918_cse, mux_3281_cse, fsm_output(0));
  and_421_nl <= (fsm_output(8)) AND (fsm_output(3)) AND (NOT mux_3252_nl);
  nor_642_nl <= NOT((fsm_output(2)) OR (fsm_output(6)) OR (fsm_output(10)));
  nor_643_nl <= NOT((NOT (fsm_output(2))) OR (fsm_output(6)) OR (fsm_output(10)));
  mux_3250_nl <= MUX_s_1_2_2(nor_642_nl, nor_643_nl, fsm_output(9));
  nand_85_nl <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND
      mux_3250_nl);
  mux_3249_nl <= MUX_s_1_2_2(or_2914_cse, or_2912_cse, fsm_output(0));
  mux_3251_nl <= MUX_s_1_2_2(nand_85_nl, mux_3249_nl, fsm_output(3));
  nor_641_nl <= NOT((fsm_output(8)) OR mux_3251_nl);
  mux_3253_nl <= MUX_s_1_2_2(and_421_nl, nor_641_nl, fsm_output(4));
  mux_3256_nl <= MUX_s_1_2_2(nor_640_nl, mux_3253_nl, fsm_output(5));
  or_2910_nl <= (NOT (fsm_output(1))) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(2)))
      OR (fsm_output(6)) OR (fsm_output(10));
  mux_3246_nl <= MUX_s_1_2_2(or_2910_nl, or_2947_cse, fsm_output(0));
  and_423_nl <= (fsm_output(3)) AND (NOT mux_3246_nl);
  nor_644_nl <= NOT((fsm_output(3)) OR mux_3245_cse);
  mux_3247_nl <= MUX_s_1_2_2(and_423_nl, nor_644_nl, fsm_output(8));
  and_422_nl <= (fsm_output(4)) AND mux_3247_nl;
  nor_645_nl <= NOT((fsm_output(4)) OR (fsm_output(8)) OR (fsm_output(3)) OR (NOT
      (fsm_output(0))) OR (fsm_output(1)) OR (fsm_output(9)) OR (fsm_output(2)) OR
      (fsm_output(6)) OR (NOT (fsm_output(10))));
  mux_3248_nl <= MUX_s_1_2_2(and_422_nl, nor_645_nl, fsm_output(5));
  mux_3257_nl <= MUX_s_1_2_2(mux_3256_nl, mux_3248_nl, fsm_output(7));
  and_323_nl <= mux_3257_nl AND COMP_LOOP_nor_11_itm;
  modExp_while_if_and_nl <= modExp_while_and_3 AND not_tmp_557;
  modExp_while_if_and_1_nl <= modExp_while_and_5 AND not_tmp_557;
  modExp_while_if_mux1h_nl <= MUX1HOT_v_64_6_2(z_out_8, STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000001"),
      COMP_LOOP_1_modExp_1_while_if_mul_mut_1, modulo_result_rem_cmp_z, modulo_qr_sva_1_mx0w6,
      COMP_LOOP_1_acc_5_mut_mx0w5, STD_LOGIC_VECTOR'( and_dcpl_237 & (NOT mux_2757_itm)
      & and_323_nl & modExp_while_if_and_nl & modExp_while_if_and_1_nl & not_tmp_441));
  and_261_nl <= and_dcpl_93 AND and_dcpl_127;
  or_2578_nl <= CONV_SL_1_1(fsm_output(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000")) OR
      (NOT nor_tmp_324);
  mux_2540_nl <= MUX_s_1_2_2(or_2578_nl, or_2541_cse, fsm_output(9));
  mux_2629_nl <= MUX_s_1_2_2((NOT or_tmp_2393), (fsm_output(5)), or_2368_cse);
  mux_2628_nl <= MUX_s_1_2_2((NOT or_tmp_2393), (fsm_output(5)), and_527_cse);
  mux_2630_nl <= MUX_s_1_2_2(mux_2629_nl, mux_2628_nl, fsm_output(9));
  mux_2541_nl <= MUX_s_1_2_2(mux_2540_nl, mux_2630_nl, fsm_output(6));
  or_2624_nl <= (NOT(and_526_cse OR (fsm_output(2)) OR (fsm_output(5)))) OR (fsm_output(10));
  mux_2609_nl <= MUX_s_1_2_2((NOT or_2534_cse), or_2624_nl, fsm_output(9));
  mux_2607_nl <= MUX_s_1_2_2(mux_2494_cse, mux_2516_cse, and_526_cse);
  or_2622_nl <= (NOT(CONV_SL_1_1(fsm_output(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))))
      OR (fsm_output(5)) OR (fsm_output(10));
  mux_2608_nl <= MUX_s_1_2_2(mux_2607_nl, or_2622_nl, fsm_output(9));
  mux_2610_nl <= MUX_s_1_2_2(mux_2609_nl, mux_2608_nl, fsm_output(6));
  mux_2542_nl <= MUX_s_1_2_2(mux_2541_nl, mux_2610_nl, fsm_output(8));
  mux_2615_nl <= MUX_s_1_2_2(nor_tmp_324, mux_2486_cse, and_527_cse);
  mux_2616_nl <= MUX_s_1_2_2((NOT or_2528_cse), mux_2615_nl, fsm_output(9));
  nor_696_nl <= NOT(nor_697_cse OR (fsm_output(5)) OR (fsm_output(10)));
  or_2627_nl <= (NOT((NOT (fsm_output(1))) OR (NOT (fsm_output(2))) OR (fsm_output(5))))
      OR (fsm_output(10));
  mux_2614_nl <= MUX_s_1_2_2(nor_696_nl, or_2627_nl, fsm_output(9));
  mux_2617_nl <= MUX_s_1_2_2(mux_2616_nl, mux_2614_nl, fsm_output(6));
  mux_2598_nl <= MUX_s_1_2_2((fsm_output(5)), nor_tmp_324, and_527_cse);
  mux_2599_nl <= MUX_s_1_2_2(mux_2598_nl, or_tmp_2474, fsm_output(9));
  mux_2600_nl <= MUX_s_1_2_2(mux_2599_nl, mux_2465_cse, fsm_output(6));
  mux_2532_nl <= MUX_s_1_2_2(mux_2617_nl, mux_2600_nl, fsm_output(8));
  mux_2543_nl <= MUX_s_1_2_2(mux_2542_nl, mux_2532_nl, fsm_output(7));
  mux_2520_nl <= MUX_s_1_2_2((fsm_output(5)), nor_tmp_324, or_2368_cse);
  mux_2623_nl <= MUX_s_1_2_2(mux_2494_cse, mux_2515_cse, fsm_output(1));
  mux_2622_nl <= MUX_s_1_2_2(mux_2516_cse, mux_2515_cse, fsm_output(1));
  mux_2624_nl <= MUX_s_1_2_2(mux_2623_nl, mux_2622_nl, fsm_output(0));
  mux_2521_nl <= MUX_s_1_2_2(mux_2520_nl, mux_2624_nl, fsm_output(9));
  mux_2619_nl <= MUX_s_1_2_2((fsm_output(5)), nor_tmp_324, or_2377_cse);
  mux_2620_nl <= MUX_s_1_2_2((NOT nand_173_cse), mux_2619_nl, fsm_output(9));
  mux_2522_nl <= MUX_s_1_2_2(mux_2521_nl, mux_2620_nl, fsm_output(6));
  mux_2603_nl <= MUX_s_1_2_2((fsm_output(5)), or_tmp_2474, fsm_output(9));
  mux_2586_nl <= MUX_s_1_2_2(or_tmp_2474, (fsm_output(5)), and_529_cse);
  or_2620_nl <= (NOT(nor_697_cse OR (fsm_output(5)))) OR (fsm_output(10));
  mux_2602_nl <= MUX_s_1_2_2((NOT mux_2586_nl), or_2620_nl, fsm_output(9));
  mux_2604_nl <= MUX_s_1_2_2(mux_2603_nl, mux_2602_nl, fsm_output(6));
  mux_2523_nl <= MUX_s_1_2_2(mux_2522_nl, mux_2604_nl, fsm_output(8));
  or_2625_nl <= (fsm_output(9)) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(1)))
      OR (NOT (fsm_output(2))) OR (fsm_output(5)) OR (fsm_output(10));
  mux_2613_nl <= MUX_s_1_2_2(mux_2465_cse, or_2625_nl, fsm_output(6));
  mux_2594_nl <= MUX_s_1_2_2(or_tmp_2474, nor_tmp_324, and_529_cse);
  mux_2595_nl <= MUX_s_1_2_2(or_2528_cse, mux_2594_nl, fsm_output(0));
  or_2616_nl <= (NOT((NOT (fsm_output(2))) OR (fsm_output(5)))) OR (fsm_output(10));
  mux_2596_nl <= MUX_s_1_2_2((NOT mux_2595_nl), or_2616_nl, fsm_output(9));
  nor_704_nl <= NOT((fsm_output(2)) OR (fsm_output(5)) OR (NOT (fsm_output(10))));
  or_2612_nl <= (NOT((fsm_output(0)) OR (fsm_output(1)) OR (fsm_output(2)) OR (fsm_output(5))))
      OR (fsm_output(10));
  mux_2593_nl <= MUX_s_1_2_2(nor_704_nl, or_2612_nl, fsm_output(9));
  mux_2597_nl <= MUX_s_1_2_2(mux_2596_nl, mux_2593_nl, fsm_output(6));
  mux_2508_nl <= MUX_s_1_2_2(mux_2613_nl, mux_2597_nl, fsm_output(8));
  mux_2524_nl <= MUX_s_1_2_2(mux_2523_nl, mux_2508_nl, fsm_output(7));
  mux_2544_nl <= MUX_s_1_2_2(mux_2543_nl, mux_2524_nl, fsm_output(4));
  mux_2495_nl <= MUX_s_1_2_2(or_2540_cse, mux_2494_cse, fsm_output(1));
  mux_2496_nl <= MUX_s_1_2_2(or_2528_cse, mux_2495_nl, fsm_output(0));
  mux_2497_nl <= MUX_s_1_2_2(mux_2496_nl, or_2540_cse, fsm_output(9));
  mux_2498_nl <= MUX_s_1_2_2(mux_2497_nl, (fsm_output(5)), fsm_output(6));
  nor_707_nl <= NOT(nor_758_cse OR (NOT (fsm_output(5))) OR (fsm_output(10)));
  or_2591_nl <= (or_3388_cse AND (fsm_output(2)) AND (fsm_output(5))) OR (fsm_output(10));
  mux_2560_nl <= MUX_s_1_2_2(nor_707_nl, or_2591_nl, fsm_output(9));
  or_2589_nl <= (NOT((fsm_output(1)) OR (fsm_output(2)) OR (NOT (fsm_output(5)))))
      OR (fsm_output(10));
  mux_2559_nl <= MUX_s_1_2_2((NOT nand_386_cse), or_2589_nl, fsm_output(9));
  mux_2561_nl <= MUX_s_1_2_2(mux_2560_nl, mux_2559_nl, fsm_output(6));
  mux_2499_nl <= MUX_s_1_2_2(mux_2498_nl, mux_2561_nl, fsm_output(8));
  mux_2574_nl <= MUX_s_1_2_2(mux_2486_cse, or_tmp_2393, or_2377_cse);
  mux_2575_nl <= MUX_s_1_2_2((NOT (fsm_output(5))), mux_2574_nl, fsm_output(9));
  mux_2570_nl <= MUX_s_1_2_2(or_tmp_2474, nor_tmp_324, or_2368_cse);
  mux_2571_nl <= MUX_s_1_2_2((NOT mux_2570_nl), nand_173_cse, fsm_output(0));
  or_2602_nl <= (fsm_output(2)) OR (NOT (fsm_output(5))) OR (fsm_output(10));
  mux_2572_nl <= MUX_s_1_2_2(mux_2571_nl, or_2602_nl, fsm_output(9));
  mux_2576_nl <= MUX_s_1_2_2(mux_2575_nl, mux_2572_nl, fsm_output(6));
  nor_709_nl <= NOT(and_526_cse OR (fsm_output(2)) OR (NOT nor_tmp_324));
  mux_2552_nl <= MUX_s_1_2_2(nor_709_nl, (fsm_output(10)), fsm_output(9));
  mux_2550_nl <= MUX_s_1_2_2((fsm_output(5)), or_tmp_2394, and_529_cse);
  mux_2551_nl <= MUX_s_1_2_2((NOT mux_2550_nl), or_tmp_2393, fsm_output(9));
  mux_2553_nl <= MUX_s_1_2_2(mux_2552_nl, mux_2551_nl, fsm_output(6));
  mux_2490_nl <= MUX_s_1_2_2(mux_2576_nl, mux_2553_nl, fsm_output(8));
  mux_2500_nl <= MUX_s_1_2_2(mux_2499_nl, mux_2490_nl, fsm_output(7));
  mux_2581_nl <= MUX_s_1_2_2((NOT nor_tmp_324), or_tmp_2474, fsm_output(2));
  mux_2582_nl <= MUX_s_1_2_2(or_2541_cse, mux_2581_nl, fsm_output(1));
  mux_2580_nl <= MUX_s_1_2_2(or_2541_cse, or_2540_cse, fsm_output(1));
  mux_2583_nl <= MUX_s_1_2_2(mux_2582_nl, mux_2580_nl, fsm_output(0));
  mux_2584_nl <= MUX_s_1_2_2(or_2540_cse, mux_2583_nl, fsm_output(9));
  or_2608_nl <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("00")) OR (NOT
      nor_tmp_324);
  or_2606_nl <= (NOT (fsm_output(1))) OR (NOT (fsm_output(2))) OR (fsm_output(5))
      OR (fsm_output(10));
  mux_2578_nl <= MUX_s_1_2_2(or_2608_nl, or_2606_nl, fsm_output(0));
  mux_2579_nl <= MUX_s_1_2_2(or_2540_cse, mux_2578_nl, fsm_output(9));
  mux_2585_nl <= MUX_s_1_2_2(mux_2584_nl, mux_2579_nl, fsm_output(6));
  mux_2556_nl <= MUX_s_1_2_2((fsm_output(5)), nor_tmp_324, and_529_cse);
  mux_2557_nl <= MUX_s_1_2_2(mux_2556_nl, or_tmp_2474, fsm_output(9));
  mux_2558_nl <= MUX_s_1_2_2(mux_2557_nl, mux_2465_cse, fsm_output(6));
  mux_2477_nl <= MUX_s_1_2_2((NOT mux_2585_nl), mux_2558_nl, fsm_output(8));
  mux_2566_nl <= MUX_s_1_2_2((fsm_output(5)), or_tmp_2394, or_2368_cse);
  mux_2567_nl <= MUX_s_1_2_2(mux_2566_nl, or_2534_cse, fsm_output(0));
  or_2598_nl <= (NOT((fsm_output(2)) OR (fsm_output(5)))) OR (fsm_output(10));
  mux_2568_nl <= MUX_s_1_2_2((NOT mux_2567_nl), or_2598_nl, fsm_output(9));
  mux_2564_nl <= MUX_s_1_2_2(or_tmp_2474, (fsm_output(5)), and_527_cse);
  mux_2565_nl <= MUX_s_1_2_2(mux_2564_nl, or_2528_cse, fsm_output(9));
  mux_2569_nl <= MUX_s_1_2_2(mux_2568_nl, mux_2565_nl, fsm_output(6));
  or_2582_nl <= (fsm_output(1)) OR (fsm_output(2)) OR (NOT (fsm_output(5))) OR (fsm_output(10));
  mux_2548_nl <= MUX_s_1_2_2(nand_386_cse, or_2582_nl, fsm_output(9));
  mux_2546_nl <= MUX_s_1_2_2((NOT or_tmp_2393), (fsm_output(5)), and_529_cse);
  or_2580_nl <= (or_2377_cse AND (fsm_output(5))) OR (fsm_output(10));
  mux_2547_nl <= MUX_s_1_2_2(mux_2546_nl, or_2580_nl, fsm_output(9));
  mux_2549_nl <= MUX_s_1_2_2(mux_2548_nl, mux_2547_nl, fsm_output(6));
  mux_2464_nl <= MUX_s_1_2_2(mux_2569_nl, mux_2549_nl, fsm_output(8));
  mux_2478_nl <= MUX_s_1_2_2(mux_2477_nl, mux_2464_nl, fsm_output(7));
  mux_2501_nl <= MUX_s_1_2_2(mux_2500_nl, mux_2478_nl, fsm_output(4));
  mux_2545_nl <= MUX_s_1_2_2(mux_2544_nl, mux_2501_nl, fsm_output(3));
  operator_64_false_mux1h_2_rgt <= MUX1HOT_v_65_3_2(z_out_6, (STD_LOGIC_VECTOR'(
      "00") & operator_64_false_slc_modExp_exp_63_1_3), ('0' & modExp_while_if_mux1h_nl),
      STD_LOGIC_VECTOR'( and_261_nl & and_dcpl_247 & (NOT mux_2545_nl)));
  or_3532_cse <= (fsm_output(6)) OR and_757_cse;
  or_3609_nl <= (NOT (fsm_output(10))) OR (fsm_output(6)) OR (NOT (fsm_output(2)))
      OR (fsm_output(9));
  mux_3935_cse <= MUX_s_1_2_2(or_2965_cse, or_3609_nl, fsm_output(1));
  mux_554_cse <= MUX_s_1_2_2((NOT (fsm_output(10))), (fsm_output(10)), fsm_output(6));
  or_181_cse <= (fsm_output(5)) OR (fsm_output(3));
  or_2644_cse <= CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00"));
  mux_544_cse <= MUX_s_1_2_2((NOT or_tmp_167), (fsm_output(10)), fsm_output(9));
  mux_2643_cse <= MUX_s_1_2_2(mux_tmp_2640, and_756_cse, fsm_output(6));
  and_273_m1c <= and_dcpl_147 AND and_dcpl_90 AND and_dcpl_107;
  and_756_cse <= (fsm_output(7)) AND (fsm_output(9)) AND (fsm_output(10));
  and_757_cse <= CONV_SL_1_1(fsm_output(10 DOWNTO 9)=STD_LOGIC_VECTOR'("11"));
  modExp_result_and_rgt <= (NOT modExp_while_and_5) AND and_273_m1c;
  modExp_result_and_1_rgt <= modExp_while_and_5 AND and_273_m1c;
  and_458_cse <= (fsm_output(7)) AND (fsm_output(9));
  and_459_cse <= CONV_SL_1_1(fsm_output(3 DOWNTO 1)=STD_LOGIC_VECTOR'("111"));
  nand_166_nl <= NOT((fsm_output(2)) AND (fsm_output(9)) AND (fsm_output(1)) AND
      (fsm_output(6)) AND (NOT (fsm_output(10))));
  mux_2769_nl <= MUX_s_1_2_2(nand_166_nl, or_tmp_2651, fsm_output(0));
  nor_678_nl <= NOT((NOT (fsm_output(4))) OR (fsm_output(8)) OR (NOT (fsm_output(3)))
      OR mux_2769_nl);
  or_2716_nl <= (NOT (fsm_output(2))) OR (NOT (fsm_output(9))) OR (fsm_output(1))
      OR not_tmp_49;
  or_2714_nl <= (fsm_output(2)) OR (fsm_output(9)) OR (fsm_output(1)) OR not_tmp_49;
  mux_2767_nl <= MUX_s_1_2_2(or_2716_nl, or_2714_nl, fsm_output(0));
  or_2717_nl <= (fsm_output(3)) OR mux_2767_nl;
  mux_2766_nl <= MUX_s_1_2_2(or_2921_cse, mux_tmp_2760, fsm_output(0));
  nand_58_nl <= NOT((fsm_output(3)) AND (NOT mux_2766_nl));
  mux_2768_nl <= MUX_s_1_2_2(or_2717_nl, nand_58_nl, fsm_output(8));
  nor_679_nl <= NOT((fsm_output(4)) OR mux_2768_nl);
  mux_2770_nl <= MUX_s_1_2_2(nor_678_nl, nor_679_nl, fsm_output(5));
  mux_2762_nl <= MUX_s_1_2_2(or_tmp_2651, or_2918_cse, fsm_output(0));
  or_2708_nl <= (fsm_output(0)) OR (fsm_output(2)) OR (fsm_output(9)) OR (fsm_output(1))
      OR not_tmp_49;
  mux_2763_nl <= MUX_s_1_2_2(mux_2762_nl, or_2708_nl, fsm_output(3));
  nor_680_nl <= NOT((fsm_output(8)) OR mux_2763_nl);
  or_2702_nl <= (fsm_output(2)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(1)))
      OR (fsm_output(6)) OR (fsm_output(10));
  mux_2761_nl <= MUX_s_1_2_2(mux_tmp_2760, or_2702_nl, fsm_output(0));
  nor_681_nl <= NOT((NOT (fsm_output(8))) OR (fsm_output(3)) OR mux_2761_nl);
  mux_2764_nl <= MUX_s_1_2_2(nor_680_nl, nor_681_nl, fsm_output(4));
  nor_682_nl <= NOT((NOT (fsm_output(0))) OR (NOT (fsm_output(2))) OR (fsm_output(9))
      OR (NOT (fsm_output(1))) OR (NOT (fsm_output(6))) OR (fsm_output(10)));
  nor_683_nl <= NOT((fsm_output(2)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(1)))
      OR (NOT (fsm_output(6))) OR (fsm_output(10)));
  nor_684_nl <= NOT((NOT (fsm_output(2))) OR (fsm_output(9)) OR (fsm_output(1)) OR
      not_tmp_49);
  mux_2758_nl <= MUX_s_1_2_2(nor_683_nl, nor_684_nl, fsm_output(0));
  mux_2759_nl <= MUX_s_1_2_2(nor_682_nl, mux_2758_nl, fsm_output(3));
  and_451_nl <= (fsm_output(4)) AND (fsm_output(8)) AND mux_2759_nl;
  mux_2765_nl <= MUX_s_1_2_2(mux_2764_nl, and_451_nl, fsm_output(5));
  mux_2771_m1c <= MUX_s_1_2_2(mux_2770_nl, mux_2765_nl, fsm_output(7));
  or_470_cse <= CONV_SL_1_1(fsm_output(9 DOWNTO 8)/=STD_LOGIC_VECTOR'("00"));
  or_469_cse <= CONV_SL_1_1(fsm_output(10 DOWNTO 8)/=STD_LOGIC_VECTOR'("100"));
  mux_2926_cse <= MUX_s_1_2_2((NOT (fsm_output(10))), (fsm_output(10)), fsm_output(7));
  mux_1036_cse <= MUX_s_1_2_2((NOT or_tmp_93), or_tmp_88, fsm_output(9));
  mux_981_cse <= MUX_s_1_2_2(or_tmp_94, or_tmp_93, fsm_output(9));
  nor_685_nl <= NOT((fsm_output(6)) OR (NOT (fsm_output(5))) OR (fsm_output(3)));
  nor_686_nl <= NOT((NOT (fsm_output(6))) OR (fsm_output(5)) OR (NOT (fsm_output(3))));
  mux_2743_nl <= MUX_s_1_2_2(nor_685_nl, nor_686_nl, fsm_output(0));
  and_317_m1c <= mux_2743_nl AND and_dcpl_245 AND (NOT (fsm_output(8))) AND (fsm_output(4))
      AND (NOT (fsm_output(1))) AND nor_609_cse;
  or_80_cse <= (fsm_output(9)) OR (fsm_output(2)) OR (fsm_output(5)) OR (NOT (fsm_output(7)))
      OR (fsm_output(3)) OR (fsm_output(8)) OR (NOT (fsm_output(6))) OR (fsm_output(10));
  nand_159_cse <= NOT((fsm_output(3)) AND (fsm_output(10)));
  nor_657_cse <= NOT((NOT (fsm_output(9))) OR (fsm_output(2)));
  nor_653_cse <= NOT((NOT((NOT (fsm_output(0))) OR (fsm_output(9)))) OR (fsm_output(2)));
  mux_498_cse <= MUX_s_1_2_2(mux_tmp_165, or_2991_cse, fsm_output(4));
  COMP_LOOP_or_32_cse <= and_dcpl_117 OR and_dcpl_130 OR and_dcpl_140 OR and_dcpl_149
      OR and_dcpl_155 OR and_dcpl_164 OR and_dcpl_171 OR and_dcpl_178 OR and_dcpl_185
      OR and_dcpl_189 OR and_dcpl_197 OR and_dcpl_202 OR and_dcpl_211 OR and_dcpl_219
      OR and_dcpl_226 OR and_dcpl_231;
  or_2855_cse <= (NOT (fsm_output(9))) OR (fsm_output(2));
  or_2991_cse <= CONV_SL_1_1(fsm_output(10 DOWNTO 8)/=STD_LOGIC_VECTOR'("001"));
  or_2998_cse <= CONV_SL_1_1(fsm_output(10 DOWNTO 8)/=STD_LOGIC_VECTOR'("000"));
  or_2947_cse <= (NOT (fsm_output(1))) OR (fsm_output(9)) OR (fsm_output(2)) OR (fsm_output(6))
      OR (fsm_output(10));
  or_3008_cse <= (fsm_output(9)) OR nand_138_cse;
  or_2962_nl <= (fsm_output(9)) OR (fsm_output(2)) OR (NOT (fsm_output(6))) OR (fsm_output(10));
  or_2961_nl <= (fsm_output(9)) OR nand_367_cse;
  mux_3281_cse <= MUX_s_1_2_2(or_2962_nl, or_2961_nl, fsm_output(1));
  or_2965_cse <= (fsm_output(9)) OR (fsm_output(2)) OR (fsm_output(6)) OR (fsm_output(10));
  nand_367_cse <= NOT((fsm_output(2)) AND (fsm_output(6)) AND (fsm_output(10)));
  and_407_cse <= CONV_SL_1_1(fsm_output(5 DOWNTO 4)=STD_LOGIC_VECTOR'("11"));
  or_3039_cse <= CONV_SL_1_1(fsm_output(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("000"));
  or_3427_cse <= (fsm_output(7)) OR (fsm_output(5));
  and_404_cse <= CONV_SL_1_1(fsm_output(8 DOWNTO 7)=STD_LOGIC_VECTOR'("11"));
  or_259_cse <= CONV_SL_1_1(fsm_output(9 DOWNTO 8)/=STD_LOGIC_VECTOR'("01"));
  and_676_cse <= (fsm_output(5)) AND (fsm_output(2));
  and_672_cse <= ((fsm_output(9)) OR (fsm_output(6))) AND (fsm_output(10));
  and_395_cse <= (fsm_output(7)) AND (fsm_output(10));
  or_3063_cse <= CONV_SL_1_1(fsm_output(5 DOWNTO 4)/=STD_LOGIC_VECTOR'("00"));
  or_352_cse <= (NOT (fsm_output(6))) OR (fsm_output(10));
  or_3417_cse <= (fsm_output(1)) OR (fsm_output(2)) OR (fsm_output(9)) OR (fsm_output(6));
  or_361_cse <= CONV_SL_1_1(fsm_output(10 DOWNTO 9)/=STD_LOGIC_VECTOR'("01"));
  or_3079_cse <= CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000"));
  or_3074_cse <= CONV_SL_1_1(fsm_output(8 DOWNTO 5)/=STD_LOGIC_VECTOR'("0000"));
  nor_609_cse <= NOT(CONV_SL_1_1(fsm_output(10 DOWNTO 9)/=STD_LOGIC_VECTOR'("00")));
  nand_142_cse <= NOT((fsm_output(8)) AND (fsm_output(6)) AND (fsm_output(10)));
  and_366_cse <= (fsm_output(2)) AND (fsm_output(4));
  nand_138_cse <= NOT((fsm_output(8)) AND (fsm_output(10)));
  mux_3555_cse <= MUX_s_1_2_2(or_tmp_93, (fsm_output(8)), fsm_output(9));
  and_350_cse <= (fsm_output(7)) AND (fsm_output(5));
  STAGE_LOOP_i_3_0_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(STAGE_LOOP_i_3_0_sva)
      + UNSIGNED'( "0001"), 4));
  COMP_LOOP_acc_psp_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_sva_11_0(11
      DOWNTO 4)) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0),
      5), 8), 8));
  COMP_LOOP_1_acc_5_mut_mx0w5 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_10_lpi_4_dfm)
      + SIGNED(COMP_LOOP_10_mul_mut), 64));
  COMP_LOOP_1_modExp_1_while_if_mul_mut_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED'(
      SIGNED(operator_64_false_acc_mut_63_0) * SIGNED(COMP_LOOP_10_mul_mut)), 64));
  operator_64_false_slc_modExp_exp_63_1_3 <= MUX_v_63_2_2((operator_66_true_div_cmp_z(63
      DOWNTO 1)), (tmp_10_lpi_4_dfm(63 DOWNTO 1)), and_dcpl_256);
  modulo_qr_sva_1_mx0w6 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_result_rem_cmp_z)
      + UNSIGNED(p_sva), 64));
  or_70_cse <= (fsm_output(2)) OR (fsm_output(6)) OR (NOT (fsm_output(1))) OR (NOT
      (fsm_output(8))) OR (fsm_output(4)) OR (NOT (fsm_output(9))) OR (fsm_output(10));
  or_56_cse <= (fsm_output(2)) OR (NOT (fsm_output(6))) OR (fsm_output(1)) OR (NOT
      (fsm_output(8))) OR (NOT (fsm_output(4))) OR (NOT (fsm_output(9))) OR (fsm_output(10));
  mux_340_cse <= MUX_s_1_2_2(mux_tmp_141, or_tmp_94, fsm_output(4));
  mux_375_cse <= MUX_s_1_2_2(mux_tmp_130, or_2998_cse, fsm_output(4));
  COMP_LOOP_acc_1_cse_6_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_sva_11_0)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0 & STD_LOGIC_VECTOR'(
      "0101")), 9), 12), 12));
  COMP_LOOP_acc_1_cse_2_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_sva_11_0)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0 & STD_LOGIC_VECTOR'(
      "0001")), 9), 12), 12));
  modExp_while_and_3 <= (NOT (modulo_result_rem_cmp_z(63))) AND COMP_LOOP_nor_11_itm;
  modExp_while_and_5 <= (modulo_result_rem_cmp_z(63)) AND COMP_LOOP_nor_11_itm;
  nor_tmp_4 <= (fsm_output(3)) AND (fsm_output(5));
  or_18_nl <= (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(5));
  mux_tmp_14 <= MUX_s_1_2_2((fsm_output(5)), or_18_nl, fsm_output(7));
  not_tmp_39 <= NOT((fsm_output(4)) AND (fsm_output(10)));
  or_tmp_68 <= (fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(3))) OR (fsm_output(8))
      OR (NOT (fsm_output(6))) OR (fsm_output(10));
  not_tmp_49 <= NOT((fsm_output(6)) AND (fsm_output(10)));
  or_84_nl <= (fsm_output(8)) OR not_tmp_49;
  or_83_nl <= (NOT (fsm_output(8))) OR (fsm_output(6)) OR (fsm_output(10));
  mux_tmp_119 <= MUX_s_1_2_2(or_84_nl, or_83_nl, fsm_output(3));
  or_tmp_88 <= (NOT (fsm_output(8))) OR (fsm_output(10));
  mux_tmp_130 <= MUX_s_1_2_2((NOT (fsm_output(8))), or_tmp_88, fsm_output(9));
  mux_tmp_131 <= MUX_s_1_2_2(or_2991_cse, mux_tmp_130, fsm_output(4));
  or_tmp_93 <= (fsm_output(8)) OR (NOT (fsm_output(10)));
  nand_tmp_4 <= NOT((fsm_output(4)) AND (NOT mux_tmp_130));
  or_tmp_94 <= (fsm_output(8)) OR (fsm_output(10));
  mux_tmp_139 <= MUX_s_1_2_2((fsm_output(8)), or_tmp_94, fsm_output(9));
  mux_tmp_141 <= MUX_s_1_2_2(nand_138_cse, or_tmp_88, fsm_output(9));
  or_tmp_96 <= (fsm_output(4)) OR mux_tmp_130;
  or_108_nl <= (NOT (fsm_output(4))) OR (fsm_output(9));
  mux_155_cse <= MUX_s_1_2_2((NOT (fsm_output(8))), or_tmp_88, or_108_nl);
  mux_161_cse <= MUX_s_1_2_2(mux_tmp_130, or_3008_cse, fsm_output(4));
  mux_tmp_165 <= MUX_s_1_2_2(or_tmp_93, or_tmp_94, fsm_output(9));
  mux_171_cse <= MUX_s_1_2_2(or_469_cse, or_tmp_88, fsm_output(4));
  or_tmp_104 <= CONV_SL_1_1(fsm_output(10 DOWNTO 9)/=STD_LOGIC_VECTOR'("10"));
  mux_tmp_214 <= MUX_s_1_2_2(and_757_cse, or_tmp_104, fsm_output(5));
  mux_tmp_215 <= MUX_s_1_2_2(or_2414_cse, and_757_cse, fsm_output(5));
  nand_tmp_7 <= NOT((fsm_output(5)) AND (NOT and_757_cse));
  mux_tmp_227 <= MUX_s_1_2_2((NOT (fsm_output(10))), (fsm_output(10)), fsm_output(9));
  nor_tmp_23 <= ((NOT (fsm_output(5))) OR (fsm_output(9))) AND (fsm_output(10));
  mux_tmp_228 <= MUX_s_1_2_2(or_tmp_104, and_757_cse, fsm_output(5));
  mux_tmp_231 <= MUX_s_1_2_2(and_757_cse, or_2414_cse, fsm_output(5));
  mux_tmp_236 <= MUX_s_1_2_2(and_757_cse, mux_tmp_227, fsm_output(5));
  or_tmp_114 <= (fsm_output(5)) OR and_757_cse;
  mux_259_cse <= MUX_s_1_2_2((fsm_output(9)), and_757_cse, fsm_output(5));
  or_163_cse <= (NOT (fsm_output(4))) OR (fsm_output(8));
  and_dcpl_1 <= (NOT (fsm_output(4))) AND (fsm_output(1));
  and_dcpl_2 <= and_dcpl_1 AND (fsm_output(0));
  and_dcpl_4 <= CONV_SL_1_1(fsm_output(8 DOWNTO 7)=STD_LOGIC_VECTOR'("01"));
  and_dcpl_5 <= and_dcpl_4 AND (fsm_output(6));
  and_dcpl_6 <= nor_tmp_4 AND (NOT (fsm_output(2)));
  nor_1580_cse <= NOT((fsm_output(5)) OR (fsm_output(7)));
  not_tmp_90 <= NOT(CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00")));
  or_tmp_167 <= (fsm_output(6)) OR (fsm_output(10));
  nor_tmp_48 <= (fsm_output(6)) AND (fsm_output(10));
  and_707_cse <= (fsm_output(5)) AND (fsm_output(8));
  mux_648_cse <= MUX_s_1_2_2((NOT (fsm_output(8))), and_707_cse, fsm_output(6));
  or_tmp_222 <= (fsm_output(5)) OR (fsm_output(8));
  not_tmp_133 <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("00")));
  nor_tmp_82 <= CONV_SL_1_1(fsm_output(9 DOWNTO 8)=STD_LOGIC_VECTOR'("11"));
  or_tmp_258 <= (fsm_output(7)) OR (fsm_output(9));
  and_dcpl_19 <= (fsm_output(4)) AND (fsm_output(1));
  and_dcpl_26 <= (fsm_output(4)) AND (NOT (fsm_output(1)));
  and_dcpl_27 <= and_dcpl_26 AND (fsm_output(0));
  and_dcpl_33 <= CONV_SL_1_1(fsm_output(10 DOWNTO 9)=STD_LOGIC_VECTOR'("01"));
  and_dcpl_34 <= NOT((fsm_output(4)) OR (fsm_output(1)));
  and_dcpl_39 <= (fsm_output(5)) AND (NOT (fsm_output(3)));
  and_dcpl_40 <= and_dcpl_39 AND (NOT (fsm_output(2)));
  and_dcpl_44 <= and_dcpl_4 AND (NOT (fsm_output(6)));
  and_dcpl_48 <= and_dcpl_1 AND (NOT (fsm_output(0)));
  and_dcpl_55 <= and_dcpl_26 AND (NOT (fsm_output(0)));
  and_dcpl_59 <= CONV_SL_1_1(fsm_output(10 DOWNTO 9)=STD_LOGIC_VECTOR'("10"));
  or_3394_nl <= (fsm_output(0)) OR (fsm_output(1)) OR (fsm_output(5)) OR (fsm_output(7))
      OR (fsm_output(9)) OR (fsm_output(10));
  mux_1077_nl <= MUX_s_1_2_2(or_3394_nl, nand_356_cse, or_491_cse);
  mux_1078_nl <= MUX_s_1_2_2(mux_1077_nl, nand_357_cse, fsm_output(6));
  not_tmp_208 <= MUX_s_1_2_2(mux_1078_nl, nand_358_cse, fsm_output(8));
  and_dcpl_87 <= and_dcpl_34 AND (NOT (fsm_output(0)));
  and_dcpl_88 <= and_dcpl_87 AND nor_609_cse;
  and_dcpl_90 <= not_tmp_133 AND (NOT (fsm_output(6)));
  and_dcpl_91 <= NOT((fsm_output(3)) OR (fsm_output(5)));
  and_dcpl_92 <= and_dcpl_91 AND (NOT (fsm_output(2)));
  and_dcpl_93 <= and_dcpl_92 AND and_dcpl_90;
  and_dcpl_98 <= and_dcpl_2 AND and_757_cse;
  and_dcpl_103 <= and_dcpl_40 AND and_dcpl_44;
  and_dcpl_107 <= and_dcpl_27 AND nor_609_cse;
  and_dcpl_108 <= and_dcpl_40 AND and_dcpl_90;
  and_dcpl_109 <= and_dcpl_108 AND and_dcpl_107;
  and_dcpl_111 <= and_dcpl_19 AND (NOT (fsm_output(0)));
  and_dcpl_112 <= and_dcpl_111 AND nor_609_cse;
  and_dcpl_113 <= not_tmp_133 AND (fsm_output(6));
  and_dcpl_114 <= (fsm_output(3)) AND (NOT (fsm_output(5)));
  and_dcpl_115 <= and_dcpl_114 AND (NOT (fsm_output(2)));
  and_dcpl_117 <= and_dcpl_115 AND and_dcpl_113 AND and_dcpl_112;
  and_dcpl_118 <= and_dcpl_91 AND (fsm_output(2));
  or_tmp_453 <= (fsm_output(1)) OR (NOT (fsm_output(6))) OR (fsm_output(4)) OR (NOT
      (fsm_output(8))) OR (fsm_output(10));
  or_510_nl <= (NOT (fsm_output(0))) OR (NOT (fsm_output(1))) OR (fsm_output(6))
      OR (NOT (fsm_output(4))) OR (fsm_output(8)) OR (fsm_output(10));
  or_508_nl <= (fsm_output(1)) OR (fsm_output(6)) OR (NOT (fsm_output(4))) OR (fsm_output(8))
      OR (NOT (fsm_output(10)));
  mux_1081_nl <= MUX_s_1_2_2(or_tmp_453, or_508_nl, fsm_output(0));
  mux_tmp_1082 <= MUX_s_1_2_2(or_510_nl, mux_1081_nl, fsm_output(3));
  and_dcpl_126 <= and_dcpl_34 AND (fsm_output(0));
  and_dcpl_127 <= and_dcpl_126 AND nor_609_cse;
  and_dcpl_130 <= and_dcpl_92 AND and_dcpl_5 AND and_dcpl_127;
  and_dcpl_135 <= CONV_SL_1_1(fsm_output(8 DOWNTO 7)=STD_LOGIC_VECTOR'("10"));
  and_dcpl_136 <= and_dcpl_135 AND (NOT (fsm_output(6)));
  and_dcpl_139 <= and_dcpl_6 AND and_dcpl_136;
  and_dcpl_140 <= and_dcpl_139 AND and_dcpl_88;
  and_dcpl_144 <= and_dcpl_2 AND nor_609_cse;
  and_dcpl_146 <= and_404_cse AND (NOT (fsm_output(6)));
  and_dcpl_147 <= and_dcpl_114 AND (fsm_output(2));
  and_dcpl_149 <= and_dcpl_147 AND and_dcpl_146 AND and_dcpl_144;
  and_dcpl_152 <= and_404_cse AND (fsm_output(6));
  and_dcpl_153 <= and_dcpl_39 AND (fsm_output(2));
  and_dcpl_155 <= and_dcpl_153 AND and_dcpl_152 AND and_dcpl_112;
  and_dcpl_162 <= and_dcpl_27 AND and_dcpl_33;
  and_dcpl_164 <= and_dcpl_147 AND and_dcpl_113 AND and_dcpl_162;
  and_dcpl_170 <= and_dcpl_118 AND and_dcpl_5;
  and_dcpl_171 <= and_dcpl_170 AND and_dcpl_87 AND and_dcpl_33;
  and_dcpl_177 <= and_dcpl_2 AND and_dcpl_33;
  and_dcpl_178 <= and_dcpl_139 AND and_dcpl_177;
  and_dcpl_185 <= and_dcpl_92 AND and_dcpl_146 AND and_dcpl_111 AND and_dcpl_33;
  and_dcpl_189 <= and_dcpl_6 AND and_dcpl_152 AND and_dcpl_162;
  and_dcpl_191 <= NOT((fsm_output(8)) OR (fsm_output(6)));
  and_dcpl_196 <= and_dcpl_40 AND and_dcpl_113;
  and_dcpl_197 <= and_dcpl_196 AND and_dcpl_87 AND and_dcpl_59;
  and_dcpl_202 <= and_dcpl_170 AND and_dcpl_2 AND and_dcpl_59;
  and_dcpl_208 <= and_dcpl_48 AND and_dcpl_59;
  and_dcpl_209 <= nor_tmp_4 AND (fsm_output(2));
  and_dcpl_211 <= and_dcpl_209 AND and_dcpl_136 AND and_dcpl_208;
  and_dcpl_219 <= and_dcpl_118 AND and_dcpl_146 AND and_dcpl_27 AND and_dcpl_59;
  and_dcpl_224 <= and_dcpl_55 AND and_dcpl_59;
  and_dcpl_226 <= and_dcpl_209 AND and_dcpl_152 AND and_dcpl_224;
  and_dcpl_231 <= and_dcpl_196 AND and_dcpl_98;
  not_tmp_248 <= NOT((fsm_output(5)) AND (fsm_output(10)));
  or_580_nl <= (fsm_output(7)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(5)))
      OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(10));
  or_579_nl <= (NOT (fsm_output(7))) OR (fsm_output(9)) OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")) OR (fsm_output(10));
  mux_tmp_1116 <= MUX_s_1_2_2(or_580_nl, or_579_nl, fsm_output(2));
  or_tmp_532 <= (NOT (fsm_output(7))) OR (fsm_output(9)) OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")) OR (NOT (fsm_output(10)));
  or_586_cse <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"));
  or_591_cse <= (VEC_LOOP_j_sva_11_0(0)) OR (fsm_output(9)) OR (fsm_output(5)) OR
      (fsm_output(10));
  nand_337_cse <= NOT((fsm_output(9)) AND (fsm_output(5)) AND (fsm_output(10)));
  not_tmp_253 <= NOT((fsm_output(2)) AND (fsm_output(10)));
  or_691_nl <= (fsm_output(7)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(5)))
      OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(10));
  or_690_nl <= (NOT (fsm_output(7))) OR (fsm_output(9)) OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0001")) OR (fsm_output(10));
  mux_tmp_1180 <= MUX_s_1_2_2(or_691_nl, or_690_nl, fsm_output(2));
  or_tmp_643 <= (NOT (fsm_output(7))) OR (fsm_output(9)) OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0001")) OR (NOT (fsm_output(10)));
  nand_334_cse <= NOT((VEC_LOOP_j_sva_11_0(0)) AND (fsm_output(9)) AND (fsm_output(5))
      AND (fsm_output(10)));
  or_702_cse <= (NOT (VEC_LOOP_j_sva_11_0(0))) OR (fsm_output(9)) OR (fsm_output(5))
      OR (fsm_output(10));
  or_802_nl <= (fsm_output(7)) OR (NOT (fsm_output(5))) OR (NOT (fsm_output(9)))
      OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(10));
  or_801_nl <= (NOT (fsm_output(7))) OR (fsm_output(5)) OR (fsm_output(9)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0010")) OR (fsm_output(10));
  mux_tmp_1244 <= MUX_s_1_2_2(or_802_nl, or_801_nl, fsm_output(2));
  or_tmp_756 <= (NOT (fsm_output(7))) OR (fsm_output(5)) OR (fsm_output(9)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0010")) OR (NOT (fsm_output(10)));
  nor_209_cse <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001")));
  or_912_nl <= (fsm_output(7)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(5)))
      OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(10));
  or_911_nl <= (NOT (fsm_output(7))) OR (fsm_output(9)) OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0011")) OR (fsm_output(10));
  mux_tmp_1308 <= MUX_s_1_2_2(or_912_nl, or_911_nl, fsm_output(2));
  or_tmp_866 <= (NOT (fsm_output(7))) OR (fsm_output(9)) OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0011")) OR (NOT (fsm_output(10)));
  or_1022_nl <= (fsm_output(7)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(5)))
      OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(10));
  or_1021_nl <= (NOT (fsm_output(7))) OR (fsm_output(9)) OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0100")) OR (fsm_output(10));
  mux_tmp_1372 <= MUX_s_1_2_2(or_1022_nl, or_1021_nl, fsm_output(2));
  or_tmp_974 <= (NOT (fsm_output(7))) OR (fsm_output(9)) OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0100")) OR (NOT (fsm_output(10)));
  or_1028_cse <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"));
  or_1133_nl <= (fsm_output(7)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(5)))
      OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(10));
  or_1132_nl <= (NOT (fsm_output(7))) OR (fsm_output(9)) OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0101")) OR (fsm_output(10));
  mux_tmp_1436 <= MUX_s_1_2_2(or_1133_nl, or_1132_nl, fsm_output(2));
  or_tmp_1085 <= (NOT (fsm_output(7))) OR (fsm_output(9)) OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0101")) OR (NOT (fsm_output(10)));
  or_1244_nl <= (fsm_output(7)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(5)))
      OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(10));
  or_1243_nl <= (NOT (fsm_output(7))) OR (fsm_output(9)) OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0110")) OR (fsm_output(10));
  mux_tmp_1500 <= MUX_s_1_2_2(or_1244_nl, or_1243_nl, fsm_output(2));
  or_tmp_1198 <= (NOT (fsm_output(7))) OR (fsm_output(9)) OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0110")) OR (NOT (fsm_output(10)));
  nor_223_cse <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011")));
  or_1354_nl <= (fsm_output(7)) OR (NOT (fsm_output(5))) OR (NOT (fsm_output(9)))
      OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(10));
  or_1353_nl <= (NOT (fsm_output(7))) OR (fsm_output(5)) OR (fsm_output(9)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0111")) OR (fsm_output(10));
  mux_tmp_1564 <= MUX_s_1_2_2(or_1354_nl, or_1353_nl, fsm_output(2));
  or_tmp_1308 <= (NOT (fsm_output(7))) OR (fsm_output(5)) OR (fsm_output(9)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0111")) OR (NOT (fsm_output(10)));
  not_tmp_318 <= NOT((COMP_LOOP_acc_10_cse_12_1_1_sva(3)) AND (fsm_output(10)));
  or_1464_nl <= (fsm_output(7)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(5)))
      OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(10));
  or_1463_nl <= (NOT (fsm_output(7))) OR (fsm_output(9)) OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1000")) OR (fsm_output(10));
  mux_tmp_1628 <= MUX_s_1_2_2(or_1464_nl, or_1463_nl, fsm_output(2));
  or_tmp_1416 <= (NOT (fsm_output(7))) OR (fsm_output(9)) OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000")) OR not_tmp_318;
  or_1470_cse <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"));
  or_1575_nl <= (fsm_output(7)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(5)))
      OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(10));
  or_1574_nl <= (NOT (fsm_output(7))) OR (fsm_output(9)) OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1001")) OR (fsm_output(10));
  mux_tmp_1692 <= MUX_s_1_2_2(or_1575_nl, or_1574_nl, fsm_output(2));
  or_tmp_1527 <= (NOT (fsm_output(7))) OR (fsm_output(9)) OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001")) OR not_tmp_318;
  or_1686_nl <= (fsm_output(7)) OR (NOT (fsm_output(5))) OR (NOT (fsm_output(9)))
      OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(10));
  or_1685_nl <= (NOT (fsm_output(7))) OR (fsm_output(5)) OR (fsm_output(9)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1010")) OR (fsm_output(10));
  mux_tmp_1756 <= MUX_s_1_2_2(or_1686_nl, or_1685_nl, fsm_output(2));
  or_tmp_1640 <= (NOT (fsm_output(7))) OR (fsm_output(5)) OR (fsm_output(9)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010")) OR not_tmp_318;
  nor_239_cse <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101")));
  or_1796_nl <= (fsm_output(7)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(5)))
      OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(10));
  or_1795_nl <= (NOT (fsm_output(7))) OR (fsm_output(9)) OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1011")) OR (fsm_output(10));
  mux_tmp_1820 <= MUX_s_1_2_2(or_1796_nl, or_1795_nl, fsm_output(2));
  or_tmp_1750 <= (NOT (fsm_output(7))) OR (fsm_output(9)) OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("011")) OR not_tmp_318;
  not_tmp_357 <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 2)=STD_LOGIC_VECTOR'("11"))
      AND (fsm_output(10)));
  or_1906_nl <= (fsm_output(7)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(5)))
      OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(10));
  or_1905_nl <= (NOT (fsm_output(7))) OR (fsm_output(9)) OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1100")) OR (fsm_output(10));
  mux_tmp_1884 <= MUX_s_1_2_2(or_1906_nl, or_1905_nl, fsm_output(2));
  or_tmp_1858 <= (NOT (fsm_output(7))) OR (fsm_output(9)) OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR not_tmp_357;
  or_1912_cse <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"));
  or_2017_nl <= (fsm_output(7)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(5)))
      OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(10));
  or_2016_nl <= (NOT (fsm_output(7))) OR (fsm_output(9)) OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1101")) OR (fsm_output(10));
  mux_tmp_1948 <= MUX_s_1_2_2(or_2017_nl, or_2016_nl, fsm_output(2));
  or_tmp_1969 <= (NOT (fsm_output(7))) OR (fsm_output(9)) OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR not_tmp_357;
  not_tmp_377 <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 1)=STD_LOGIC_VECTOR'("111"))
      AND (fsm_output(10)));
  or_2128_nl <= (fsm_output(7)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(5)))
      OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(10));
  or_2127_nl <= (NOT (fsm_output(7))) OR (fsm_output(9)) OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1110")) OR (fsm_output(10));
  mux_tmp_2012 <= MUX_s_1_2_2(or_2128_nl, or_2127_nl, fsm_output(2));
  or_tmp_2082 <= (NOT (fsm_output(7))) OR (fsm_output(9)) OR (fsm_output(5)) OR (COMP_LOOP_acc_10_cse_12_1_1_sva(0))
      OR not_tmp_377;
  and_564_cse <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"));
  not_tmp_387 <= NOT((fsm_output(5)) AND CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)=STD_LOGIC_VECTOR'("1111")) AND (fsm_output(10)));
  nand_225_nl <= NOT((NOT (fsm_output(7))) AND (fsm_output(9)) AND (fsm_output(5))
      AND CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (NOT (fsm_output(10))));
  or_2237_nl <= (NOT (fsm_output(7))) OR (fsm_output(9)) OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1111")) OR (fsm_output(10));
  mux_tmp_2076 <= MUX_s_1_2_2(nand_225_nl, or_2237_nl, fsm_output(2));
  not_tmp_390 <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (fsm_output(10)));
  or_tmp_2192 <= (NOT (fsm_output(7))) OR (fsm_output(9)) OR (fsm_output(5)) OR not_tmp_390;
  nor_tmp_265 <= (fsm_output(9)) AND (fsm_output(5)) AND CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)=STD_LOGIC_VECTOR'("1111")) AND (fsm_output(10));
  and_dcpl_235 <= and_dcpl_48 AND nor_609_cse;
  and_dcpl_236 <= and_dcpl_115 AND and_dcpl_90;
  and_dcpl_237 <= and_dcpl_236 AND and_dcpl_235;
  or_tmp_2274 <= (NOT (fsm_output(1))) OR (NOT (fsm_output(2))) OR (fsm_output(7))
      OR (fsm_output(10));
  or_tmp_2276 <= (fsm_output(7)) OR (fsm_output(10));
  or_tmp_2277 <= and_526_cse OR (fsm_output(2)) OR (NOT (fsm_output(7))) OR (fsm_output(10));
  or_tmp_2280 <= (NOT (fsm_output(7))) OR (fsm_output(10));
  or_tmp_2281 <= (fsm_output(7)) OR (NOT (fsm_output(10)));
  mux_tmp_2159 <= MUX_s_1_2_2((NOT (fsm_output(7))), or_tmp_2280, fsm_output(9));
  or_tmp_2294 <= nor_753_cse OR (NOT (fsm_output(2))) OR (NOT (fsm_output(7))) OR
      (fsm_output(10));
  mux_tmp_2172 <= MUX_s_1_2_2((fsm_output(7)), and_395_cse, and_529_cse);
  or_tmp_2297 <= nor_758_cse OR (fsm_output(7)) OR (fsm_output(10));
  mux_2175_nl <= MUX_s_1_2_2(or_tmp_2276, (fsm_output(7)), and_529_cse);
  mux_tmp_2176 <= MUX_s_1_2_2(or_tmp_2297, mux_2175_nl, fsm_output(0));
  mux_tmp_2178 <= MUX_s_1_2_2((NOT and_395_cse), or_tmp_2276, fsm_output(2));
  or_tmp_2302 <= (NOT (fsm_output(2))) OR (fsm_output(7)) OR (fsm_output(10));
  mux_2234_nl <= MUX_s_1_2_2(mux_tmp_139, mux_tmp_165, or_3388_cse);
  mux_tmp_2235 <= MUX_s_1_2_2(mux_tmp_139, mux_2234_nl, fsm_output(3));
  mux_2239_nl <= MUX_s_1_2_2(mux_tmp_141, or_3008_cse, fsm_output(1));
  mux_tmp_2241 <= MUX_s_1_2_2(mux_tmp_130, mux_2239_nl, fsm_output(3));
  or_tmp_2340 <= nor_303_cse OR (fsm_output(8)) OR (fsm_output(10));
  or_tmp_2341 <= (NOT (fsm_output(1))) OR (fsm_output(9)) OR (fsm_output(8)) OR (fsm_output(10));
  mux_tmp_2262 <= MUX_s_1_2_2(mux_tmp_141, or_3008_cse, and_526_cse);
  and_524_cse <= (fsm_output(3)) AND (fsm_output(0)) AND (fsm_output(1));
  mux_tmp_2287 <= MUX_s_1_2_2(mux_tmp_130, mux_tmp_141, and_524_cse);
  mux_tmp_2289 <= MUX_s_1_2_2(or_tmp_93, (fsm_output(8)), nor_303_cse);
  mux_tmp_2293 <= MUX_s_1_2_2(or_259_cse, or_2991_cse, fsm_output(1));
  or_tmp_2360 <= (fsm_output(1)) OR (fsm_output(9)) OR nand_138_cse;
  mux_tmp_2311 <= MUX_s_1_2_2(or_3008_cse, or_2991_cse, fsm_output(1));
  or_tmp_2376 <= (fsm_output(4)) OR (NOT (fsm_output(7))) OR (fsm_output(3)) OR (fsm_output(8))
      OR (NOT (fsm_output(6))) OR (fsm_output(10));
  or_tmp_2389 <= (NOT (fsm_output(8))) OR (NOT (fsm_output(5))) OR (fsm_output(10));
  nand_188_nl <= NOT((fsm_output(8)) AND (fsm_output(5)));
  mux_tmp_2347 <= MUX_s_1_2_2(nand_188_nl, or_tmp_2389, fsm_output(9));
  or_tmp_2390 <= (NOT (fsm_output(8))) OR (fsm_output(5)) OR (fsm_output(10));
  or_2447_nl <= (NOT (fsm_output(8))) OR (fsm_output(5));
  mux_tmp_2348 <= MUX_s_1_2_2(or_2447_nl, or_tmp_2390, fsm_output(9));
  mux_tmp_2350 <= MUX_s_1_2_2(mux_tmp_2348, or_tmp_2389, fsm_output(6));
  not_tmp_431 <= NOT((fsm_output(8)) AND (fsm_output(5)) AND (fsm_output(10)));
  mux_2352_nl <= MUX_s_1_2_2(not_tmp_431, or_tmp_2389, fsm_output(9));
  or_2448_nl <= (fsm_output(9)) OR (fsm_output(8)) OR (fsm_output(5)) OR (fsm_output(10));
  mux_tmp_2353 <= MUX_s_1_2_2(mux_2352_nl, or_2448_nl, fsm_output(6));
  or_tmp_2393 <= (NOT (fsm_output(5))) OR (fsm_output(10));
  or_tmp_2394 <= (fsm_output(5)) OR (NOT (fsm_output(10)));
  mux_tmp_2355 <= MUX_s_1_2_2(or_tmp_2394, or_tmp_2393, fsm_output(8));
  or_2451_nl <= (fsm_output(9)) OR mux_tmp_2355;
  mux_tmp_2356 <= MUX_s_1_2_2(mux_tmp_2348, or_2451_nl, fsm_output(6));
  or_tmp_2396 <= (fsm_output(6)) OR mux_tmp_2347;
  or_tmp_2397 <= (fsm_output(8)) OR (fsm_output(5)) OR (fsm_output(10));
  or_tmp_2399 <= (fsm_output(8)) OR (fsm_output(5)) OR (NOT (fsm_output(10)));
  mux_tmp_2359 <= MUX_s_1_2_2(or_tmp_2399, or_tmp_2397, fsm_output(9));
  or_2457_nl <= CONV_SL_1_1(fsm_output(9 DOWNTO 8)/=STD_LOGIC_VECTOR'("10")) OR not_tmp_248;
  mux_tmp_2361 <= MUX_s_1_2_2(mux_tmp_2347, or_2457_nl, fsm_output(6));
  mux_tmp_2363 <= MUX_s_1_2_2(or_tmp_222, or_tmp_2397, fsm_output(9));
  or_2459_nl <= (fsm_output(9)) OR (NOT (fsm_output(8))) OR (fsm_output(5)) OR (fsm_output(10));
  mux_tmp_2364 <= MUX_s_1_2_2(or_2459_nl, mux_tmp_2363, fsm_output(6));
  or_tmp_2404 <= (fsm_output(8)) OR not_tmp_248;
  mux_tmp_2365 <= MUX_s_1_2_2(mux_tmp_2347, or_tmp_2404, fsm_output(6));
  nand_tmp_54 <= NOT((fsm_output(6)) AND (NOT mux_tmp_2363));
  or_tmp_2405 <= (fsm_output(8)) OR (NOT (fsm_output(5)));
  mux_tmp_2369 <= MUX_s_1_2_2(or_tmp_2404, or_tmp_2405, fsm_output(9));
  mux_tmp_2370 <= MUX_s_1_2_2(or_tmp_2389, mux_tmp_2355, fsm_output(9));
  mux_tmp_2371 <= MUX_s_1_2_2(mux_tmp_2370, mux_tmp_2369, fsm_output(6));
  mux_2375_nl <= MUX_s_1_2_2(mux_tmp_2355, or_tmp_2399, fsm_output(9));
  mux_tmp_2376 <= MUX_s_1_2_2(mux_2375_nl, or_tmp_2405, fsm_output(6));
  mux_tmp_2377 <= MUX_s_1_2_2(or_tmp_2399, or_tmp_222, fsm_output(9));
  mux_tmp_2378 <= MUX_s_1_2_2(mux_tmp_2377, or_tmp_2405, fsm_output(6));
  or_2462_nl <= (fsm_output(9)) OR not_tmp_431;
  mux_tmp_2382 <= MUX_s_1_2_2(or_2462_nl, or_tmp_2397, fsm_output(6));
  or_tmp_2407 <= (fsm_output(8)) OR (NOT (fsm_output(5))) OR (fsm_output(10));
  mux_2385_nl <= MUX_s_1_2_2(or_tmp_2405, or_tmp_2407, fsm_output(9));
  mux_tmp_2386 <= MUX_s_1_2_2(mux_tmp_2377, mux_2385_nl, fsm_output(6));
  mux_2387_nl <= MUX_s_1_2_2(or_tmp_2393, or_tmp_2394, fsm_output(8));
  mux_2388_nl <= MUX_s_1_2_2(mux_2387_nl, or_tmp_2407, fsm_output(9));
  mux_tmp_2389 <= MUX_s_1_2_2(mux_tmp_2377, mux_2388_nl, fsm_output(6));
  or_2475_nl <= (NOT (fsm_output(1))) OR (NOT (fsm_output(6))) OR (fsm_output(10));
  or_2474_nl <= (fsm_output(1)) OR not_tmp_49;
  mux_tmp_2424 <= MUX_s_1_2_2(or_2475_nl, or_2474_nl, fsm_output(3));
  nand_183_cse <= NOT((fsm_output(1)) AND (fsm_output(6)) AND (fsm_output(10)));
  or_2488_nl <= (NOT (fsm_output(9))) OR (NOT (fsm_output(2))) OR (fsm_output(7))
      OR (NOT (fsm_output(3))) OR (fsm_output(1)) OR (fsm_output(6)) OR (fsm_output(10));
  or_2487_nl <= (fsm_output(9)) OR (NOT (fsm_output(2))) OR (fsm_output(7)) OR (NOT
      (fsm_output(3))) OR (NOT (fsm_output(1))) OR (fsm_output(6)) OR (NOT (fsm_output(10)));
  mux_2430_nl <= MUX_s_1_2_2(or_2488_nl, or_2487_nl, fsm_output(0));
  nor_741_nl <= NOT((fsm_output(5)) OR mux_2430_nl);
  or_2484_nl <= (fsm_output(3)) OR (NOT (fsm_output(1))) OR (fsm_output(6)) OR (NOT
      (fsm_output(10)));
  nand_182_nl <= NOT((fsm_output(3)) AND (fsm_output(1)) AND (fsm_output(6)) AND
      (NOT (fsm_output(10))));
  mux_2427_nl <= MUX_s_1_2_2(or_2484_nl, nand_182_nl, fsm_output(7));
  nor_742_nl <= NOT((NOT (fsm_output(9))) OR (fsm_output(2)) OR mux_2427_nl);
  nor_743_nl <= NOT((fsm_output(9)) OR (NOT (fsm_output(2))) OR (NOT (fsm_output(7)))
      OR mux_tmp_2424);
  mux_2428_nl <= MUX_s_1_2_2(nor_742_nl, nor_743_nl, fsm_output(0));
  or_2479_nl <= (fsm_output(7)) OR (fsm_output(3)) OR (fsm_output(1)) OR (NOT (fsm_output(6)))
      OR (fsm_output(10));
  or_2478_nl <= (fsm_output(7)) OR (fsm_output(3)) OR nand_183_cse;
  mux_2425_nl <= MUX_s_1_2_2(or_2479_nl, or_2478_nl, fsm_output(2));
  nor_744_nl <= NOT((fsm_output(9)) OR mux_2425_nl);
  nor_745_nl <= NOT((NOT (fsm_output(9))) OR (fsm_output(2)) OR (fsm_output(7)) OR
      mux_tmp_2424);
  mux_2426_nl <= MUX_s_1_2_2(nor_744_nl, nor_745_nl, fsm_output(0));
  mux_2429_nl <= MUX_s_1_2_2(mux_2428_nl, mux_2426_nl, fsm_output(5));
  mux_2431_nl <= MUX_s_1_2_2(nor_741_nl, mux_2429_nl, fsm_output(4));
  nor_746_nl <= NOT((fsm_output(9)) OR (NOT (fsm_output(2))) OR (fsm_output(7)) OR
      (fsm_output(3)) OR (fsm_output(1)) OR not_tmp_49);
  nor_747_nl <= NOT((NOT (fsm_output(9))) OR (fsm_output(2)) OR (fsm_output(7)) OR
      (fsm_output(3)) OR (fsm_output(1)) OR (NOT (fsm_output(6))) OR (fsm_output(10)));
  mux_2421_nl <= MUX_s_1_2_2(nor_746_nl, nor_747_nl, fsm_output(0));
  nor_748_nl <= NOT((NOT (fsm_output(9))) OR (fsm_output(2)) OR (NOT (fsm_output(7)))
      OR (NOT (fsm_output(3))) OR (fsm_output(1)) OR (fsm_output(6)) OR (fsm_output(10)));
  nand_388_nl <= NOT((fsm_output(7)) AND (fsm_output(3)) AND (fsm_output(1)) AND
      (NOT (fsm_output(6))) AND (fsm_output(10)));
  or_2465_nl <= (NOT (fsm_output(7))) OR (fsm_output(3)) OR (fsm_output(1)) OR (fsm_output(6))
      OR (fsm_output(10));
  mux_2419_nl <= MUX_s_1_2_2(nand_388_nl, or_2465_nl, fsm_output(2));
  nor_749_nl <= NOT((fsm_output(9)) OR mux_2419_nl);
  mux_2420_nl <= MUX_s_1_2_2(nor_748_nl, nor_749_nl, fsm_output(0));
  mux_2422_nl <= MUX_s_1_2_2(mux_2421_nl, mux_2420_nl, fsm_output(5));
  nor_750_nl <= NOT((NOT (fsm_output(5))) OR (fsm_output(0)) OR (fsm_output(9)) OR
      (NOT (fsm_output(2))) OR (fsm_output(7)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(1)))
      OR (fsm_output(6)) OR (fsm_output(10)));
  mux_2423_nl <= MUX_s_1_2_2(mux_2422_nl, nor_750_nl, fsm_output(4));
  not_tmp_441 <= MUX_s_1_2_2(mux_2431_nl, mux_2423_nl, fsm_output(8));
  or_tmp_2436 <= NOT((fsm_output(3)) AND (fsm_output(8)) AND (fsm_output(6)) AND
      (NOT (fsm_output(10))));
  or_2512_nl <= (fsm_output(3)) OR (fsm_output(8)) OR (fsm_output(6)) OR (NOT (fsm_output(10)));
  mux_2442_nl <= MUX_s_1_2_2(or_tmp_2436, or_2512_nl, fsm_output(7));
  nor_729_nl <= NOT((fsm_output(2)) OR (NOT (fsm_output(5))) OR mux_2442_nl);
  nor_730_nl <= NOT((NOT (fsm_output(2))) OR (fsm_output(5)) OR (fsm_output(7)) OR
      (fsm_output(3)) OR (NOT (fsm_output(8))) OR (fsm_output(6)) OR (fsm_output(10)));
  mux_2443_nl <= MUX_s_1_2_2(nor_729_nl, nor_730_nl, fsm_output(9));
  nor_1628_nl <= NOT((NOT (fsm_output(2))) OR (NOT (fsm_output(5))) OR (NOT (fsm_output(9)))
      OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (fsm_output(8)) OR (fsm_output(7))
      OR (NOT (fsm_output(10))));
  mux_2444_nl <= MUX_s_1_2_2(mux_2443_nl, nor_1628_nl, fsm_output(4));
  nor_732_nl <= NOT((fsm_output(9)) OR (NOT (fsm_output(2))) OR (NOT (fsm_output(5)))
      OR (fsm_output(7)) OR (NOT((fsm_output(3)) AND (fsm_output(8)) AND (fsm_output(6))
      AND (fsm_output(10)))));
  nor_733_nl <= NOT((fsm_output(2)) OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR
      (NOT (fsm_output(3))) OR (fsm_output(8)) OR (fsm_output(6)) OR (fsm_output(10)));
  nor_734_nl <= NOT((fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(3)) OR
      (NOT (fsm_output(8))) OR (NOT (fsm_output(6))) OR (fsm_output(10)));
  nor_735_nl <= NOT((NOT (fsm_output(5))) OR (fsm_output(7)) OR (fsm_output(3)) OR
      (fsm_output(8)) OR (fsm_output(6)) OR (fsm_output(10)));
  mux_2439_nl <= MUX_s_1_2_2(nor_734_nl, nor_735_nl, fsm_output(2));
  mux_2440_nl <= MUX_s_1_2_2(nor_733_nl, mux_2439_nl, fsm_output(9));
  mux_2441_nl <= MUX_s_1_2_2(nor_732_nl, mux_2440_nl, fsm_output(4));
  mux_2445_nl <= MUX_s_1_2_2(mux_2444_nl, mux_2441_nl, fsm_output(1));
  nor_736_nl <= NOT((fsm_output(9)) OR (fsm_output(2)) OR (fsm_output(5)) OR (fsm_output(7))
      OR (fsm_output(3)) OR (NOT (fsm_output(8))) OR (fsm_output(6)) OR (fsm_output(10)));
  nor_737_nl <= NOT((NOT (fsm_output(5))) OR (fsm_output(7)) OR (NOT (fsm_output(3)))
      OR (fsm_output(8)) OR (fsm_output(6)) OR (NOT (fsm_output(10))));
  nor_738_nl <= NOT((fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(3)) OR
      nand_142_cse);
  mux_2435_nl <= MUX_s_1_2_2(nor_737_nl, nor_738_nl, fsm_output(2));
  nor_739_nl <= NOT((NOT (fsm_output(2))) OR (fsm_output(5)) OR (NOT (fsm_output(7)))
      OR (NOT (fsm_output(3))) OR (fsm_output(8)) OR (fsm_output(6)) OR (fsm_output(10)));
  mux_2436_nl <= MUX_s_1_2_2(mux_2435_nl, nor_739_nl, fsm_output(9));
  mux_2437_nl <= MUX_s_1_2_2(nor_736_nl, mux_2436_nl, fsm_output(4));
  or_2494_nl <= (fsm_output(3)) OR (NOT (fsm_output(8))) OR (fsm_output(6)) OR (NOT
      (fsm_output(10)));
  mux_2433_nl <= MUX_s_1_2_2(or_2494_nl, or_tmp_2436, fsm_output(7));
  or_2495_nl <= (NOT (fsm_output(2))) OR (fsm_output(5)) OR mux_2433_nl;
  or_2490_nl <= (fsm_output(2)) OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (NOT
      (fsm_output(3))) OR (NOT (fsm_output(8))) OR (NOT (fsm_output(6))) OR (fsm_output(10));
  mux_2434_nl <= MUX_s_1_2_2(or_2495_nl, or_2490_nl, fsm_output(9));
  nor_740_nl <= NOT((fsm_output(4)) OR mux_2434_nl);
  mux_2438_nl <= MUX_s_1_2_2(mux_2437_nl, nor_740_nl, fsm_output(1));
  not_tmp_446 <= MUX_s_1_2_2(mux_2445_nl, mux_2438_nl, fsm_output(0));
  mux_2447_nl <= MUX_s_1_2_2((fsm_output(3)), (NOT (fsm_output(3))), or_2368_cse);
  nor_1612_nl <= NOT(nor_758_cse OR (fsm_output(3)));
  mux_2448_nl <= MUX_s_1_2_2(mux_2447_nl, nor_1612_nl, fsm_output(0));
  and_dcpl_241 <= mux_2448_nl AND nor_1580_cse AND and_dcpl_191 AND (NOT (fsm_output(4)))
      AND nor_609_cse;
  and_dcpl_245 <= NOT((fsm_output(2)) OR (fsm_output(7)));
  nor_726_nl <= NOT(CONV_SL_1_1(fsm_output(5 DOWNTO 3)/=STD_LOGIC_VECTOR'("110")));
  nor_727_nl <= NOT(CONV_SL_1_1(fsm_output(5 DOWNTO 3)/=STD_LOGIC_VECTOR'("001")));
  mux_2453_nl <= MUX_s_1_2_2(nor_726_nl, nor_727_nl, fsm_output(0));
  and_dcpl_247 <= mux_2453_nl AND and_dcpl_245 AND and_dcpl_191 AND (NOT (fsm_output(1)))
      AND nor_609_cse;
  nor_tmp_324 <= (fsm_output(5)) AND (fsm_output(10));
  nand_386_cse <= NOT((NOT(or_3388_cse AND (fsm_output(2)))) AND nor_tmp_324);
  or_2528_cse <= nor_758_cse OR (fsm_output(5)) OR (fsm_output(10));
  or_tmp_2474 <= (fsm_output(5)) OR (fsm_output(10));
  or_2534_cse <= and_529_cse OR (fsm_output(5)) OR (NOT (fsm_output(10)));
  mux_2465_cse <= MUX_s_1_2_2((NOT (fsm_output(5))), or_tmp_2393, fsm_output(9));
  or_2540_cse <= (NOT (fsm_output(2))) OR (fsm_output(5)) OR (fsm_output(10));
  or_2541_cse <= (fsm_output(2)) OR (NOT nor_tmp_324);
  nand_173_cse <= NOT(nand_196_cse AND nor_tmp_324);
  mux_2486_cse <= MUX_s_1_2_2((NOT (fsm_output(10))), (fsm_output(10)), fsm_output(5));
  mux_2494_cse <= MUX_s_1_2_2(or_tmp_2474, (fsm_output(5)), fsm_output(2));
  mux_2515_cse <= MUX_s_1_2_2((fsm_output(5)), nor_tmp_324, fsm_output(2));
  mux_2516_cse <= MUX_s_1_2_2(or_tmp_2474, nor_tmp_324, fsm_output(2));
  mux_tmp_2640 <= MUX_s_1_2_2(nor_609_cse, and_757_cse, fsm_output(7));
  nor_694_cse <= NOT((fsm_output(7)) OR (fsm_output(9)) OR (fsm_output(10)));
  and_465_cse <= (fsm_output(5)) AND (fsm_output(7)) AND (fsm_output(9)) AND (fsm_output(10));
  mux_tmp_2659 <= MUX_s_1_2_2(nor_694_cse, and_756_cse, fsm_output(5));
  and_dcpl_256 <= and_dcpl_108 AND and_dcpl_55 AND nor_609_cse;
  mux_tmp_2669 <= MUX_s_1_2_2((NOT (fsm_output(6))), or_352_cse, fsm_output(9));
  mux_tmp_2672 <= MUX_s_1_2_2(and_757_cse, mux_tmp_2669, fsm_output(7));
  mux_tmp_2675 <= MUX_s_1_2_2((fsm_output(6)), or_tmp_167, fsm_output(9));
  not_tmp_500 <= MUX_s_1_2_2(or_tmp_167, (NOT mux_554_cse), fsm_output(9));
  mux_2681_nl <= MUX_s_1_2_2(mux_554_cse, nor_tmp_48, fsm_output(9));
  mux_tmp_2682 <= MUX_s_1_2_2((NOT mux_2681_nl), mux_tmp_2675, fsm_output(7));
  mux_tmp_2690 <= MUX_s_1_2_2(mux_tmp_2675, and_757_cse, fsm_output(7));
  mux_tmp_2691 <= MUX_s_1_2_2(mux_tmp_2675, and_672_cse, fsm_output(7));
  mux_tmp_2693 <= MUX_s_1_2_2(nor_tmp_48, or_tmp_167, fsm_output(9));
  or_tmp_2603 <= (fsm_output(6)) OR (NOT (fsm_output(10)));
  mux_2698_itm <= MUX_s_1_2_2(or_tmp_2603, (fsm_output(6)), fsm_output(9));
  or_tmp_2604 <= (fsm_output(9)) OR (NOT mux_554_cse);
  mux_tmp_2700 <= MUX_s_1_2_2((NOT mux_2698_itm), or_tmp_2604, fsm_output(7));
  mux_tmp_2702 <= MUX_s_1_2_2((NOT nor_tmp_48), or_352_cse, fsm_output(9));
  mux_tmp_2703 <= MUX_s_1_2_2((NOT mux_2698_itm), mux_tmp_2702, fsm_output(7));
  mux_tmp_2706 <= MUX_s_1_2_2((NOT mux_2698_itm), mux_tmp_2669, fsm_output(7));
  mux_2708_nl <= MUX_s_1_2_2(or_tmp_2603, or_tmp_167, fsm_output(9));
  mux_tmp_2709 <= MUX_s_1_2_2((NOT mux_2708_nl), mux_tmp_2669, fsm_output(7));
  mux_tmp_2715 <= MUX_s_1_2_2(and_672_cse, mux_tmp_2669, fsm_output(7));
  nor_1575_nl <= NOT((fsm_output(9)) OR (fsm_output(6)) OR (fsm_output(10)));
  mux_tmp_2736 <= MUX_s_1_2_2(nor_1575_nl, mux_tmp_2669, fsm_output(7));
  and_dcpl_257 <= and_dcpl_108 AND and_dcpl_112;
  and_dcpl_260 <= and_dcpl_92 AND and_dcpl_136;
  and_dcpl_262 <= and_dcpl_135 AND (fsm_output(6));
  and_dcpl_270 <= and_dcpl_147 AND and_dcpl_44;
  and_dcpl_278 <= and_dcpl_6 AND and_dcpl_90;
  and_dcpl_280 <= and_dcpl_19 AND (fsm_output(0));
  or_2678_nl <= (NOT (fsm_output(1))) OR (NOT (fsm_output(2))) OR (NOT (fsm_output(6)))
      OR (NOT (fsm_output(8))) OR (fsm_output(4)) OR (fsm_output(10));
  or_2677_nl <= (fsm_output(1)) OR (NOT (fsm_output(2))) OR (fsm_output(6)) OR (fsm_output(8))
      OR (NOT (fsm_output(4))) OR (fsm_output(10));
  mux_tmp_2745 <= MUX_s_1_2_2(or_2678_nl, or_2677_nl, fsm_output(9));
  or_2694_nl <= (fsm_output(2)) OR (fsm_output(6)) OR (NOT (fsm_output(8))) OR (fsm_output(4))
      OR (fsm_output(10));
  or_2693_nl <= (NOT (fsm_output(2))) OR (fsm_output(6)) OR (NOT (fsm_output(8)))
      OR (fsm_output(4)) OR (NOT (fsm_output(10)));
  mux_2754_nl <= MUX_s_1_2_2(or_2694_nl, or_2693_nl, fsm_output(1));
  or_2695_nl <= (fsm_output(9)) OR mux_2754_nl;
  mux_2755_nl <= MUX_s_1_2_2(or_2695_nl, or_70_cse, fsm_output(0));
  or_2696_nl <= (fsm_output(3)) OR mux_2755_nl;
  or_2690_nl <= (fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(2)) OR (fsm_output(6))
      OR (fsm_output(8)) OR (NOT (fsm_output(4))) OR (fsm_output(10));
  mux_2752_nl <= MUX_s_1_2_2(or_2690_nl, mux_tmp_2745, fsm_output(0));
  or_2689_nl <= (fsm_output(1)) OR (fsm_output(2)) OR (fsm_output(6)) OR (fsm_output(8))
      OR not_tmp_39;
  or_2687_nl <= (NOT (fsm_output(1))) OR (fsm_output(2)) OR (NOT (fsm_output(6)))
      OR (NOT (fsm_output(8))) OR (fsm_output(4)) OR (fsm_output(10));
  mux_2750_nl <= MUX_s_1_2_2(or_2689_nl, or_2687_nl, fsm_output(9));
  or_2686_nl <= (fsm_output(1)) OR (NOT (fsm_output(2))) OR (NOT (fsm_output(6)))
      OR (NOT (fsm_output(8))) OR (fsm_output(4)) OR (NOT (fsm_output(10)));
  or_2684_nl <= (NOT (fsm_output(1))) OR (fsm_output(2)) OR (fsm_output(6)) OR (fsm_output(8))
      OR not_tmp_39;
  mux_2749_nl <= MUX_s_1_2_2(or_2686_nl, or_2684_nl, fsm_output(9));
  mux_2751_nl <= MUX_s_1_2_2(mux_2750_nl, mux_2749_nl, fsm_output(0));
  mux_2753_nl <= MUX_s_1_2_2(mux_2752_nl, mux_2751_nl, fsm_output(3));
  mux_2756_nl <= MUX_s_1_2_2(or_2696_nl, mux_2753_nl, fsm_output(5));
  or_2681_nl <= (fsm_output(9)) OR (fsm_output(1)) OR (NOT((fsm_output(2)) AND (fsm_output(6))
      AND (fsm_output(8)) AND (fsm_output(4)) AND (fsm_output(10))));
  mux_2747_nl <= MUX_s_1_2_2(or_2681_nl, or_56_cse, fsm_output(0));
  or_2675_nl <= (fsm_output(2)) OR (fsm_output(6)) OR (fsm_output(8)) OR (NOT (fsm_output(4)))
      OR (fsm_output(10));
  or_2674_nl <= (NOT (fsm_output(2))) OR (fsm_output(6)) OR (fsm_output(8)) OR not_tmp_39;
  mux_2744_nl <= MUX_s_1_2_2(or_2675_nl, or_2674_nl, fsm_output(1));
  or_2676_nl <= (fsm_output(9)) OR mux_2744_nl;
  mux_2746_nl <= MUX_s_1_2_2(mux_tmp_2745, or_2676_nl, fsm_output(0));
  mux_2748_nl <= MUX_s_1_2_2(mux_2747_nl, mux_2746_nl, fsm_output(3));
  or_2682_nl <= (fsm_output(5)) OR mux_2748_nl;
  mux_2757_itm <= MUX_s_1_2_2(mux_2756_nl, or_2682_nl, fsm_output(7));
  or_2705_nl <= (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(6)) OR (fsm_output(10));
  or_2704_nl <= (fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(6)) OR (NOT
      (fsm_output(10)));
  mux_tmp_2760 <= MUX_s_1_2_2(or_2705_nl, or_2704_nl, fsm_output(2));
  or_tmp_2651 <= (fsm_output(2)) OR (fsm_output(9)) OR (NOT (fsm_output(1))) OR (NOT
      (fsm_output(6))) OR (fsm_output(10));
  or_tmp_2682 <= CONV_SL_1_1(fsm_output(10 DOWNTO 7)/=STD_LOGIC_VECTOR'("0110"));
  or_tmp_2683 <= NOT(CONV_SL_1_1(fsm_output(10 DOWNTO 7)=STD_LOGIC_VECTOR'("0111")));
  or_tmp_2690 <= (fsm_output(7)) OR (fsm_output(9)) OR nand_138_cse;
  or_tmp_2693 <= CONV_SL_1_1(fsm_output(10 DOWNTO 7)/=STD_LOGIC_VECTOR'("0010"));
  or_tmp_2696 <= CONV_SL_1_1(fsm_output(10 DOWNTO 7)/=STD_LOGIC_VECTOR'("0011"));
  or_tmp_2697 <= CONV_SL_1_1(fsm_output(10 DOWNTO 7)/=STD_LOGIC_VECTOR'("0100"));
  mux_tmp_2796 <= MUX_s_1_2_2(or_3008_cse, or_2998_cse, fsm_output(7));
  or_tmp_2701 <= CONV_SL_1_1(fsm_output(10 DOWNTO 7)/=STD_LOGIC_VECTOR'("0001"));
  or_tmp_2703 <= CONV_SL_1_1(fsm_output(10 DOWNTO 7)/=STD_LOGIC_VECTOR'("1000"));
  or_tmp_2704 <= CONV_SL_1_1(fsm_output(10 DOWNTO 7)/=STD_LOGIC_VECTOR'("0101"));
  or_tmp_2706 <= CONV_SL_1_1(fsm_output(10 DOWNTO 7)/=STD_LOGIC_VECTOR'("1100"));
  or_tmp_2709 <= CONV_SL_1_1(fsm_output(10 DOWNTO 7)/=STD_LOGIC_VECTOR'("1001"));
  or_tmp_2714 <= (NOT (fsm_output(7))) OR (fsm_output(9)) OR nand_138_cse;
  or_2785_nl <= (fsm_output(4)) OR (fsm_output(3)) OR (fsm_output(7)) OR (NOT (fsm_output(9)))
      OR (NOT (fsm_output(8))) OR (fsm_output(10));
  or_2784_nl <= (NOT((fsm_output(3)) AND (fsm_output(6)) AND (fsm_output(7)) AND
      (NOT (fsm_output(9))))) OR nand_138_cse;
  mux_2834_nl <= MUX_s_1_2_2(or_tmp_2704, or_tmp_2709, fsm_output(6));
  mux_2832_nl <= MUX_s_1_2_2(or_2387_cse, or_2991_cse, fsm_output(7));
  mux_2833_nl <= MUX_s_1_2_2(mux_2832_nl, or_tmp_2706, fsm_output(6));
  mux_2835_nl <= MUX_s_1_2_2(mux_2834_nl, mux_2833_nl, fsm_output(3));
  mux_2836_nl <= MUX_s_1_2_2(or_2784_nl, mux_2835_nl, fsm_output(4));
  mux_2837_nl <= MUX_s_1_2_2(or_2785_nl, mux_2836_nl, fsm_output(5));
  nand_394_nl <= NOT(CONV_SL_1_1(fsm_output(10 DOWNTO 7)=STD_LOGIC_VECTOR'("1101")));
  mux_2829_nl <= MUX_s_1_2_2(nand_394_nl, or_tmp_2703, fsm_output(6));
  nand_65_nl <= NOT((fsm_output(3)) AND (NOT mux_2829_nl));
  mux_2827_nl <= MUX_s_1_2_2(or_tmp_2693, or_tmp_2682, fsm_output(6));
  mux_2828_nl <= MUX_s_1_2_2(mux_2827_nl, or_tmp_2709, fsm_output(3));
  mux_2830_nl <= MUX_s_1_2_2(nand_65_nl, mux_2828_nl, fsm_output(4));
  mux_2826_nl <= MUX_s_1_2_2(or_tmp_2696, or_tmp_2693, fsm_output(6));
  or_2780_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("00")) OR mux_2826_nl;
  mux_2831_nl <= MUX_s_1_2_2(mux_2830_nl, or_2780_nl, fsm_output(5));
  mux_2838_nl <= MUX_s_1_2_2(mux_2837_nl, mux_2831_nl, fsm_output(2));
  or_2778_nl <= (NOT (fsm_output(4))) OR (NOT (fsm_output(3))) OR (fsm_output(6))
      OR (fsm_output(7)) OR (fsm_output(9)) OR nand_138_cse;
  mux_2821_nl <= MUX_s_1_2_2(or_tmp_2703, or_tmp_2696, fsm_output(6));
  mux_2820_nl <= MUX_s_1_2_2(or_tmp_2714, mux_tmp_2796, fsm_output(6));
  mux_2822_nl <= MUX_s_1_2_2(mux_2821_nl, mux_2820_nl, fsm_output(3));
  or_2776_nl <= (fsm_output(3)) OR (fsm_output(7)) OR (NOT (fsm_output(9))) OR (fsm_output(8))
      OR (fsm_output(10));
  mux_2823_nl <= MUX_s_1_2_2(mux_2822_nl, or_2776_nl, fsm_output(4));
  mux_2824_nl <= MUX_s_1_2_2(or_2778_nl, mux_2823_nl, fsm_output(5));
  or_2775_nl <= CONV_SL_1_1(fsm_output(10 DOWNTO 6)/=STD_LOGIC_VECTOR'("01010"));
  mux_2816_nl <= MUX_s_1_2_2(or_tmp_2703, or_tmp_2683, fsm_output(6));
  mux_2817_nl <= MUX_s_1_2_2(or_2775_nl, mux_2816_nl, fsm_output(3));
  or_2774_nl <= (fsm_output(3)) OR (NOT (fsm_output(7))) OR (fsm_output(9)) OR (fsm_output(8))
      OR (fsm_output(10));
  mux_2818_nl <= MUX_s_1_2_2(mux_2817_nl, or_2774_nl, fsm_output(4));
  mux_2815_nl <= MUX_s_1_2_2(or_tmp_2714, or_tmp_2682, fsm_output(6));
  nand_64_nl <= NOT(CONV_SL_1_1(fsm_output(4 DOWNTO 3)=STD_LOGIC_VECTOR'("11")) AND
      (NOT mux_2815_nl));
  mux_2819_nl <= MUX_s_1_2_2(mux_2818_nl, nand_64_nl, fsm_output(5));
  mux_2825_nl <= MUX_s_1_2_2(mux_2824_nl, mux_2819_nl, fsm_output(2));
  mux_2839_nl <= MUX_s_1_2_2(mux_2838_nl, mux_2825_nl, fsm_output(1));
  or_2770_nl <= (fsm_output(6)) OR (NOT (fsm_output(7))) OR (fsm_output(9)) OR nand_138_cse;
  mux_2810_nl <= MUX_s_1_2_2(or_tmp_2709, or_tmp_2697, fsm_output(6));
  mux_2811_nl <= MUX_s_1_2_2(or_2770_nl, mux_2810_nl, fsm_output(3));
  mux_2807_nl <= MUX_s_1_2_2(or_2991_cse, or_3008_cse, fsm_output(7));
  mux_2808_nl <= MUX_s_1_2_2(or_tmp_2706, mux_2807_nl, fsm_output(6));
  mux_2809_nl <= MUX_s_1_2_2(mux_2808_nl, or_tmp_2704, fsm_output(3));
  mux_2812_nl <= MUX_s_1_2_2(mux_2811_nl, mux_2809_nl, fsm_output(4));
  or_2771_nl <= (fsm_output(5)) OR mux_2812_nl;
  mux_2804_nl <= MUX_s_1_2_2(or_tmp_2706, or_tmp_2683, fsm_output(6));
  mux_2803_nl <= MUX_s_1_2_2(or_tmp_2701, or_tmp_2704, fsm_output(6));
  mux_2805_nl <= MUX_s_1_2_2(mux_2804_nl, mux_2803_nl, fsm_output(3));
  mux_2801_nl <= MUX_s_1_2_2(or_tmp_2693, or_tmp_2701, fsm_output(6));
  mux_2802_nl <= MUX_s_1_2_2(or_tmp_2703, mux_2801_nl, fsm_output(3));
  mux_2806_nl <= MUX_s_1_2_2(mux_2805_nl, mux_2802_nl, fsm_output(4));
  nand_63_nl <= NOT((fsm_output(5)) AND (NOT mux_2806_nl));
  mux_2813_nl <= MUX_s_1_2_2(or_2771_nl, nand_63_nl, fsm_output(2));
  mux_2797_nl <= MUX_s_1_2_2(mux_tmp_2796, or_tmp_2690, fsm_output(6));
  mux_2795_nl <= MUX_s_1_2_2(or_tmp_2697, or_tmp_2696, fsm_output(6));
  mux_2798_nl <= MUX_s_1_2_2(mux_2797_nl, mux_2795_nl, fsm_output(3));
  or_2759_nl <= (fsm_output(4)) OR mux_2798_nl;
  or_2754_nl <= CONV_SL_1_1(fsm_output(10 DOWNTO 6)/=STD_LOGIC_VECTOR'("10010"));
  mux_2793_nl <= MUX_s_1_2_2(or_tmp_2683, or_tmp_2693, fsm_output(6));
  mux_2794_nl <= MUX_s_1_2_2(or_2754_nl, mux_2793_nl, fsm_output(3));
  nand_62_nl <= NOT((fsm_output(4)) AND (NOT mux_2794_nl));
  mux_2799_nl <= MUX_s_1_2_2(or_2759_nl, nand_62_nl, fsm_output(5));
  or_2751_nl <= (NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(7))
      OR (NOT (fsm_output(9))) OR (fsm_output(8)) OR (NOT (fsm_output(10)));
  mux_2789_nl <= MUX_s_1_2_2(or_tmp_2682, or_tmp_2690, fsm_output(6));
  mux_2788_nl <= MUX_s_1_2_2(or_2407_cse, or_2387_cse, fsm_output(7));
  or_2747_nl <= (fsm_output(6)) OR mux_2788_nl;
  mux_2790_nl <= MUX_s_1_2_2(mux_2789_nl, or_2747_nl, fsm_output(3));
  mux_2791_nl <= MUX_s_1_2_2(or_2751_nl, mux_2790_nl, fsm_output(4));
  mux_2786_nl <= MUX_s_1_2_2(or_tmp_2683, or_tmp_2682, fsm_output(6));
  or_2740_nl <= CONV_SL_1_1(fsm_output(10 DOWNTO 6)/=STD_LOGIC_VECTOR'("00001"));
  mux_2787_nl <= MUX_s_1_2_2(mux_2786_nl, or_2740_nl, fsm_output(3));
  or_2743_nl <= (fsm_output(4)) OR mux_2787_nl;
  mux_2792_nl <= MUX_s_1_2_2(mux_2791_nl, or_2743_nl, fsm_output(5));
  mux_2800_nl <= MUX_s_1_2_2(mux_2799_nl, mux_2792_nl, fsm_output(2));
  mux_2814_nl <= MUX_s_1_2_2(mux_2813_nl, mux_2800_nl, fsm_output(1));
  mux_2840_itm <= MUX_s_1_2_2(mux_2839_nl, mux_2814_nl, fsm_output(0));
  mux_tmp_2841 <= MUX_s_1_2_2((NOT or_tmp_2281), (fsm_output(10)), fsm_output(9));
  or_tmp_2729 <= (fsm_output(9)) OR (fsm_output(7)) OR (NOT (fsm_output(10)));
  or_tmp_2731 <= (NOT((NOT (fsm_output(9))) OR (fsm_output(7)))) OR (fsm_output(10));
  mux_tmp_2843 <= MUX_s_1_2_2(or_tmp_2281, or_tmp_2276, fsm_output(9));
  mux_tmp_2844 <= MUX_s_1_2_2(mux_tmp_2843, or_tmp_2731, fsm_output(6));
  or_tmp_2734 <= (fsm_output(6)) OR mux_tmp_2159;
  mux_tmp_2848 <= MUX_s_1_2_2((NOT and_395_cse), or_tmp_2280, fsm_output(9));
  mux_tmp_2850 <= MUX_s_1_2_2(mux_2171_cse, mux_tmp_2848, fsm_output(6));
  or_tmp_2736 <= (NOT (fsm_output(9))) OR (fsm_output(7)) OR (NOT (fsm_output(10)));
  mux_tmp_2851 <= MUX_s_1_2_2((NOT (fsm_output(7))), (fsm_output(10)), fsm_output(9));
  mux_tmp_2856 <= MUX_s_1_2_2((fsm_output(7)), or_tmp_2281, fsm_output(9));
  mux_2858_nl <= MUX_s_1_2_2((fsm_output(10)), (NOT and_395_cse), fsm_output(9));
  nand_tmp_67 <= NOT((fsm_output(6)) AND mux_2858_nl);
  mux_tmp_2862 <= MUX_s_1_2_2(or_tmp_2276, mux_tmp_2159, fsm_output(6));
  mux_tmp_2863 <= MUX_s_1_2_2((NOT or_tmp_2276), or_tmp_2280, fsm_output(9));
  or_tmp_2739 <= (fsm_output(9)) OR (NOT (fsm_output(7))) OR (fsm_output(10));
  mux_tmp_2867 <= MUX_s_1_2_2(or_tmp_2739, mux_2203_cse, fsm_output(6));
  or_tmp_2740 <= CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"));
  mux_2875_nl <= MUX_s_1_2_2((NOT or_tmp_2276), (fsm_output(10)), fsm_output(9));
  mux_tmp_2876 <= MUX_s_1_2_2(or_tmp_2736, mux_2875_nl, fsm_output(6));
  or_2800_nl <= (fsm_output(6)) OR mux_tmp_2863;
  mux_tmp_2878 <= MUX_s_1_2_2(or_tmp_2734, or_2800_nl, fsm_output(0));
  mux_tmp_2879 <= MUX_s_1_2_2(mux_2203_cse, or_tmp_2280, fsm_output(6));
  or_tmp_2742 <= (fsm_output(9)) OR (NOT (fsm_output(7)));
  mux_tmp_2880 <= MUX_s_1_2_2(mux_2203_cse, or_tmp_2742, fsm_output(6));
  mux_tmp_2886 <= MUX_s_1_2_2(mux_2171_cse, or_tmp_2742, fsm_output(6));
  mux_tmp_2888 <= MUX_s_1_2_2(mux_2171_cse, mux_tmp_2159, fsm_output(6));
  mux_tmp_2890 <= MUX_s_1_2_2(or_tmp_2280, or_tmp_2281, fsm_output(6));
  or_tmp_2743 <= (fsm_output(6)) OR mux_tmp_2841;
  nand_tmp_68 <= NOT((fsm_output(6)) AND (NOT mux_2203_cse));
  mux_tmp_2895 <= MUX_s_1_2_2((NOT (fsm_output(10))), (fsm_output(7)), fsm_output(9));
  or_tmp_2745 <= (fsm_output(6)) OR (fsm_output(9)) OR (NOT (fsm_output(7)));
  or_tmp_2746 <= (NOT (fsm_output(9))) OR (NOT (fsm_output(7))) OR (fsm_output(10));
  mux_2901_nl <= MUX_s_1_2_2(or_tmp_2276, (NOT and_395_cse), fsm_output(9));
  nand_tmp_69 <= NOT((fsm_output(6)) AND mux_2901_nl);
  mux_tmp_2906 <= MUX_s_1_2_2(mux_tmp_2843, mux_tmp_2159, fsm_output(6));
  mux_2909_nl <= MUX_s_1_2_2((NOT or_tmp_2280), (fsm_output(10)), fsm_output(9));
  mux_tmp_2910 <= MUX_s_1_2_2(mux_2909_nl, or_tmp_2739, fsm_output(6));
  nand_tmp_70 <= NOT((fsm_output(6)) AND (NOT mux_2171_cse));
  mux_tmp_2912 <= MUX_s_1_2_2(or_tmp_2276, (fsm_output(7)), fsm_output(9));
  nand_tmp_71 <= NOT((fsm_output(6)) AND (NOT mux_tmp_2912));
  mux_tmp_2916 <= MUX_s_1_2_2(or_tmp_2281, mux_tmp_2851, fsm_output(6));
  mux_tmp_2920 <= MUX_s_1_2_2(mux_2203_cse, mux_tmp_2848, fsm_output(6));
  or_tmp_2749 <= (fsm_output(9)) OR (NOT and_395_cse);
  or_tmp_2774 <= (NOT (fsm_output(1))) OR (NOT (fsm_output(8))) OR (fsm_output(6))
      OR (fsm_output(10));
  or_2835_cse <= (NOT (fsm_output(1))) OR (fsm_output(8)) OR not_tmp_49;
  mux_tmp_2996 <= MUX_s_1_2_2(or_2835_cse, or_tmp_2774, fsm_output(3));
  nor_667_cse <= NOT((NOT (fsm_output(7))) OR (fsm_output(3)) OR (fsm_output(1))
      OR (NOT (fsm_output(8))) OR (NOT (fsm_output(6))) OR (fsm_output(10)));
  or_2840_nl <= (fsm_output(1)) OR (NOT (fsm_output(8))) OR (fsm_output(6)) OR (NOT
      (fsm_output(10)));
  mux_2998_cse <= MUX_s_1_2_2(or_tmp_2774, or_2840_nl, fsm_output(3));
  nor_661_nl <= NOT((fsm_output(0)) OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR
      (fsm_output(3)) OR (fsm_output(1)) OR (fsm_output(8)) OR (NOT (fsm_output(6)))
      OR (fsm_output(10)));
  or_2842_nl <= (fsm_output(3)) OR (NOT (fsm_output(1))) OR (fsm_output(8)) OR (NOT
      (fsm_output(6))) OR (fsm_output(10));
  mux_2999_nl <= MUX_s_1_2_2(or_2842_nl, mux_tmp_2996, fsm_output(7));
  nor_662_nl <= NOT((fsm_output(5)) OR mux_2999_nl);
  nor_663_nl <= NOT((NOT (fsm_output(5))) OR (fsm_output(7)) OR mux_2998_cse);
  mux_3000_nl <= MUX_s_1_2_2(nor_662_nl, nor_663_nl, fsm_output(0));
  mux_3001_nl <= MUX_s_1_2_2(nor_661_nl, mux_3000_nl, fsm_output(2));
  or_2836_nl <= (NOT (fsm_output(5))) OR (fsm_output(7)) OR mux_tmp_2996;
  or_2831_nl <= (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(3)) OR (NOT
      (fsm_output(1))) OR (fsm_output(8)) OR (NOT (fsm_output(6))) OR (fsm_output(10));
  mux_2997_nl <= MUX_s_1_2_2(or_2836_nl, or_2831_nl, fsm_output(0));
  nor_664_nl <= NOT((fsm_output(2)) OR mux_2997_nl);
  mux_3002_nl <= MUX_s_1_2_2(mux_3001_nl, nor_664_nl, fsm_output(9));
  and_445_nl <= (fsm_output(0)) AND (fsm_output(5)) AND (fsm_output(7)) AND (fsm_output(3))
      AND (fsm_output(1)) AND (fsm_output(8)) AND (fsm_output(6)) AND (fsm_output(10));
  nor_665_nl <= NOT((fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(3)) OR
      (fsm_output(1)) OR (NOT (fsm_output(8))) OR (fsm_output(6)) OR (NOT (fsm_output(10))));
  nor_666_nl <= NOT((fsm_output(7)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(1)))
      OR (fsm_output(8)) OR not_tmp_49);
  mux_2992_nl <= MUX_s_1_2_2(nor_666_nl, nor_667_cse, fsm_output(5));
  mux_2993_nl <= MUX_s_1_2_2(nor_665_nl, mux_2992_nl, fsm_output(0));
  mux_2994_nl <= MUX_s_1_2_2(and_445_nl, mux_2993_nl, fsm_output(2));
  and_446_nl <= (fsm_output(5)) AND (fsm_output(7)) AND (fsm_output(3)) AND (NOT
      (fsm_output(1))) AND (fsm_output(8)) AND (fsm_output(6)) AND (NOT (fsm_output(10)));
  nor_668_nl <= NOT((fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(3)) OR
      (fsm_output(1)) OR (NOT (fsm_output(8))) OR (fsm_output(6)) OR (fsm_output(10)));
  mux_2990_nl <= MUX_s_1_2_2(and_446_nl, nor_668_nl, fsm_output(0));
  nor_669_nl <= NOT((fsm_output(0)) OR (fsm_output(5)) OR (fsm_output(7)) OR (NOT
      (fsm_output(3))) OR (fsm_output(1)) OR (fsm_output(8)) OR (NOT (fsm_output(6)))
      OR (fsm_output(10)));
  mux_2991_nl <= MUX_s_1_2_2(mux_2990_nl, nor_669_nl, fsm_output(2));
  mux_2995_nl <= MUX_s_1_2_2(mux_2994_nl, mux_2991_nl, fsm_output(9));
  not_tmp_557 <= MUX_s_1_2_2(mux_3002_nl, mux_2995_nl, fsm_output(4));
  nor_tmp_405 <= (fsm_output(8)) AND (fsm_output(10));
  mux_3799_nl <= MUX_s_1_2_2(or_tmp_88, (NOT (fsm_output(8))), fsm_output(2));
  mux_tmp_3007 <= MUX_s_1_2_2(mux_3799_nl, or_tmp_88, fsm_output(9));
  mux_3006_nl <= MUX_s_1_2_2(or_tmp_88, (NOT (fsm_output(8))), fsm_output(2));
  or_2848_nl <= (NOT (fsm_output(2))) OR (NOT (fsm_output(8))) OR (fsm_output(10));
  mux_tmp_3008 <= MUX_s_1_2_2(mux_3006_nl, or_2848_nl, fsm_output(9));
  or_tmp_2791 <= nor_657_cse OR (NOT (fsm_output(8))) OR (fsm_output(10));
  mux_tmp_3014 <= MUX_s_1_2_2((fsm_output(8)), or_tmp_93, fsm_output(2));
  or_tmp_2795 <= (fsm_output(2)) OR (fsm_output(8)) OR (NOT (fsm_output(10)));
  or_tmp_2802 <= (fsm_output(9)) OR (fsm_output(2)) OR (NOT nor_tmp_405);
  or_tmp_2803 <= (fsm_output(2)) OR (NOT (fsm_output(8))) OR (fsm_output(10));
  or_2863_nl <= (fsm_output(2)) OR (NOT nor_tmp_405);
  mux_tmp_3024 <= MUX_s_1_2_2(or_2863_nl, or_tmp_2803, fsm_output(9));
  mux_3031_nl <= MUX_s_1_2_2((fsm_output(8)), nor_tmp_405, fsm_output(2));
  mux_tmp_3032 <= MUX_s_1_2_2((NOT mux_3031_nl), or_tmp_88, fsm_output(9));
  mux_tmp_3049 <= MUX_s_1_2_2(or_tmp_2791, mux_tmp_3008, fsm_output(0));
  or_tmp_2814 <= (fsm_output(2)) OR (fsm_output(8)) OR (fsm_output(10));
  nor_tmp_410 <= (fsm_output(1)) AND (fsm_output(4)) AND (fsm_output(3)) AND (fsm_output(10));
  and_dcpl_304 <= and_dcpl_108 AND and_dcpl_280 AND nor_609_cse;
  or_3025_nl <= (fsm_output(2)) OR (fsm_output(1)) OR (fsm_output(3)) OR (fsm_output(6))
      OR (fsm_output(7)) OR (fsm_output(8));
  mux_3321_nl <= MUX_s_1_2_2(or_3079_cse, or_3025_nl, and_407_cse);
  or_3367_nl <= (fsm_output(10)) OR mux_3321_nl;
  or_3023_nl <= and_524_cse OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000"));
  or_3022_nl <= (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(7)) OR (fsm_output(8));
  mux_3319_nl <= MUX_s_1_2_2(or_3023_nl, or_3022_nl, fsm_output(2));
  mux_3320_nl <= MUX_s_1_2_2(or_3079_cse, mux_3319_nl, and_407_cse);
  nand_149_nl <= NOT((fsm_output(10)) AND mux_3320_nl);
  not_tmp_619 <= MUX_s_1_2_2(or_3367_nl, nand_149_nl, fsm_output(9));
  mux_tmp_3329 <= MUX_s_1_2_2(nor_694_cse, and_757_cse, fsm_output(6));
  nor_tmp_457 <= CONV_SL_1_1(fsm_output(7 DOWNTO 6)=STD_LOGIC_VECTOR'("11"));
  mux_tmp_3341 <= MUX_s_1_2_2((NOT (fsm_output(7))), (fsm_output(7)), fsm_output(6));
  mux_3342_nl <= MUX_s_1_2_2(not_tmp_90, mux_tmp_3341, fsm_output(3));
  mux_tmp_3343 <= MUX_s_1_2_2(mux_3342_nl, nor_tmp_457, fsm_output(4));
  mux_tmp_3361 <= MUX_s_1_2_2(nor_tmp_4, (fsm_output(5)), fsm_output(2));
  or_tmp_2988 <= (NOT((fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(7)) OR (fsm_output(8))
      OR (fsm_output(9)))) OR (fsm_output(10));
  or_3061_nl <= CONV_SL_1_1(fsm_output(9 DOWNTO 6)/=STD_LOGIC_VECTOR'("0000"));
  mux_tmp_3378 <= MUX_s_1_2_2((NOT (fsm_output(10))), (fsm_output(10)), or_3061_nl);
  not_tmp_647 <= NOT((fsm_output(6)) OR (fsm_output(7)) OR (fsm_output(10)));
  or_3087_nl <= CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("00")) OR (NOT
      and_dcpl_209);
  or_12_nl <= (fsm_output(8)) OR (fsm_output(7)) OR (fsm_output(5));
  mux_tmp_3410 <= MUX_s_1_2_2(or_3087_nl, or_12_nl, fsm_output(6));
  mux_tmp_3414 <= MUX_s_1_2_2((NOT (fsm_output(3))), (fsm_output(3)), fsm_output(5));
  mux_tmp_3415 <= MUX_s_1_2_2(mux_tmp_3414, nor_tmp_4, fsm_output(2));
  mux_tmp_3417 <= MUX_s_1_2_2((fsm_output(5)), or_181_cse, fsm_output(2));
  or_tmp_3023 <= (fsm_output(7)) OR mux_tmp_3417;
  mux_3416_nl <= MUX_s_1_2_2((NOT (fsm_output(5))), mux_tmp_3415, fsm_output(7));
  mux_tmp_3418 <= MUX_s_1_2_2(or_tmp_3023, mux_3416_nl, fsm_output(8));
  mux_tmp_3420 <= MUX_s_1_2_2(nor_tmp_4, (fsm_output(5)), fsm_output(7));
  mux_tmp_3421 <= MUX_s_1_2_2((NOT mux_tmp_3420), mux_tmp_14, fsm_output(8));
  mux_tmp_3423 <= MUX_s_1_2_2(and_dcpl_209, (fsm_output(5)), fsm_output(7));
  mux_tmp_3424 <= MUX_s_1_2_2((NOT mux_tmp_14), mux_tmp_3423, fsm_output(8));
  mux_tmp_3425 <= MUX_s_1_2_2(and_dcpl_91, nor_tmp_4, fsm_output(2));
  mux_3426_nl <= MUX_s_1_2_2(mux_tmp_3425, (fsm_output(5)), fsm_output(7));
  mux_3427_nl <= MUX_s_1_2_2((NOT and_350_cse), mux_3426_nl, fsm_output(8));
  not_tmp_663 <= MUX_s_1_2_2(mux_3427_nl, (NOT mux_tmp_3424), fsm_output(6));
  mux_3422_nl <= MUX_s_1_2_2(mux_tmp_3421, mux_tmp_3418, fsm_output(6));
  mux_tmp_3429 <= MUX_s_1_2_2(not_tmp_663, mux_3422_nl, fsm_output(4));
  mux_3430_nl <= MUX_s_1_2_2((NOT (fsm_output(5))), mux_tmp_3425, fsm_output(7));
  mux_3431_nl <= MUX_s_1_2_2(or_3427_cse, mux_3430_nl, fsm_output(8));
  mux_tmp_3432 <= MUX_s_1_2_2(mux_tmp_3421, mux_3431_nl, fsm_output(6));
  mux_3433_nl <= MUX_s_1_2_2((fsm_output(5)), or_181_cse, fsm_output(7));
  mux_tmp_3434 <= MUX_s_1_2_2((NOT mux_3433_nl), and_350_cse, fsm_output(8));
  mux_tmp_3435 <= MUX_s_1_2_2(and_dcpl_91, mux_tmp_3414, fsm_output(2));
  mux_3436_nl <= MUX_s_1_2_2(mux_tmp_3435, (fsm_output(5)), fsm_output(7));
  not_tmp_665 <= MUX_s_1_2_2(and_350_cse, (NOT mux_3436_nl), fsm_output(8));
  mux_3447_nl <= MUX_s_1_2_2(and_dcpl_91, (fsm_output(5)), fsm_output(7));
  mux_3448_nl <= MUX_s_1_2_2(and_350_cse, (NOT mux_3447_nl), fsm_output(8));
  mux_3449_nl <= MUX_s_1_2_2(mux_3448_nl, mux_tmp_3434, fsm_output(6));
  mux_3445_nl <= MUX_s_1_2_2((NOT mux_tmp_3423), mux_tmp_14, fsm_output(8));
  mux_3443_nl <= MUX_s_1_2_2((NOT (fsm_output(5))), mux_tmp_3435, fsm_output(7));
  mux_3444_nl <= MUX_s_1_2_2(or_3427_cse, mux_3443_nl, fsm_output(8));
  mux_3446_nl <= MUX_s_1_2_2(mux_3445_nl, mux_3444_nl, fsm_output(6));
  mux_3450_nl <= MUX_s_1_2_2((NOT mux_3449_nl), mux_3446_nl, fsm_output(4));
  mux_3441_nl <= MUX_s_1_2_2(not_tmp_665, mux_tmp_3424, fsm_output(6));
  mux_3442_nl <= MUX_s_1_2_2((NOT mux_3441_nl), mux_tmp_3432, fsm_output(4));
  mux_3451_nl <= MUX_s_1_2_2(mux_3450_nl, mux_3442_nl, fsm_output(1));
  mux_3438_nl <= MUX_s_1_2_2(not_tmp_665, mux_tmp_3434, fsm_output(6));
  mux_3439_nl <= MUX_s_1_2_2((NOT mux_3438_nl), mux_tmp_3432, fsm_output(4));
  mux_3440_nl <= MUX_s_1_2_2(mux_3439_nl, mux_tmp_3429, fsm_output(1));
  mux_3452_nl <= MUX_s_1_2_2(mux_3451_nl, mux_3440_nl, fsm_output(0));
  or_3090_nl <= CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001")) OR
      mux_tmp_3361;
  mux_3412_nl <= MUX_s_1_2_2(or_3090_nl, mux_tmp_3410, fsm_output(4));
  or_3088_nl <= CONV_SL_1_1(fsm_output(8 DOWNTO 5)/=STD_LOGIC_VECTOR'("0010"));
  mux_3411_nl <= MUX_s_1_2_2(or_3088_nl, mux_tmp_3410, fsm_output(4));
  mux_3413_nl <= MUX_s_1_2_2(mux_3412_nl, mux_3411_nl, fsm_output(1));
  mux_tmp_3453 <= MUX_s_1_2_2(mux_3452_nl, mux_3413_nl, fsm_output(9));
  mux_tmp_3456 <= MUX_s_1_2_2(mux_tmp_3361, mux_tmp_3417, fsm_output(7));
  mux_tmp_3457 <= MUX_s_1_2_2((NOT mux_tmp_3456), or_3427_cse, fsm_output(8));
  mux_3454_nl <= MUX_s_1_2_2((NOT (fsm_output(5))), nor_tmp_4, fsm_output(7));
  mux_3455_nl <= MUX_s_1_2_2(or_tmp_3023, mux_3454_nl, fsm_output(8));
  mux_tmp_3458 <= MUX_s_1_2_2(mux_tmp_3457, mux_3455_nl, fsm_output(6));
  mux_tmp_3459 <= MUX_s_1_2_2(nor_1580_cse, mux_tmp_3420, fsm_output(8));
  mux_3460_nl <= MUX_s_1_2_2(mux_tmp_3415, (fsm_output(5)), fsm_output(7));
  not_tmp_672 <= MUX_s_1_2_2(and_350_cse, (NOT mux_3460_nl), fsm_output(8));
  mux_3462_nl <= MUX_s_1_2_2(not_tmp_672, mux_tmp_3459, fsm_output(6));
  mux_tmp_3463 <= MUX_s_1_2_2((NOT mux_3462_nl), mux_tmp_3458, fsm_output(4));
  mux_tmp_3464 <= MUX_s_1_2_2(nor_tmp_4, mux_tmp_3417, fsm_output(7));
  mux_3469_nl <= MUX_s_1_2_2(not_tmp_672, mux_tmp_3424, fsm_output(6));
  mux_3470_nl <= MUX_s_1_2_2((NOT mux_3469_nl), mux_tmp_3458, fsm_output(4));
  mux_3471_nl <= MUX_s_1_2_2(mux_tmp_3429, mux_3470_nl, fsm_output(1));
  mux_3465_nl <= MUX_s_1_2_2((NOT mux_tmp_3464), or_3427_cse, fsm_output(8));
  mux_3466_nl <= MUX_s_1_2_2(mux_3465_nl, mux_tmp_3418, fsm_output(6));
  mux_3467_nl <= MUX_s_1_2_2(not_tmp_663, mux_3466_nl, fsm_output(4));
  mux_3468_nl <= MUX_s_1_2_2(mux_3467_nl, mux_tmp_3463, fsm_output(1));
  mux_tmp_3472 <= MUX_s_1_2_2(mux_3471_nl, mux_3468_nl, fsm_output(0));
  mux_tmp_3473 <= MUX_s_1_2_2((NOT (fsm_output(5))), mux_tmp_3361, fsm_output(7));
  or_3095_nl <= (fsm_output(7)) OR (fsm_output(5)) OR (fsm_output(3));
  mux_tmp_3474 <= MUX_s_1_2_2(or_3095_nl, mux_tmp_3473, fsm_output(8));
  mux_3475_nl <= MUX_s_1_2_2(mux_tmp_3361, or_181_cse, fsm_output(7));
  mux_3476_nl <= MUX_s_1_2_2((NOT mux_3475_nl), or_3427_cse, fsm_output(8));
  mux_tmp_3477 <= MUX_s_1_2_2(mux_3476_nl, mux_tmp_3474, fsm_output(6));
  mux_3479_nl <= MUX_s_1_2_2(and_350_cse, (NOT mux_tmp_3456), fsm_output(8));
  mux_3478_nl <= MUX_s_1_2_2(nor_1580_cse, mux_tmp_3464, fsm_output(8));
  mux_3480_nl <= MUX_s_1_2_2(mux_3479_nl, mux_3478_nl, fsm_output(6));
  mux_tmp_3481 <= MUX_s_1_2_2((NOT mux_3480_nl), mux_tmp_3477, fsm_output(4));
  mux_3484_nl <= MUX_s_1_2_2(and_350_cse, (NOT mux_tmp_3420), fsm_output(8));
  mux_3485_itm <= MUX_s_1_2_2(mux_3484_nl, mux_tmp_3459, fsm_output(6));
  mux_3488_nl <= MUX_s_1_2_2(and_350_cse, (NOT mux_tmp_3464), fsm_output(8));
  mux_3489_nl <= MUX_s_1_2_2(mux_3488_nl, mux_tmp_3459, fsm_output(6));
  mux_3490_nl <= MUX_s_1_2_2((NOT mux_3489_nl), mux_tmp_3477, fsm_output(4));
  mux_tmp_3491 <= MUX_s_1_2_2(mux_tmp_3463, mux_3490_nl, fsm_output(1));
  mux_3482_nl <= MUX_s_1_2_2(or_tmp_3023, mux_tmp_3473, fsm_output(8));
  mux_3483_nl <= MUX_s_1_2_2(mux_tmp_3457, mux_3482_nl, fsm_output(6));
  mux_3486_nl <= MUX_s_1_2_2((NOT mux_3485_itm), mux_3483_nl, fsm_output(4));
  mux_3487_nl <= MUX_s_1_2_2(mux_3486_nl, mux_tmp_3481, fsm_output(1));
  mux_3492_nl <= MUX_s_1_2_2(mux_tmp_3491, mux_3487_nl, fsm_output(0));
  mux_3493_nl <= MUX_s_1_2_2(mux_3492_nl, mux_tmp_3472, fsm_output(9));
  mux_3494_itm <= MUX_s_1_2_2(mux_3493_nl, mux_tmp_3453, fsm_output(10));
  or_3116_nl <= (fsm_output(1)) OR (fsm_output(6)) OR (NOT (fsm_output(8))) OR (fsm_output(4))
      OR (fsm_output(10));
  or_3115_nl <= (NOT (fsm_output(1))) OR (fsm_output(6)) OR (NOT (fsm_output(8)))
      OR (fsm_output(4)) OR (NOT (fsm_output(10)));
  mux_3504_nl <= MUX_s_1_2_2(or_3116_nl, or_3115_nl, fsm_output(2));
  or_3117_nl <= (fsm_output(9)) OR mux_3504_nl;
  mux_3505_nl <= MUX_s_1_2_2(or_3117_nl, or_70_cse, fsm_output(0));
  nor_603_nl <= NOT((fsm_output(3)) OR mux_3505_nl);
  and_376_nl <= (fsm_output(0)) AND (NOT mux_tmp_2745);
  nor_604_nl <= NOT((fsm_output(2)) OR (fsm_output(1)) OR (fsm_output(6)) OR (fsm_output(8))
      OR not_tmp_39);
  nor_605_nl <= NOT((fsm_output(2)) OR (NOT (fsm_output(1))) OR (NOT (fsm_output(6)))
      OR (NOT (fsm_output(8))) OR (fsm_output(4)) OR (fsm_output(10)));
  mux_3501_nl <= MUX_s_1_2_2(nor_604_nl, nor_605_nl, fsm_output(9));
  nor_606_nl <= NOT((NOT (fsm_output(2))) OR (fsm_output(1)) OR (NOT (fsm_output(6)))
      OR (NOT (fsm_output(8))) OR (fsm_output(4)) OR (NOT (fsm_output(10))));
  nor_607_nl <= NOT((fsm_output(2)) OR (NOT (fsm_output(1))) OR (fsm_output(6)) OR
      (fsm_output(8)) OR not_tmp_39);
  mux_3500_nl <= MUX_s_1_2_2(nor_606_nl, nor_607_nl, fsm_output(9));
  mux_3502_nl <= MUX_s_1_2_2(mux_3501_nl, mux_3500_nl, fsm_output(0));
  mux_3503_nl <= MUX_s_1_2_2(and_376_nl, mux_3502_nl, fsm_output(3));
  mux_3506_nl <= MUX_s_1_2_2(nor_603_nl, mux_3503_nl, fsm_output(5));
  or_3104_nl <= (fsm_output(9)) OR (NOT (fsm_output(2))) OR (fsm_output(1)) OR (NOT((fsm_output(6))
      AND (fsm_output(8)) AND (fsm_output(4)) AND (fsm_output(10))));
  mux_3498_nl <= MUX_s_1_2_2(or_3104_nl, or_56_cse, fsm_output(0));
  or_3098_nl <= (fsm_output(1)) OR (fsm_output(6)) OR (fsm_output(8)) OR (NOT (fsm_output(4)))
      OR (fsm_output(10));
  or_3097_nl <= (NOT (fsm_output(1))) OR (fsm_output(6)) OR (fsm_output(8)) OR not_tmp_39;
  mux_3495_nl <= MUX_s_1_2_2(or_3098_nl, or_3097_nl, fsm_output(2));
  or_3099_nl <= (fsm_output(9)) OR mux_3495_nl;
  mux_3497_nl <= MUX_s_1_2_2(mux_tmp_2745, or_3099_nl, fsm_output(0));
  mux_3499_nl <= MUX_s_1_2_2(mux_3498_nl, mux_3497_nl, fsm_output(3));
  nor_608_nl <= NOT((fsm_output(5)) OR mux_3499_nl);
  not_tmp_688 <= MUX_s_1_2_2(mux_3506_nl, nor_608_nl, fsm_output(7));
  or_tmp_3053 <= (fsm_output(5)) OR (fsm_output(9)) OR (NOT (fsm_output(2))) OR (fsm_output(8))
      OR not_tmp_49;
  or_3154_nl <= (fsm_output(8)) OR nand_183_cse;
  mux_tmp_3529 <= MUX_s_1_2_2(or_3154_nl, or_tmp_2774, fsm_output(3));
  nor_584_nl <= NOT((fsm_output(5)) OR (fsm_output(4)) OR (NOT (fsm_output(7))) OR
      (fsm_output(3)) OR (fsm_output(8)) OR (fsm_output(1)) OR (NOT (fsm_output(6)))
      OR (fsm_output(10)));
  nand_103_nl <= NOT((fsm_output(7)) AND (NOT mux_tmp_3529));
  or_3157_nl <= (NOT (fsm_output(7))) OR (fsm_output(3)) OR (NOT (fsm_output(8)))
      OR (fsm_output(1)) OR (fsm_output(6)) OR (NOT (fsm_output(10)));
  mux_3532_nl <= MUX_s_1_2_2(nand_103_nl, or_3157_nl, fsm_output(4));
  nor_585_nl <= NOT((fsm_output(5)) OR mux_3532_nl);
  mux_3533_nl <= MUX_s_1_2_2(nor_584_nl, nor_585_nl, fsm_output(2));
  nor_586_nl <= NOT((fsm_output(7)) OR mux_tmp_3529);
  nor_587_nl <= NOT((NOT (fsm_output(7))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(8)))
      OR (fsm_output(1)) OR (NOT (fsm_output(6))) OR (fsm_output(10)));
  mux_3530_nl <= MUX_s_1_2_2(nor_586_nl, nor_587_nl, fsm_output(4));
  and_371_nl <= (fsm_output(5)) AND mux_3530_nl;
  nor_588_nl <= NOT((fsm_output(5)) OR (NOT (fsm_output(4))) OR (fsm_output(7)) OR
      (NOT (fsm_output(3))) OR (fsm_output(8)) OR (fsm_output(1)) OR (NOT (fsm_output(6)))
      OR (fsm_output(10)));
  mux_3531_nl <= MUX_s_1_2_2(and_371_nl, nor_588_nl, fsm_output(2));
  mux_3534_nl <= MUX_s_1_2_2(mux_3533_nl, mux_3531_nl, fsm_output(9));
  nor_589_nl <= NOT((fsm_output(3)) OR (fsm_output(8)) OR (NOT (fsm_output(1))) OR
      (fsm_output(6)) OR (fsm_output(10)));
  and_373_nl <= (fsm_output(3)) AND (fsm_output(8)) AND (fsm_output(1)) AND (fsm_output(6))
      AND (fsm_output(10));
  mux_3526_nl <= MUX_s_1_2_2(nor_589_nl, and_373_nl, fsm_output(7));
  and_372_nl <= CONV_SL_1_1(fsm_output(5 DOWNTO 4)=STD_LOGIC_VECTOR'("11")) AND mux_3526_nl;
  nor_590_nl <= NOT((NOT (fsm_output(4))) OR (fsm_output(7)) OR (NOT (fsm_output(3)))
      OR (fsm_output(8)) OR nand_183_cse);
  nor_591_nl <= NOT((fsm_output(7)) OR mux_2998_cse);
  mux_3524_nl <= MUX_s_1_2_2(nor_591_nl, nor_667_cse, fsm_output(4));
  mux_3525_nl <= MUX_s_1_2_2(nor_590_nl, mux_3524_nl, fsm_output(5));
  mux_3527_nl <= MUX_s_1_2_2(and_372_nl, mux_3525_nl, fsm_output(2));
  or_3142_nl <= (NOT (fsm_output(7))) OR (fsm_output(3)) OR (fsm_output(8)) OR (NOT
      (fsm_output(1))) OR (NOT (fsm_output(6))) OR (fsm_output(10));
  or_3141_nl <= (NOT (fsm_output(7))) OR (fsm_output(3)) OR (NOT (fsm_output(8)))
      OR (fsm_output(1)) OR (fsm_output(6)) OR (fsm_output(10));
  mux_3522_nl <= MUX_s_1_2_2(or_3142_nl, or_3141_nl, fsm_output(4));
  nor_593_nl <= NOT((fsm_output(2)) OR (fsm_output(5)) OR mux_3522_nl);
  mux_3528_nl <= MUX_s_1_2_2(mux_3527_nl, nor_593_nl, fsm_output(9));
  not_tmp_701 <= MUX_s_1_2_2(mux_3534_nl, mux_3528_nl, fsm_output(0));
  or_tmp_3095 <= (NOT (fsm_output(4))) OR (fsm_output(9)) OR (fsm_output(6)) OR (fsm_output(8))
      OR (fsm_output(10));
  or_3178_nl <= (fsm_output(2)) OR (fsm_output(4));
  mux_tmp_3547 <= MUX_s_1_2_2(or_2991_cse, mux_tmp_130, or_3178_nl);
  mux_tmp_3551 <= MUX_s_1_2_2(mux_tmp_131, mux_155_cse, fsm_output(2));
  mux_tmp_3574 <= MUX_s_1_2_2(mux_375_cse, mux_340_cse, fsm_output(2));
  mux_460_nl <= MUX_s_1_2_2(mux_tmp_130, or_tmp_94, fsm_output(4));
  mux_tmp_3576 <= MUX_s_1_2_2(or_tmp_96, mux_460_nl, fsm_output(2));
  mux_tmp_3577 <= MUX_s_1_2_2(or_tmp_96, mux_375_cse, fsm_output(2));
  or_3199_nl <= (fsm_output(1)) OR (fsm_output(8)) OR (NOT (fsm_output(6))) OR (fsm_output(10));
  mux_tmp_3618 <= MUX_s_1_2_2(or_3199_nl, or_2835_cse, fsm_output(2));
  or_tmp_3135 <= (NOT (fsm_output(2))) OR (NOT (fsm_output(1))) OR (NOT (fsm_output(8)))
      OR (fsm_output(6)) OR (fsm_output(10));
  or_3222_nl <= (fsm_output(7)) OR (fsm_output(3)) OR (NOT (fsm_output(8))) OR (fsm_output(4))
      OR (fsm_output(10));
  or_3221_nl <= (fsm_output(7)) OR (NOT (fsm_output(3))) OR (fsm_output(8)) OR not_tmp_39;
  mux_tmp_3632 <= MUX_s_1_2_2(or_3222_nl, or_3221_nl, fsm_output(5));
  or_tmp_3176 <= (NOT (fsm_output(4))) OR (fsm_output(8)) OR (NOT (fsm_output(9)))
      OR (fsm_output(6)) OR (fsm_output(10));
  or_tmp_3190 <= (fsm_output(1)) OR (NOT (fsm_output(2))) OR (fsm_output(6)) OR (NOT
      (fsm_output(9)));
  mux_tmp_3673 <= MUX_s_1_2_2(mux_tmp_215, mux_tmp_214, fsm_output(7));
  mux_tmp_3674 <= MUX_s_1_2_2(mux_tmp_215, or_tmp_114, fsm_output(7));
  or_127_nl <= (NOT((fsm_output(5)) OR (NOT (fsm_output(9))))) OR (fsm_output(10));
  mux_tmp_3679 <= MUX_s_1_2_2(or_127_nl, nand_tmp_7, fsm_output(7));
  mux_tmp_3681 <= MUX_s_1_2_2(or_2414_cse, nand_tmp_7, fsm_output(7));
  and_tmp_28 <= (fsm_output(5)) AND or_tmp_104;
  mux_tmp_3691 <= MUX_s_1_2_2(and_tmp_28, or_361_cse, fsm_output(7));
  or_tmp_3224 <= (fsm_output(7)) OR mux_tmp_231;
  or_134_nl <= (fsm_output(5)) OR mux_tmp_227;
  mux_tmp_3698 <= MUX_s_1_2_2(mux_tmp_231, or_134_nl, fsm_output(7));
  mux_262_nl <= MUX_s_1_2_2(and_757_cse, (fsm_output(9)), fsm_output(5));
  mux_tmp_3701 <= MUX_s_1_2_2(mux_262_nl, or_tmp_114, fsm_output(7));
  mux_tmp_3705 <= MUX_s_1_2_2(mux_tmp_236, or_tmp_114, fsm_output(7));
  mux_tmp_3720 <= MUX_s_1_2_2((NOT mux_tmp_214), mux_tmp_228, fsm_output(7));
  mux_tmp_3724 <= MUX_s_1_2_2((NOT and_757_cse), mux_tmp_228, fsm_output(7));
  mux_tmp_3736 <= MUX_s_1_2_2(mux_tmp_227, or_361_cse, fsm_output(5));
  mux_tmp_3737 <= MUX_s_1_2_2(and_tmp_28, mux_tmp_3736, fsm_output(7));
  mux_3738_nl <= MUX_s_1_2_2(or_tmp_104, or_361_cse, fsm_output(5));
  mux_tmp_3739 <= MUX_s_1_2_2(and_tmp_28, mux_3738_nl, fsm_output(7));
  mux_tmp_3753 <= MUX_s_1_2_2(nor_tmp_23, or_tmp_114, fsm_output(7));
  STAGE_LOOP_i_3_0_sva_mx0c1 <= and_dcpl_103 AND and_dcpl_98;
  VEC_LOOP_j_sva_11_0_mx0c1 <= and_dcpl_103 AND and_dcpl_48 AND and_757_cse;
  nor_693_nl <= NOT((fsm_output(2)) OR (fsm_output(1)) OR (fsm_output(7)) OR (fsm_output(9))
      OR (fsm_output(10)));
  mux_2654_nl <= MUX_s_1_2_2(nor_694_cse, nor_693_nl, fsm_output(3));
  and_467_nl <= (fsm_output(0)) AND (fsm_output(1)) AND (fsm_output(7)) AND (fsm_output(9))
      AND (fsm_output(10));
  mux_2653_nl <= MUX_s_1_2_2(and_467_nl, and_756_cse, or_2644_cse);
  mux_2655_nl <= MUX_s_1_2_2(mux_2654_nl, mux_2653_nl, fsm_output(5));
  mux_2656_nl <= MUX_s_1_2_2(mux_2655_nl, and_465_cse, fsm_output(4));
  mux_2657_nl <= MUX_s_1_2_2(mux_2656_nl, and_756_cse, fsm_output(6));
  modExp_result_sva_mx0c0 <= MUX_s_1_2_2(mux_2657_nl, and_757_cse, fsm_output(8));
  STAGE_LOOP_acc_nl <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(STAGE_LOOP_i_3_0_sva_2(3
      DOWNTO 1)) + SIGNED'( "011"), 3));
  STAGE_LOOP_acc_itm_2_1 <= STAGE_LOOP_acc_nl(2);
  and_279_m1c <= and_dcpl_115 AND and_dcpl_44 AND and_dcpl_107;
  and_281_m1c <= and_dcpl_260 AND and_dcpl_88;
  and_284_m1c <= and_dcpl_153 AND and_dcpl_262 AND and_dcpl_144;
  and_286_m1c <= and_dcpl_147 AND and_dcpl_152 AND and_dcpl_235;
  and_288_m1c <= and_dcpl_153 AND and_dcpl_90 AND and_dcpl_162;
  and_291_m1c <= and_dcpl_270 AND and_dcpl_55 AND and_dcpl_33;
  and_292_m1c <= and_dcpl_260 AND and_dcpl_177;
  and_295_m1c <= and_dcpl_6 AND and_dcpl_262 AND and_dcpl_48 AND and_dcpl_33;
  and_297_m1c <= and_dcpl_92 AND and_dcpl_152 AND and_dcpl_162;
  and_299_m1c <= and_dcpl_278 AND and_dcpl_224;
  and_302_m1c <= and_dcpl_270 AND and_dcpl_280 AND and_dcpl_59;
  and_304_m1c <= and_dcpl_118 AND and_dcpl_136 AND and_dcpl_208;
  and_307_m1c <= and_dcpl_209 AND and_dcpl_262 AND and_dcpl_126 AND and_dcpl_59;
  and_309_m1c <= and_dcpl_118 AND and_dcpl_152 AND and_dcpl_224;
  and_311_m1c <= and_dcpl_278 AND and_dcpl_280 AND and_757_cse;
  and_139_nl <= and_dcpl_118 AND and_dcpl_44 AND and_dcpl_88;
  or_522_nl <= (NOT (fsm_output(7))) OR (fsm_output(3)) OR (fsm_output(0)) OR (NOT((fsm_output(1))
      AND (fsm_output(6)) AND (fsm_output(4)) AND (fsm_output(8)) AND (fsm_output(10))));
  or_520_nl <= (fsm_output(7)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(0)))
      OR (NOT (fsm_output(1))) OR (NOT (fsm_output(6))) OR (fsm_output(4)) OR nand_138_cse;
  mux_1091_nl <= MUX_s_1_2_2(or_522_nl, or_520_nl, fsm_output(5));
  or_518_nl <= (fsm_output(3)) OR (fsm_output(0)) OR (fsm_output(1)) OR (fsm_output(6))
      OR (fsm_output(4)) OR nand_138_cse;
  mux_1089_nl <= MUX_s_1_2_2(or_518_nl, mux_tmp_1082, fsm_output(7));
  or_515_nl <= (NOT (fsm_output(1))) OR (fsm_output(6)) OR (NOT (fsm_output(4)))
      OR (fsm_output(8)) OR (NOT (fsm_output(10)));
  mux_1087_nl <= MUX_s_1_2_2(or_515_nl, or_tmp_453, fsm_output(0));
  or_516_nl <= (fsm_output(3)) OR mux_1087_nl;
  or_513_nl <= (NOT (fsm_output(3))) OR (fsm_output(0)) OR (NOT (fsm_output(1)))
      OR (NOT (fsm_output(6))) OR (NOT (fsm_output(4))) OR (fsm_output(8)) OR (fsm_output(10));
  mux_1088_nl <= MUX_s_1_2_2(or_516_nl, or_513_nl, fsm_output(7));
  mux_1090_nl <= MUX_s_1_2_2(mux_1089_nl, mux_1088_nl, fsm_output(5));
  mux_1092_nl <= MUX_s_1_2_2(mux_1091_nl, mux_1090_nl, fsm_output(2));
  or_512_nl <= (fsm_output(3)) OR (NOT (fsm_output(0))) OR (fsm_output(1)) OR (fsm_output(6))
      OR (fsm_output(4)) OR (NOT (fsm_output(8))) OR (fsm_output(10));
  or_511_nl <= (NOT (fsm_output(3))) OR (fsm_output(0)) OR (NOT (fsm_output(1)))
      OR (fsm_output(6)) OR (NOT (fsm_output(4))) OR (fsm_output(8)) OR (fsm_output(10));
  mux_1084_nl <= MUX_s_1_2_2(or_512_nl, or_511_nl, fsm_output(7));
  or_506_nl <= (fsm_output(3)) OR (fsm_output(0)) OR (fsm_output(1)) OR (fsm_output(6))
      OR (fsm_output(4)) OR (fsm_output(8)) OR (NOT (fsm_output(10)));
  mux_1083_nl <= MUX_s_1_2_2(mux_tmp_1082, or_506_nl, fsm_output(7));
  mux_1085_nl <= MUX_s_1_2_2(mux_1084_nl, mux_1083_nl, fsm_output(5));
  or_504_nl <= (fsm_output(5)) OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3)))
      OR (NOT (fsm_output(0))) OR (NOT (fsm_output(1))) OR (NOT (fsm_output(6)))
      OR (fsm_output(4)) OR (NOT (fsm_output(8))) OR (fsm_output(10));
  mux_1086_nl <= MUX_s_1_2_2(mux_1085_nl, or_504_nl, fsm_output(2));
  mux_1093_nl <= MUX_s_1_2_2(mux_1092_nl, mux_1086_nl, fsm_output(9));
  nor_1513_nl <= NOT((fsm_output(1)) OR (NOT (fsm_output(4))) OR (fsm_output(6))
      OR (fsm_output(5)));
  nor_1514_nl <= NOT((NOT (fsm_output(1))) OR (fsm_output(4)) OR (NOT(CONV_SL_1_1(fsm_output(6
      DOWNTO 5)=STD_LOGIC_VECTOR'("11")))));
  mux_1094_nl <= MUX_s_1_2_2(nor_1513_nl, nor_1514_nl, fsm_output(0));
  and_144_nl <= mux_1094_nl AND (fsm_output(3)) AND (NOT (fsm_output(2))) AND (fsm_output(7))
      AND (NOT (fsm_output(8))) AND nor_609_cse;
  nor_1511_nl <= NOT((NOT (fsm_output(8))) OR (fsm_output(7)) OR (fsm_output(2))
      OR (fsm_output(5)) OR (fsm_output(3)));
  nor_1512_nl <= NOT((fsm_output(8)) OR (NOT((fsm_output(7)) AND (fsm_output(2))
      AND (fsm_output(5)) AND (fsm_output(3)))));
  mux_1095_nl <= MUX_s_1_2_2(nor_1511_nl, nor_1512_nl, fsm_output(0));
  and_153_nl <= mux_1095_nl AND (fsm_output(6)) AND (fsm_output(4)) AND (fsm_output(1))
      AND nor_609_cse;
  nor_1509_nl <= NOT((NOT (fsm_output(1))) OR (fsm_output(4)) OR (NOT (fsm_output(6)))
      OR (fsm_output(7)) OR (NOT (fsm_output(2))) OR (fsm_output(3)));
  nor_1510_nl <= NOT((fsm_output(1)) OR (NOT (fsm_output(4))) OR (fsm_output(6))
      OR (NOT (fsm_output(7))) OR (fsm_output(2)) OR (NOT (fsm_output(3))));
  mux_1096_nl <= MUX_s_1_2_2(nor_1509_nl, nor_1510_nl, fsm_output(0));
  and_162_nl <= mux_1096_nl AND and_707_cse AND nor_609_cse;
  and_758_nl <= (fsm_output(0)) AND (fsm_output(6)) AND (fsm_output(8)) AND (fsm_output(7))
      AND (fsm_output(2)) AND (NOT (fsm_output(5))) AND (fsm_output(3));
  nor_1508_nl <= NOT((fsm_output(0)) OR (fsm_output(6)) OR (fsm_output(8)) OR (fsm_output(7))
      OR (fsm_output(2)) OR (NOT (fsm_output(5))) OR (fsm_output(3)));
  mux_1097_nl <= MUX_s_1_2_2(and_758_nl, nor_1508_nl, fsm_output(9));
  and_170_nl <= mux_1097_nl AND and_dcpl_34 AND (NOT (fsm_output(10)));
  nor_1505_nl <= NOT((fsm_output(1)) OR (NOT (fsm_output(4))) OR (fsm_output(7))
      OR (NOT (fsm_output(5))));
  nor_1506_nl <= NOT((NOT (fsm_output(1))) OR (fsm_output(4)) OR (NOT (fsm_output(7)))
      OR (fsm_output(5)));
  mux_1098_nl <= MUX_s_1_2_2(nor_1505_nl, nor_1506_nl, fsm_output(0));
  and_180_nl <= mux_1098_nl AND (NOT (fsm_output(3))) AND (fsm_output(2)) AND (NOT
      (fsm_output(8))) AND (NOT (fsm_output(6))) AND and_dcpl_33;
  nor_1503_nl <= NOT((fsm_output(4)) OR (NOT((fsm_output(6)) AND (fsm_output(2))
      AND (fsm_output(5)))));
  nor_1504_nl <= NOT((NOT (fsm_output(4))) OR (fsm_output(6)) OR (fsm_output(2))
      OR (fsm_output(5)));
  mux_1099_nl <= MUX_s_1_2_2(nor_1503_nl, nor_1504_nl, fsm_output(0));
  and_187_nl <= mux_1099_nl AND (fsm_output(3)) AND and_dcpl_4 AND (fsm_output(1))
      AND and_dcpl_33;
  nor_1501_nl <= NOT((NOT (fsm_output(1))) OR (fsm_output(4)) OR (fsm_output(6))
      OR (fsm_output(2)));
  nor_1502_nl <= NOT((fsm_output(1)) OR (NOT((fsm_output(4)) AND (fsm_output(6))
      AND (fsm_output(2)))));
  mux_1100_nl <= MUX_s_1_2_2(nor_1501_nl, nor_1502_nl, fsm_output(0));
  and_195_nl <= mux_1100_nl AND (NOT (fsm_output(3))) AND nor_1580_cse AND (fsm_output(8))
      AND and_dcpl_33;
  nor_1499_nl <= NOT((NOT (fsm_output(4))) OR (fsm_output(6)) OR (NOT((fsm_output(7))
      AND (fsm_output(2)))));
  nor_1500_nl <= NOT((fsm_output(4)) OR (NOT (fsm_output(6))) OR (fsm_output(7))
      OR (fsm_output(2)));
  mux_1101_nl <= MUX_s_1_2_2(nor_1499_nl, nor_1500_nl, fsm_output(0));
  and_201_nl <= mux_1101_nl AND (fsm_output(3)) AND and_707_cse AND (NOT (fsm_output(1)))
      AND and_dcpl_33;
  or_3445_nl <= (NOT (fsm_output(9))) OR (fsm_output(0)) OR (fsm_output(1)) OR (NOT
      (fsm_output(4))) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(8))) OR (NOT
      (fsm_output(7))) OR (fsm_output(5));
  or_3446_nl <= (fsm_output(9)) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(1)))
      OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(8)) OR (fsm_output(7))
      OR (NOT (fsm_output(5)));
  mux_1102_nl <= MUX_s_1_2_2(or_3445_nl, or_3446_nl, fsm_output(10));
  nor_1625_nl <= NOT(mux_1102_nl OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00")));
  nor_1495_nl <= NOT((fsm_output(4)) OR (NOT (fsm_output(7))) OR (fsm_output(2))
      OR (fsm_output(5)) OR (NOT (fsm_output(3))));
  nor_1496_nl <= NOT((NOT (fsm_output(4))) OR (fsm_output(7)) OR (NOT (fsm_output(2)))
      OR (NOT (fsm_output(5))) OR (fsm_output(3)));
  mux_1103_nl <= MUX_s_1_2_2(nor_1495_nl, nor_1496_nl, fsm_output(0));
  and_213_nl <= mux_1103_nl AND and_dcpl_191 AND (fsm_output(1)) AND and_dcpl_59;
  nor_1493_nl <= NOT((NOT (fsm_output(1))) OR (fsm_output(6)) OR (NOT (fsm_output(2)))
      OR (fsm_output(5)) OR (NOT (fsm_output(3))));
  nor_1494_nl <= NOT((fsm_output(1)) OR (NOT (fsm_output(6))) OR (fsm_output(2))
      OR (NOT (fsm_output(5))) OR (fsm_output(3)));
  mux_1104_nl <= MUX_s_1_2_2(nor_1493_nl, nor_1494_nl, fsm_output(0));
  and_219_nl <= mux_1104_nl AND and_dcpl_4 AND (fsm_output(4)) AND and_dcpl_59;
  and_760_nl <= (fsm_output(4)) AND (fsm_output(6)) AND (NOT (fsm_output(2))) AND
      (fsm_output(3));
  nor_1492_nl <= NOT((fsm_output(4)) OR (fsm_output(6)) OR (NOT (fsm_output(2)))
      OR (fsm_output(3)));
  mux_1105_nl <= MUX_s_1_2_2(and_760_nl, nor_1492_nl, fsm_output(0));
  and_225_nl <= mux_1105_nl AND (NOT (fsm_output(5))) AND and_dcpl_135 AND (NOT (fsm_output(1)))
      AND and_dcpl_59;
  nor_1489_nl <= NOT((fsm_output(1)) OR (fsm_output(4)) OR (NOT (fsm_output(6)))
      OR (fsm_output(7)));
  and_748_nl <= (fsm_output(1)) AND (fsm_output(4)) AND (NOT (fsm_output(6))) AND
      (fsm_output(7));
  mux_1106_nl <= MUX_s_1_2_2(nor_1489_nl, and_748_nl, fsm_output(0));
  and_235_nl <= mux_1106_nl AND (fsm_output(3)) AND and_676_cse AND (fsm_output(8))
      AND and_dcpl_59;
  and_627_nl <= (fsm_output(0)) AND (fsm_output(4)) AND (fsm_output(6)) AND (fsm_output(8))
      AND (fsm_output(7)) AND (NOT (fsm_output(2))) AND (NOT (fsm_output(5)));
  nor_1488_nl <= NOT((fsm_output(0)) OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(8))
      OR (fsm_output(7)) OR (NOT and_676_cse));
  mux_1107_nl <= MUX_s_1_2_2(and_627_nl, nor_1488_nl, fsm_output(9));
  and_241_nl <= mux_1107_nl AND (NOT (fsm_output(3))) AND (fsm_output(1)) AND (fsm_output(10));
  nor_1486_nl <= NOT((NOT (fsm_output(1))) OR (NOT (fsm_output(4))) OR (fsm_output(7))
      OR (fsm_output(2)) OR (NOT (fsm_output(5))));
  nor_1487_nl <= NOT((fsm_output(1)) OR (fsm_output(4)) OR (NOT (fsm_output(7)))
      OR (NOT (fsm_output(2))) OR (fsm_output(5)));
  mux_1108_nl <= MUX_s_1_2_2(nor_1486_nl, nor_1487_nl, fsm_output(0));
  and_249_nl <= mux_1108_nl AND (fsm_output(3)) AND (NOT (fsm_output(8))) AND (NOT
      (fsm_output(6))) AND and_757_cse;
  vec_rsc_0_0_i_adra_d_pff <= MUX1HOT_v_8_19_2(COMP_LOOP_acc_psp_sva_1, (z_out_2_12_1(11
      DOWNTO 4)), COMP_LOOP_acc_psp_sva, (COMP_LOOP_acc_10_cse_12_1_1_sva(11 DOWNTO
      4)), (COMP_LOOP_acc_1_cse_2_sva(11 DOWNTO 4)), (COMP_LOOP_acc_11_psp_sva(10
      DOWNTO 3)), (COMP_LOOP_acc_1_cse_4_sva(11 DOWNTO 4)), (COMP_LOOP_acc_13_psp_sva(9
      DOWNTO 2)), (COMP_LOOP_acc_1_cse_6_sva(11 DOWNTO 4)), (COMP_LOOP_acc_14_psp_sva(10
      DOWNTO 3)), (COMP_LOOP_acc_1_cse_8_sva(11 DOWNTO 4)), (COMP_LOOP_acc_16_psp_sva(8
      DOWNTO 1)), (COMP_LOOP_acc_1_cse_10_sva(11 DOWNTO 4)), (COMP_LOOP_acc_17_psp_sva(10
      DOWNTO 3)), (COMP_LOOP_acc_1_cse_12_sva(11 DOWNTO 4)), (COMP_LOOP_acc_19_psp_sva(9
      DOWNTO 2)), (COMP_LOOP_acc_1_cse_14_sva(11 DOWNTO 4)), (COMP_LOOP_acc_20_psp_sva(10
      DOWNTO 3)), (COMP_LOOP_acc_1_cse_sva(11 DOWNTO 4)), STD_LOGIC_VECTOR'( and_dcpl_109
      & COMP_LOOP_or_32_cse & and_139_nl & (NOT mux_1093_nl) & and_144_nl & and_153_nl
      & and_162_nl & and_170_nl & and_180_nl & and_187_nl & and_195_nl & and_201_nl
      & nor_1625_nl & and_213_nl & and_219_nl & and_225_nl & and_235_nl & and_241_nl
      & and_249_nl));
  vec_rsc_0_0_i_da_d_pff <= COMP_LOOP_10_mul_mut;
  or_618_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR
      (NOT (fsm_output(9))) OR (NOT (fsm_output(5))) OR (fsm_output(10));
  or_617_nl <= (NOT (fsm_output(9))) OR (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")) OR (NOT (fsm_output(10)));
  mux_1134_nl <= MUX_s_1_2_2(or_618_nl, or_617_nl, fsm_output(7));
  or_615_nl <= CONV_SL_1_1(VEC_LOOP_j_sva_11_0(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT (fsm_output(7))) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (fsm_output(9)) OR (fsm_output(5)) OR (fsm_output(10));
  mux_1135_nl <= MUX_s_1_2_2(mux_1134_nl, or_615_nl, fsm_output(2));
  nor_1471_nl <= NOT((fsm_output(6)) OR (fsm_output(4)) OR mux_1135_nl);
  nor_1472_nl <= NOT((fsm_output(6)) OR (fsm_output(4)) OR (NOT (fsm_output(2)))
      OR (fsm_output(7)) OR (fsm_output(9)) OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")) OR (NOT (fsm_output(10))));
  mux_1136_nl <= MUX_s_1_2_2(nor_1471_nl, nor_1472_nl, fsm_output(8));
  nor_1473_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT (fsm_output(6))) OR (NOT (fsm_output(4))) OR (fsm_output(2)) OR (NOT
      (fsm_output(7))) OR (fsm_output(9)) OR not_tmp_248);
  nor_1474_nl <= NOT((fsm_output(4)) OR (fsm_output(2)) OR (fsm_output(7)) OR (NOT
      (fsm_output(9))) OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")) OR (fsm_output(10)));
  nor_1475_nl <= NOT((NOT (fsm_output(2))) OR (fsm_output(7)) OR (fsm_output(9))
      OR (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("0000")) OR (fsm_output(10)));
  nor_1476_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT (fsm_output(2))) OR (fsm_output(7)) OR (NOT (fsm_output(9))) OR (fsm_output(5))
      OR (fsm_output(10)));
  mux_1131_nl <= MUX_s_1_2_2(nor_1475_nl, nor_1476_nl, fsm_output(4));
  mux_1132_nl <= MUX_s_1_2_2(nor_1474_nl, mux_1131_nl, fsm_output(6));
  mux_1133_nl <= MUX_s_1_2_2(nor_1473_nl, mux_1132_nl, fsm_output(8));
  mux_1137_nl <= MUX_s_1_2_2(mux_1136_nl, mux_1133_nl, fsm_output(0));
  or_606_nl <= (COMP_LOOP_acc_16_psp_sva(0)) OR (NOT (fsm_output(4))) OR (NOT (fsm_output(2)))
      OR (VEC_LOOP_j_sva_11_0(2)) OR (NOT (fsm_output(7))) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(5)))
      OR (fsm_output(10));
  or_605_nl <= CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (fsm_output(2)) OR (fsm_output(7)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR (fsm_output(9)) OR (fsm_output(5)) OR
      (NOT (fsm_output(10)));
  mux_1128_nl <= MUX_s_1_2_2(mux_tmp_1116, or_605_nl, fsm_output(4));
  mux_1129_nl <= MUX_s_1_2_2(or_606_nl, mux_1128_nl, fsm_output(6));
  and_626_nl <= (fsm_output(8)) AND (NOT mux_1129_nl);
  or_602_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(7))) OR (NOT (fsm_output(9)))
      OR (fsm_output(5)) OR (NOT (fsm_output(10)));
  or_600_nl <= (fsm_output(7)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(5)))
      OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT (fsm_output(10)));
  mux_1125_nl <= MUX_s_1_2_2(or_600_nl, or_tmp_532, fsm_output(2));
  mux_1126_nl <= MUX_s_1_2_2(or_602_nl, mux_1125_nl, fsm_output(4));
  nor_1477_nl <= NOT((fsm_output(6)) OR mux_1126_nl);
  nor_1478_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(6)) OR (NOT (fsm_output(4))) OR (fsm_output(2)) OR (NOT (fsm_output(7)))
      OR (fsm_output(9)) OR (NOT (fsm_output(5))) OR (fsm_output(10)));
  mux_1127_nl <= MUX_s_1_2_2(nor_1477_nl, nor_1478_nl, fsm_output(8));
  mux_1130_nl <= MUX_s_1_2_2(and_626_nl, mux_1127_nl, fsm_output(0));
  mux_1138_nl <= MUX_s_1_2_2(mux_1137_nl, mux_1130_nl, fsm_output(3));
  or_596_nl <= CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (NOT (fsm_output(2))) OR (fsm_output(7)) OR (VEC_LOOP_j_sva_11_0(0)) OR
      nand_337_cse;
  or_594_nl <= (NOT (fsm_output(2))) OR (fsm_output(7)) OR (fsm_output(9)) OR (NOT
      (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT (fsm_output(10)));
  mux_1121_nl <= MUX_s_1_2_2(or_596_nl, or_594_nl, fsm_output(4));
  nor_1479_nl <= NOT((fsm_output(6)) OR mux_1121_nl);
  or_590_nl <= (fsm_output(9)) OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")) OR (NOT (fsm_output(10)));
  mux_1119_nl <= MUX_s_1_2_2(or_591_cse, or_590_nl, fsm_output(7));
  mux_1120_nl <= MUX_s_1_2_2(mux_1119_nl, or_tmp_532, or_586_cse);
  nor_1480_nl <= NOT((NOT (fsm_output(6))) OR (NOT (fsm_output(4))) OR (fsm_output(2))
      OR mux_1120_nl);
  mux_1122_nl <= MUX_s_1_2_2(nor_1479_nl, nor_1480_nl, fsm_output(8));
  or_583_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(7)) OR (fsm_output(9)) OR not_tmp_248;
  or_581_nl <= (NOT (fsm_output(7))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("0000")) OR (NOT (fsm_output(9))) OR (fsm_output(5))
      OR (fsm_output(10));
  mux_1117_nl <= MUX_s_1_2_2(or_583_nl, or_581_nl, fsm_output(2));
  mux_1118_nl <= MUX_s_1_2_2(mux_1117_nl, mux_tmp_1116, fsm_output(4));
  nor_1481_nl <= NOT((fsm_output(8)) OR (fsm_output(6)) OR mux_1118_nl);
  mux_1123_nl <= MUX_s_1_2_2(mux_1122_nl, nor_1481_nl, fsm_output(0));
  or_576_nl <= CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (fsm_output(2)) OR (NOT (fsm_output(7))) OR (VEC_LOOP_j_sva_11_0(0)) OR
      (fsm_output(9)) OR (fsm_output(5)) OR (NOT (fsm_output(10)));
  or_574_nl <= (fsm_output(2)) OR (NOT (fsm_output(7))) OR (NOT (fsm_output(9)))
      OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("0000")) OR (fsm_output(10));
  mux_1113_nl <= MUX_s_1_2_2(or_576_nl, or_574_nl, fsm_output(4));
  or_573_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(7))) OR (VEC_LOOP_j_sva_11_0(0))
      OR (NOT (fsm_output(9))) OR (NOT (fsm_output(5))) OR (fsm_output(10));
  or_572_nl <= (NOT (fsm_output(2))) OR (NOT (fsm_output(7))) OR (fsm_output(9))
      OR (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("0000")) OR (fsm_output(10));
  mux_1112_nl <= MUX_s_1_2_2(or_573_nl, or_572_nl, fsm_output(4));
  mux_1114_nl <= MUX_s_1_2_2(mux_1113_nl, mux_1112_nl, fsm_output(6));
  nor_1482_nl <= NOT((fsm_output(8)) OR mux_1114_nl);
  nor_1483_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT (fsm_output(6))) OR (fsm_output(4)) OR (fsm_output(2)) OR (NOT (fsm_output(7)))
      OR (fsm_output(9)) OR (NOT (fsm_output(5))) OR (fsm_output(10)));
  nor_1484_nl <= NOT((NOT (fsm_output(4))) OR (NOT (fsm_output(2))) OR (NOT (fsm_output(7)))
      OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(9)) OR not_tmp_248);
  or_567_nl <= (fsm_output(7)) OR (fsm_output(9)) OR (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")) OR (NOT (fsm_output(10)));
  or_565_nl <= (NOT (fsm_output(7))) OR (NOT (fsm_output(9))) OR (fsm_output(5))
      OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(10));
  mux_1109_nl <= MUX_s_1_2_2(or_567_nl, or_565_nl, fsm_output(2));
  nor_1485_nl <= NOT((fsm_output(4)) OR mux_1109_nl);
  mux_1110_nl <= MUX_s_1_2_2(nor_1484_nl, nor_1485_nl, fsm_output(6));
  mux_1111_nl <= MUX_s_1_2_2(nor_1483_nl, mux_1110_nl, fsm_output(8));
  mux_1115_nl <= MUX_s_1_2_2(nor_1482_nl, mux_1111_nl, fsm_output(0));
  mux_1124_nl <= MUX_s_1_2_2(mux_1123_nl, mux_1115_nl, fsm_output(3));
  vec_rsc_0_0_i_wea_d_pff <= MUX_s_1_2_2(mux_1138_nl, mux_1124_nl, fsm_output(1));
  or_674_nl <= (NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(2))) OR (fsm_output(10));
  or_673_nl <= (fsm_output(7)) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(2)) OR (NOT (fsm_output(10)));
  mux_1169_nl <= MUX_s_1_2_2(or_674_nl, or_673_nl, fsm_output(5));
  nor_1440_nl <= NOT((fsm_output(1)) OR mux_1169_nl);
  nor_1441_nl <= NOT((fsm_output(5)) OR (NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")) OR (fsm_output(3)) OR (fsm_output(9))
      OR (fsm_output(2)) OR (fsm_output(10)));
  nor_1442_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT (fsm_output(7))) OR (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_253);
  nor_1443_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(7)) OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (fsm_output(2))
      OR (NOT (fsm_output(10))));
  mux_1167_nl <= MUX_s_1_2_2(nor_1442_nl, nor_1443_nl, fsm_output(5));
  mux_1168_nl <= MUX_s_1_2_2(nor_1441_nl, mux_1167_nl, fsm_output(1));
  mux_1170_nl <= MUX_s_1_2_2(nor_1440_nl, mux_1168_nl, fsm_output(0));
  and_623_nl <= (fsm_output(6)) AND mux_1170_nl;
  nor_1444_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR (fsm_output(2)) OR (fsm_output(10)));
  nor_1446_nl <= NOT((fsm_output(7)) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR not_tmp_253);
  mux_1162_nl <= MUX_s_1_2_2(nor_1445_cse, nor_1446_nl, fsm_output(5));
  nor_1447_nl <= NOT((NOT (fsm_output(5))) OR (fsm_output(7)) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR not_tmp_253);
  or_660_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm);
  mux_1163_nl <= MUX_s_1_2_2(mux_1162_nl, nor_1447_nl, or_660_nl);
  mux_1164_nl <= MUX_s_1_2_2(nor_1444_nl, mux_1163_nl, fsm_output(1));
  nor_1448_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR
      (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_253);
  nor_1449_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (NOT
      (fsm_output(2))) OR (fsm_output(10)));
  nor_1450_nl <= NOT((fsm_output(7)) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9))) OR (fsm_output(2)) OR (fsm_output(10)));
  mux_1160_nl <= MUX_s_1_2_2(nor_1449_nl, nor_1450_nl, fsm_output(5));
  mux_1161_nl <= MUX_s_1_2_2(nor_1448_nl, mux_1160_nl, fsm_output(1));
  mux_1165_nl <= MUX_s_1_2_2(mux_1164_nl, mux_1161_nl, fsm_output(0));
  nor_1451_nl <= NOT((NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (NOT (fsm_output(5)))
      OR (fsm_output(7)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR not_tmp_253);
  nor_1452_nl <= NOT((NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (NOT (fsm_output(5)))
      OR (fsm_output(7)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(3)) OR (fsm_output(9)) OR (NOT (fsm_output(2))) OR (fsm_output(10)));
  mux_1158_nl <= MUX_s_1_2_2(nor_1451_nl, nor_1452_nl, fsm_output(1));
  nor_1453_nl <= NOT((fsm_output(1)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO
      0)/=STD_LOGIC_VECTOR'("00")) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR mux_1157_cse);
  mux_1159_nl <= MUX_s_1_2_2(mux_1158_nl, nor_1453_nl, fsm_output(0));
  mux_1166_nl <= MUX_s_1_2_2(mux_1165_nl, mux_1159_nl, fsm_output(6));
  mux_1171_nl <= MUX_s_1_2_2(and_623_nl, mux_1166_nl, fsm_output(8));
  nor_1454_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (fsm_output(2))
      OR (fsm_output(10)));
  nor_1455_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(7)) OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(2)))
      OR (fsm_output(10)));
  mux_1152_nl <= MUX_s_1_2_2(nor_1454_nl, nor_1455_nl, fsm_output(5));
  and_624_nl <= COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm AND mux_1152_nl;
  nor_1456_nl <= NOT((NOT (fsm_output(7))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR not_tmp_253);
  nor_1457_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(7)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9))) OR (fsm_output(2))
      OR (NOT (fsm_output(10))));
  mux_1151_nl <= MUX_s_1_2_2(nor_1456_nl, nor_1457_nl, fsm_output(5));
  and_625_nl <= COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm AND mux_1151_nl;
  mux_1153_nl <= MUX_s_1_2_2(and_624_nl, and_625_nl, fsm_output(1));
  nor_1458_nl <= NOT((VEC_LOOP_j_sva_11_0(3)) OR (VEC_LOOP_j_sva_11_0(1)) OR (VEC_LOOP_j_sva_11_0(0))
      OR (NOT (fsm_output(5))) OR (VEC_LOOP_j_sva_11_0(2)) OR (fsm_output(7)) OR
      (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(2)) OR (fsm_output(10)));
  nor_1459_nl <= NOT((VEC_LOOP_j_sva_11_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR mux_1149_cse);
  mux_1150_nl <= MUX_s_1_2_2(nor_1458_nl, nor_1459_nl, fsm_output(1));
  mux_1154_nl <= MUX_s_1_2_2(mux_1153_nl, mux_1150_nl, fsm_output(0));
  nor_1460_nl <= NOT((NOT (fsm_output(1))) OR (fsm_output(5)) OR (fsm_output(7))
      OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")) OR (NOT
      (fsm_output(3))) OR (fsm_output(9)) OR (fsm_output(2)) OR (fsm_output(10)));
  nor_1461_nl <= NOT((fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(3)))
      OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")) OR (NOT
      (fsm_output(9))) OR (NOT (fsm_output(2))) OR (fsm_output(10)));
  nor_1462_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (VEC_LOOP_j_sva_11_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR
      (NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3))) OR
      (fsm_output(9)) OR (NOT (fsm_output(2))) OR (fsm_output(10)));
  mux_1147_nl <= MUX_s_1_2_2(nor_1461_nl, nor_1462_nl, fsm_output(1));
  mux_1148_nl <= MUX_s_1_2_2(nor_1460_nl, mux_1147_nl, fsm_output(0));
  mux_1155_nl <= MUX_s_1_2_2(mux_1154_nl, mux_1148_nl, fsm_output(6));
  nor_1463_nl <= NOT((NOT (fsm_output(1))) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(3)) OR (NOT (fsm_output(9)))
      OR (fsm_output(2)) OR (fsm_output(10)));
  nor_1464_nl <= NOT((fsm_output(1)) OR (fsm_output(5)) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")) OR (NOT (fsm_output(7))) OR (fsm_output(3))
      OR (fsm_output(9)) OR not_tmp_253);
  mux_1145_nl <= MUX_s_1_2_2(nor_1463_nl, nor_1464_nl, fsm_output(0));
  nor_1465_nl <= NOT((NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR not_tmp_253);
  nor_1466_nl <= NOT((NOT (fsm_output(7))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")) OR (fsm_output(3)) OR (NOT (fsm_output(9)))
      OR (fsm_output(2)) OR (fsm_output(10)));
  nor_1467_nl <= NOT((NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR not_tmp_253);
  mux_1141_nl <= MUX_s_1_2_2(nor_1466_nl, nor_1467_nl, fsm_output(5));
  mux_1142_nl <= MUX_s_1_2_2(nor_1465_nl, mux_1141_nl, COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm);
  nor_1468_nl <= NOT((NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")) OR (fsm_output(3)) OR (fsm_output(9))
      OR (NOT (fsm_output(2))) OR (fsm_output(10)));
  mux_1143_nl <= MUX_s_1_2_2(mux_1142_nl, nor_1468_nl, fsm_output(1));
  nor_1469_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3)))
      OR (NOT (fsm_output(9))) OR (fsm_output(2)) OR (fsm_output(10)));
  nor_1470_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (VEC_LOOP_j_sva_11_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR
      (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(3)) OR (fsm_output(9))
      OR (fsm_output(2)) OR (NOT (fsm_output(10))));
  mux_1140_nl <= MUX_s_1_2_2(nor_1469_nl, nor_1470_nl, fsm_output(1));
  mux_1144_nl <= MUX_s_1_2_2(mux_1143_nl, mux_1140_nl, fsm_output(0));
  mux_1146_nl <= MUX_s_1_2_2(mux_1145_nl, mux_1144_nl, fsm_output(6));
  mux_1156_nl <= MUX_s_1_2_2(mux_1155_nl, mux_1146_nl, fsm_output(8));
  vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_1171_nl, mux_1156_nl,
      fsm_output(4));
  or_729_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR
      (NOT (fsm_output(9))) OR (NOT (fsm_output(5))) OR (fsm_output(10));
  or_728_nl <= (NOT (fsm_output(9))) OR (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0001")) OR (NOT (fsm_output(10)));
  mux_1198_nl <= MUX_s_1_2_2(or_729_nl, or_728_nl, fsm_output(7));
  or_726_nl <= CONV_SL_1_1(VEC_LOOP_j_sva_11_0(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT (fsm_output(7))) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR (fsm_output(9)) OR (fsm_output(5)) OR (fsm_output(10));
  mux_1199_nl <= MUX_s_1_2_2(mux_1198_nl, or_726_nl, fsm_output(2));
  nor_1425_nl <= NOT((fsm_output(6)) OR (fsm_output(4)) OR mux_1199_nl);
  nor_1426_nl <= NOT((fsm_output(6)) OR (fsm_output(4)) OR (NOT (fsm_output(2)))
      OR (fsm_output(7)) OR (fsm_output(9)) OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0001")) OR (NOT (fsm_output(10))));
  mux_1200_nl <= MUX_s_1_2_2(nor_1425_nl, nor_1426_nl, fsm_output(8));
  nor_1427_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT (fsm_output(6))) OR (NOT (fsm_output(4))) OR (fsm_output(2)) OR (NOT
      (fsm_output(7))) OR (fsm_output(9)) OR not_tmp_248);
  nor_1428_nl <= NOT((fsm_output(4)) OR (fsm_output(2)) OR (fsm_output(7)) OR (NOT
      (fsm_output(9))) OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0001")) OR (fsm_output(10)));
  nor_1429_nl <= NOT((NOT (fsm_output(2))) OR (fsm_output(7)) OR (fsm_output(9))
      OR (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("0001")) OR (fsm_output(10)));
  nor_1430_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT (fsm_output(2))) OR (fsm_output(7)) OR (NOT (fsm_output(9))) OR (fsm_output(5))
      OR (fsm_output(10)));
  mux_1195_nl <= MUX_s_1_2_2(nor_1429_nl, nor_1430_nl, fsm_output(4));
  mux_1196_nl <= MUX_s_1_2_2(nor_1428_nl, mux_1195_nl, fsm_output(6));
  mux_1197_nl <= MUX_s_1_2_2(nor_1427_nl, mux_1196_nl, fsm_output(8));
  mux_1201_nl <= MUX_s_1_2_2(mux_1200_nl, mux_1197_nl, fsm_output(0));
  or_717_nl <= (COMP_LOOP_acc_16_psp_sva(0)) OR (NOT (fsm_output(4))) OR (NOT (fsm_output(2)))
      OR (VEC_LOOP_j_sva_11_0(2)) OR (NOT (fsm_output(7))) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(5)))
      OR (fsm_output(10));
  or_716_nl <= CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (fsm_output(2)) OR (fsm_output(7)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR (fsm_output(9)) OR (fsm_output(5)) OR
      (NOT (fsm_output(10)));
  mux_1192_nl <= MUX_s_1_2_2(mux_tmp_1180, or_716_nl, fsm_output(4));
  mux_1193_nl <= MUX_s_1_2_2(or_717_nl, mux_1192_nl, fsm_output(6));
  and_622_nl <= (fsm_output(8)) AND (NOT mux_1193_nl);
  or_713_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(7))) OR (NOT (fsm_output(9)))
      OR (fsm_output(5)) OR (NOT (fsm_output(10)));
  or_711_nl <= (fsm_output(7)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(5)))
      OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT (fsm_output(10)));
  mux_1189_nl <= MUX_s_1_2_2(or_711_nl, or_tmp_643, fsm_output(2));
  mux_1190_nl <= MUX_s_1_2_2(or_713_nl, mux_1189_nl, fsm_output(4));
  nor_1431_nl <= NOT((fsm_output(6)) OR mux_1190_nl);
  nor_1432_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(6)) OR (NOT (fsm_output(4))) OR (fsm_output(2)) OR (NOT (fsm_output(7)))
      OR (fsm_output(9)) OR (NOT (fsm_output(5))) OR (fsm_output(10)));
  mux_1191_nl <= MUX_s_1_2_2(nor_1431_nl, nor_1432_nl, fsm_output(8));
  mux_1194_nl <= MUX_s_1_2_2(and_622_nl, mux_1191_nl, fsm_output(0));
  mux_1202_nl <= MUX_s_1_2_2(mux_1201_nl, mux_1194_nl, fsm_output(3));
  or_707_nl <= CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (NOT (fsm_output(2))) OR (fsm_output(7)) OR nand_334_cse;
  or_705_nl <= (NOT (fsm_output(2))) OR (fsm_output(7)) OR (fsm_output(9)) OR (NOT
      (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT (fsm_output(10)));
  mux_1185_nl <= MUX_s_1_2_2(or_707_nl, or_705_nl, fsm_output(4));
  nor_1433_nl <= NOT((fsm_output(6)) OR mux_1185_nl);
  or_701_nl <= (fsm_output(9)) OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0001")) OR (NOT (fsm_output(10)));
  mux_1183_nl <= MUX_s_1_2_2(or_702_cse, or_701_nl, fsm_output(7));
  mux_1184_nl <= MUX_s_1_2_2(mux_1183_nl, or_tmp_643, or_586_cse);
  nor_1434_nl <= NOT((NOT (fsm_output(6))) OR (NOT (fsm_output(4))) OR (fsm_output(2))
      OR mux_1184_nl);
  mux_1186_nl <= MUX_s_1_2_2(nor_1433_nl, nor_1434_nl, fsm_output(8));
  or_694_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(7)) OR (fsm_output(9)) OR not_tmp_248;
  or_692_nl <= (NOT (fsm_output(7))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("0001")) OR (NOT (fsm_output(9))) OR (fsm_output(5))
      OR (fsm_output(10));
  mux_1181_nl <= MUX_s_1_2_2(or_694_nl, or_692_nl, fsm_output(2));
  mux_1182_nl <= MUX_s_1_2_2(mux_1181_nl, mux_tmp_1180, fsm_output(4));
  nor_1435_nl <= NOT((fsm_output(8)) OR (fsm_output(6)) OR mux_1182_nl);
  mux_1187_nl <= MUX_s_1_2_2(mux_1186_nl, nor_1435_nl, fsm_output(0));
  or_687_nl <= CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (fsm_output(2)) OR (NOT (fsm_output(7))) OR (NOT (VEC_LOOP_j_sva_11_0(0)))
      OR (fsm_output(9)) OR (fsm_output(5)) OR (NOT (fsm_output(10)));
  or_685_nl <= (fsm_output(2)) OR (NOT (fsm_output(7))) OR (NOT (fsm_output(9)))
      OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("0001")) OR (fsm_output(10));
  mux_1177_nl <= MUX_s_1_2_2(or_687_nl, or_685_nl, fsm_output(4));
  or_684_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(7))) OR (NOT (VEC_LOOP_j_sva_11_0(0)))
      OR (NOT (fsm_output(9))) OR (NOT (fsm_output(5))) OR (fsm_output(10));
  or_683_nl <= (NOT (fsm_output(2))) OR (NOT (fsm_output(7))) OR (fsm_output(9))
      OR (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("0001")) OR (fsm_output(10));
  mux_1176_nl <= MUX_s_1_2_2(or_684_nl, or_683_nl, fsm_output(4));
  mux_1178_nl <= MUX_s_1_2_2(mux_1177_nl, mux_1176_nl, fsm_output(6));
  nor_1436_nl <= NOT((fsm_output(8)) OR mux_1178_nl);
  nor_1437_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT (fsm_output(6))) OR (fsm_output(4)) OR (fsm_output(2)) OR (NOT (fsm_output(7)))
      OR (fsm_output(9)) OR (NOT (fsm_output(5))) OR (fsm_output(10)));
  nor_1438_nl <= NOT((NOT (fsm_output(4))) OR (NOT (fsm_output(2))) OR (NOT (fsm_output(7)))
      OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(9)) OR not_tmp_248);
  or_678_nl <= (fsm_output(7)) OR (fsm_output(9)) OR (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0001")) OR (NOT (fsm_output(10)));
  or_676_nl <= (NOT (fsm_output(7))) OR (NOT (fsm_output(9))) OR (fsm_output(5))
      OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(10));
  mux_1173_nl <= MUX_s_1_2_2(or_678_nl, or_676_nl, fsm_output(2));
  nor_1439_nl <= NOT((fsm_output(4)) OR mux_1173_nl);
  mux_1174_nl <= MUX_s_1_2_2(nor_1438_nl, nor_1439_nl, fsm_output(6));
  mux_1175_nl <= MUX_s_1_2_2(nor_1437_nl, mux_1174_nl, fsm_output(8));
  mux_1179_nl <= MUX_s_1_2_2(nor_1436_nl, mux_1175_nl, fsm_output(0));
  mux_1188_nl <= MUX_s_1_2_2(mux_1187_nl, mux_1179_nl, fsm_output(3));
  vec_rsc_0_1_i_wea_d_pff <= MUX_s_1_2_2(mux_1202_nl, mux_1188_nl, fsm_output(1));
  or_785_nl <= (NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(2))) OR (fsm_output(10));
  or_784_nl <= (fsm_output(7)) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(2)) OR (NOT (fsm_output(10)));
  mux_1233_nl <= MUX_s_1_2_2(or_785_nl, or_784_nl, fsm_output(5));
  nor_1394_nl <= NOT((fsm_output(1)) OR mux_1233_nl);
  nor_1395_nl <= NOT((fsm_output(5)) OR (NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0001")) OR (fsm_output(3)) OR (fsm_output(9))
      OR (fsm_output(2)) OR (fsm_output(10)));
  nor_1396_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT (fsm_output(7))) OR (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_253);
  nor_1397_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(7)) OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (fsm_output(2))
      OR (NOT (fsm_output(10))));
  mux_1231_nl <= MUX_s_1_2_2(nor_1396_nl, nor_1397_nl, fsm_output(5));
  mux_1232_nl <= MUX_s_1_2_2(nor_1395_nl, mux_1231_nl, fsm_output(1));
  mux_1234_nl <= MUX_s_1_2_2(nor_1394_nl, mux_1232_nl, fsm_output(0));
  and_619_nl <= (fsm_output(6)) AND mux_1234_nl;
  nor_1398_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR (fsm_output(2)) OR (fsm_output(10)));
  nor_1400_nl <= NOT((fsm_output(7)) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR not_tmp_253);
  mux_1226_nl <= MUX_s_1_2_2(nor_1445_cse, nor_1400_nl, fsm_output(5));
  nor_1401_nl <= NOT((NOT (fsm_output(5))) OR (fsm_output(7)) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0001")) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR not_tmp_253);
  or_771_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm);
  mux_1227_nl <= MUX_s_1_2_2(mux_1226_nl, nor_1401_nl, or_771_nl);
  mux_1228_nl <= MUX_s_1_2_2(nor_1398_nl, mux_1227_nl, fsm_output(1));
  nor_1402_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR
      (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_253);
  nor_1403_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (NOT
      (fsm_output(2))) OR (fsm_output(10)));
  nor_1404_nl <= NOT((fsm_output(7)) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9))) OR (fsm_output(2)) OR (fsm_output(10)));
  mux_1224_nl <= MUX_s_1_2_2(nor_1403_nl, nor_1404_nl, fsm_output(5));
  mux_1225_nl <= MUX_s_1_2_2(nor_1402_nl, mux_1224_nl, fsm_output(1));
  mux_1229_nl <= MUX_s_1_2_2(mux_1228_nl, mux_1225_nl, fsm_output(0));
  nor_1405_nl <= NOT((NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (NOT (fsm_output(5)))
      OR (fsm_output(7)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR not_tmp_253);
  nor_1406_nl <= NOT((NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (NOT (fsm_output(5)))
      OR (fsm_output(7)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(3)) OR (fsm_output(9)) OR (NOT (fsm_output(2))) OR (fsm_output(10)));
  mux_1222_nl <= MUX_s_1_2_2(nor_1405_nl, nor_1406_nl, fsm_output(1));
  nor_1407_nl <= NOT((fsm_output(1)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO
      0)/=STD_LOGIC_VECTOR'("01")) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR mux_1157_cse);
  mux_1223_nl <= MUX_s_1_2_2(mux_1222_nl, nor_1407_nl, fsm_output(0));
  mux_1230_nl <= MUX_s_1_2_2(mux_1229_nl, mux_1223_nl, fsm_output(6));
  mux_1235_nl <= MUX_s_1_2_2(and_619_nl, mux_1230_nl, fsm_output(8));
  nor_1408_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (fsm_output(2))
      OR (fsm_output(10)));
  nor_1409_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(7)) OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(2)))
      OR (fsm_output(10)));
  mux_1216_nl <= MUX_s_1_2_2(nor_1408_nl, nor_1409_nl, fsm_output(5));
  and_620_nl <= COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm AND mux_1216_nl;
  nor_1410_nl <= NOT((NOT (fsm_output(7))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0001")) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR not_tmp_253);
  nor_1411_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(7)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9))) OR (fsm_output(2))
      OR (NOT (fsm_output(10))));
  mux_1215_nl <= MUX_s_1_2_2(nor_1410_nl, nor_1411_nl, fsm_output(5));
  and_621_nl <= COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm AND mux_1215_nl;
  mux_1217_nl <= MUX_s_1_2_2(and_620_nl, and_621_nl, fsm_output(1));
  nor_1412_nl <= NOT((VEC_LOOP_j_sva_11_0(3)) OR (VEC_LOOP_j_sva_11_0(1)) OR (NOT
      (VEC_LOOP_j_sva_11_0(0))) OR (NOT (fsm_output(5))) OR (VEC_LOOP_j_sva_11_0(2))
      OR (fsm_output(7)) OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(2))
      OR (fsm_output(10)));
  nor_1413_nl <= NOT(nand_332_cse OR mux_1149_cse);
  mux_1214_nl <= MUX_s_1_2_2(nor_1412_nl, nor_1413_nl, fsm_output(1));
  mux_1218_nl <= MUX_s_1_2_2(mux_1217_nl, mux_1214_nl, fsm_output(0));
  nor_1414_nl <= NOT((NOT (fsm_output(1))) OR (fsm_output(5)) OR (fsm_output(7))
      OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001")) OR (NOT
      (fsm_output(3))) OR (fsm_output(9)) OR (fsm_output(2)) OR (fsm_output(10)));
  nor_1415_nl <= NOT((fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(3)))
      OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001")) OR (NOT
      (fsm_output(9))) OR (NOT (fsm_output(2))) OR (fsm_output(10)));
  nor_1416_nl <= NOT((NOT (VEC_LOOP_j_sva_11_0(0))) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (NOT
      (fsm_output(2))) OR (fsm_output(10)));
  mux_1211_nl <= MUX_s_1_2_2(nor_1415_nl, nor_1416_nl, fsm_output(1));
  mux_1212_nl <= MUX_s_1_2_2(nor_1414_nl, mux_1211_nl, fsm_output(0));
  mux_1219_nl <= MUX_s_1_2_2(mux_1218_nl, mux_1212_nl, fsm_output(6));
  nor_1417_nl <= NOT((NOT (fsm_output(1))) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(3)) OR (NOT (fsm_output(9)))
      OR (fsm_output(2)) OR (fsm_output(10)));
  nor_1418_nl <= NOT((fsm_output(1)) OR (fsm_output(5)) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0001")) OR (NOT (fsm_output(7))) OR (fsm_output(3))
      OR (fsm_output(9)) OR not_tmp_253);
  mux_1209_nl <= MUX_s_1_2_2(nor_1417_nl, nor_1418_nl, fsm_output(0));
  nor_1419_nl <= NOT((NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0001")) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR not_tmp_253);
  nor_1420_nl <= NOT((NOT (fsm_output(7))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0001")) OR (fsm_output(3)) OR (NOT (fsm_output(9)))
      OR (fsm_output(2)) OR (fsm_output(10)));
  nor_1421_nl <= NOT((NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR not_tmp_253);
  mux_1205_nl <= MUX_s_1_2_2(nor_1420_nl, nor_1421_nl, fsm_output(5));
  mux_1206_nl <= MUX_s_1_2_2(nor_1419_nl, mux_1205_nl, COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm);
  nor_1422_nl <= NOT((NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0001")) OR (fsm_output(3)) OR (fsm_output(9))
      OR (NOT (fsm_output(2))) OR (fsm_output(10)));
  mux_1207_nl <= MUX_s_1_2_2(mux_1206_nl, nor_1422_nl, fsm_output(1));
  nor_1423_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3)))
      OR (NOT (fsm_output(9))) OR (fsm_output(2)) OR (fsm_output(10)));
  nor_1424_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(3)) OR (fsm_output(9))
      OR (fsm_output(2)) OR (NOT (fsm_output(10))));
  mux_1204_nl <= MUX_s_1_2_2(nor_1423_nl, nor_1424_nl, fsm_output(1));
  mux_1208_nl <= MUX_s_1_2_2(mux_1207_nl, mux_1204_nl, fsm_output(0));
  mux_1210_nl <= MUX_s_1_2_2(mux_1209_nl, mux_1208_nl, fsm_output(6));
  mux_1220_nl <= MUX_s_1_2_2(mux_1219_nl, mux_1210_nl, fsm_output(8));
  vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_1235_nl, mux_1220_nl,
      fsm_output(4));
  or_839_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT (VEC_LOOP_j_sva_11_0(1))) OR (NOT (fsm_output(5))) OR (VEC_LOOP_j_sva_11_0(0))
      OR CONV_SL_1_1(fsm_output(10 DOWNTO 9)/=STD_LOGIC_VECTOR'("01"));
  or_838_nl <= (NOT (fsm_output(5))) OR (NOT (fsm_output(9))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0010")) OR (NOT (fsm_output(10)));
  mux_1262_nl <= MUX_s_1_2_2(or_839_nl, or_838_nl, fsm_output(7));
  or_836_nl <= CONV_SL_1_1(VEC_LOOP_j_sva_11_0(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT (fsm_output(7))) OR (NOT (VEC_LOOP_j_sva_11_0(1))) OR (fsm_output(5))
      OR (VEC_LOOP_j_sva_11_0(0)) OR CONV_SL_1_1(fsm_output(10 DOWNTO 9)/=STD_LOGIC_VECTOR'("00"));
  mux_1263_nl <= MUX_s_1_2_2(mux_1262_nl, or_836_nl, fsm_output(2));
  nor_1379_nl <= NOT((fsm_output(6)) OR (fsm_output(4)) OR mux_1263_nl);
  nor_1380_nl <= NOT((fsm_output(6)) OR (fsm_output(4)) OR (NOT (fsm_output(2)))
      OR (fsm_output(7)) OR (fsm_output(5)) OR (fsm_output(9)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0010")) OR (NOT (fsm_output(10))));
  mux_1264_nl <= MUX_s_1_2_2(nor_1379_nl, nor_1380_nl, fsm_output(8));
  nor_1381_nl <= NOT((NOT (fsm_output(6))) OR (NOT (fsm_output(4))) OR (fsm_output(2))
      OR (NOT (fsm_output(7))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("0010")) OR (NOT (fsm_output(5))) OR (fsm_output(9))
      OR (NOT (fsm_output(10))));
  nor_1382_nl <= NOT((fsm_output(4)) OR (fsm_output(2)) OR (fsm_output(7)) OR (fsm_output(5))
      OR (NOT (fsm_output(9))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("0010")) OR (fsm_output(10)));
  nor_1383_nl <= NOT((NOT (fsm_output(2))) OR (fsm_output(7)) OR (NOT (fsm_output(5)))
      OR (fsm_output(9)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("0010")) OR (fsm_output(10)));
  nor_1384_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT (fsm_output(2))) OR (fsm_output(7)) OR (fsm_output(5)) OR (NOT (fsm_output(9)))
      OR (fsm_output(10)));
  mux_1259_nl <= MUX_s_1_2_2(nor_1383_nl, nor_1384_nl, fsm_output(4));
  mux_1260_nl <= MUX_s_1_2_2(nor_1382_nl, mux_1259_nl, fsm_output(6));
  mux_1261_nl <= MUX_s_1_2_2(nor_1381_nl, mux_1260_nl, fsm_output(8));
  mux_1265_nl <= MUX_s_1_2_2(mux_1264_nl, mux_1261_nl, fsm_output(0));
  or_827_nl <= (COMP_LOOP_acc_16_psp_sva(0)) OR (NOT (fsm_output(4))) OR (NOT (fsm_output(2)))
      OR (VEC_LOOP_j_sva_11_0(2)) OR (NOT (fsm_output(7))) OR (NOT (VEC_LOOP_j_sva_11_0(1)))
      OR (NOT (fsm_output(5))) OR (VEC_LOOP_j_sva_11_0(0)) OR CONV_SL_1_1(fsm_output(10
      DOWNTO 9)/=STD_LOGIC_VECTOR'("01"));
  or_826_nl <= CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (fsm_output(2)) OR (fsm_output(7)) OR (NOT (VEC_LOOP_j_sva_11_0(1))) OR
      (fsm_output(5)) OR (VEC_LOOP_j_sva_11_0(0)) OR CONV_SL_1_1(fsm_output(10 DOWNTO
      9)/=STD_LOGIC_VECTOR'("10"));
  mux_1256_nl <= MUX_s_1_2_2(mux_tmp_1244, or_826_nl, fsm_output(4));
  mux_1257_nl <= MUX_s_1_2_2(or_827_nl, mux_1256_nl, fsm_output(6));
  and_618_nl <= (fsm_output(8)) AND (NOT mux_1257_nl);
  or_823_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(7))) OR (fsm_output(5)) OR nand_358_cse;
  or_821_nl <= (fsm_output(7)) OR (NOT (fsm_output(5))) OR (NOT (fsm_output(9)))
      OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT (fsm_output(10)));
  mux_1253_nl <= MUX_s_1_2_2(or_821_nl, or_tmp_756, fsm_output(2));
  mux_1254_nl <= MUX_s_1_2_2(or_823_nl, mux_1253_nl, fsm_output(4));
  nor_1385_nl <= NOT((fsm_output(6)) OR mux_1254_nl);
  nor_1386_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(6)) OR (NOT (fsm_output(4))) OR (fsm_output(2)) OR (NOT (fsm_output(7)))
      OR (NOT (fsm_output(5))) OR (fsm_output(9)) OR (fsm_output(10)));
  mux_1255_nl <= MUX_s_1_2_2(nor_1385_nl, nor_1386_nl, fsm_output(8));
  mux_1258_nl <= MUX_s_1_2_2(and_618_nl, mux_1255_nl, fsm_output(0));
  mux_1266_nl <= MUX_s_1_2_2(mux_1265_nl, mux_1258_nl, fsm_output(3));
  or_817_nl <= CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (NOT (fsm_output(2))) OR (fsm_output(7)) OR (NOT (fsm_output(5))) OR (VEC_LOOP_j_sva_11_0(0))
      OR nand_358_cse;
  or_815_nl <= (NOT (fsm_output(2))) OR (fsm_output(7)) OR (NOT (fsm_output(5)))
      OR (fsm_output(9)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("0010")) OR (NOT (fsm_output(10)));
  mux_1249_nl <= MUX_s_1_2_2(or_817_nl, or_815_nl, fsm_output(4));
  nor_1387_nl <= NOT((fsm_output(6)) OR mux_1249_nl);
  or_809_nl <= (fsm_output(5)) OR (fsm_output(9)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0010")) OR (NOT (fsm_output(10)));
  mux_1247_nl <= MUX_s_1_2_2(or_591_cse, or_809_nl, fsm_output(7));
  mux_1248_nl <= MUX_s_1_2_2(or_tmp_756, mux_1247_nl, nor_209_cse);
  nor_1388_nl <= NOT((NOT (fsm_output(6))) OR (NOT (fsm_output(4))) OR (fsm_output(2))
      OR mux_1248_nl);
  mux_1250_nl <= MUX_s_1_2_2(nor_1387_nl, nor_1388_nl, fsm_output(8));
  or_805_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(7)) OR (NOT (fsm_output(5))) OR (fsm_output(9)) OR (NOT (fsm_output(10)));
  or_803_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT (fsm_output(7))) OR (fsm_output(5)) OR (NOT (fsm_output(9))) OR (fsm_output(10));
  mux_1245_nl <= MUX_s_1_2_2(or_805_nl, or_803_nl, fsm_output(2));
  mux_1246_nl <= MUX_s_1_2_2(mux_1245_nl, mux_tmp_1244, fsm_output(4));
  nor_1389_nl <= NOT((fsm_output(8)) OR (fsm_output(6)) OR mux_1246_nl);
  mux_1251_nl <= MUX_s_1_2_2(mux_1250_nl, nor_1389_nl, fsm_output(0));
  or_798_nl <= CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (fsm_output(2)) OR (NOT (fsm_output(7))) OR (fsm_output(5)) OR (VEC_LOOP_j_sva_11_0(0))
      OR CONV_SL_1_1(fsm_output(10 DOWNTO 9)/=STD_LOGIC_VECTOR'("10"));
  or_796_nl <= (fsm_output(2)) OR (NOT (fsm_output(7))) OR (fsm_output(5)) OR (NOT
      (fsm_output(9))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(10));
  mux_1241_nl <= MUX_s_1_2_2(or_798_nl, or_796_nl, fsm_output(4));
  or_795_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(7))) OR (NOT (fsm_output(5)))
      OR (VEC_LOOP_j_sva_11_0(0)) OR CONV_SL_1_1(fsm_output(10 DOWNTO 9)/=STD_LOGIC_VECTOR'("01"));
  or_794_nl <= (NOT (fsm_output(2))) OR (NOT (fsm_output(7))) OR (NOT (fsm_output(5)))
      OR (fsm_output(9)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("0010")) OR (fsm_output(10));
  mux_1240_nl <= MUX_s_1_2_2(or_795_nl, or_794_nl, fsm_output(4));
  mux_1242_nl <= MUX_s_1_2_2(mux_1241_nl, mux_1240_nl, fsm_output(6));
  nor_1390_nl <= NOT((fsm_output(8)) OR mux_1242_nl);
  nor_1391_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT (fsm_output(6))) OR (fsm_output(4)) OR (fsm_output(2)) OR (NOT (fsm_output(7)))
      OR (NOT (fsm_output(5))) OR (fsm_output(9)) OR (fsm_output(10)));
  nor_1392_nl <= NOT((NOT (fsm_output(4))) OR (NOT (fsm_output(2))) OR (NOT (fsm_output(7)))
      OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT (fsm_output(5))) OR (fsm_output(9)) OR (NOT (fsm_output(10))));
  or_789_nl <= (fsm_output(7)) OR (NOT (fsm_output(5))) OR (fsm_output(9)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0010")) OR (NOT (fsm_output(10)));
  or_787_nl <= (NOT (fsm_output(7))) OR (fsm_output(5)) OR (NOT (fsm_output(9)))
      OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(10));
  mux_1237_nl <= MUX_s_1_2_2(or_789_nl, or_787_nl, fsm_output(2));
  nor_1393_nl <= NOT((fsm_output(4)) OR mux_1237_nl);
  mux_1238_nl <= MUX_s_1_2_2(nor_1392_nl, nor_1393_nl, fsm_output(6));
  mux_1239_nl <= MUX_s_1_2_2(nor_1391_nl, mux_1238_nl, fsm_output(8));
  mux_1243_nl <= MUX_s_1_2_2(nor_1390_nl, mux_1239_nl, fsm_output(0));
  mux_1252_nl <= MUX_s_1_2_2(mux_1251_nl, mux_1243_nl, fsm_output(3));
  vec_rsc_0_2_i_wea_d_pff <= MUX_s_1_2_2(mux_1266_nl, mux_1252_nl, fsm_output(1));
  or_895_nl <= (NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(2))) OR (fsm_output(10));
  or_894_nl <= (fsm_output(7)) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(2)) OR (NOT (fsm_output(10)));
  mux_1297_nl <= MUX_s_1_2_2(or_895_nl, or_894_nl, fsm_output(5));
  nor_1348_nl <= NOT((fsm_output(1)) OR mux_1297_nl);
  nor_1349_nl <= NOT((fsm_output(5)) OR (NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0010")) OR (fsm_output(3)) OR (fsm_output(9))
      OR (fsm_output(2)) OR (fsm_output(10)));
  nor_1350_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT (fsm_output(7))) OR (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_253);
  nor_1351_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(7)) OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (fsm_output(2))
      OR (NOT (fsm_output(10))));
  mux_1295_nl <= MUX_s_1_2_2(nor_1350_nl, nor_1351_nl, fsm_output(5));
  mux_1296_nl <= MUX_s_1_2_2(nor_1349_nl, mux_1295_nl, fsm_output(1));
  mux_1298_nl <= MUX_s_1_2_2(nor_1348_nl, mux_1296_nl, fsm_output(0));
  and_615_nl <= (fsm_output(6)) AND mux_1298_nl;
  nor_1352_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR (fsm_output(2)) OR (fsm_output(10)));
  nor_1354_nl <= NOT((fsm_output(7)) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR not_tmp_253);
  mux_1290_nl <= MUX_s_1_2_2(nor_1445_cse, nor_1354_nl, fsm_output(5));
  nor_1355_nl <= NOT((NOT (fsm_output(5))) OR (fsm_output(7)) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0010")) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR not_tmp_253);
  or_881_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm);
  mux_1291_nl <= MUX_s_1_2_2(mux_1290_nl, nor_1355_nl, or_881_nl);
  mux_1292_nl <= MUX_s_1_2_2(nor_1352_nl, mux_1291_nl, fsm_output(1));
  nor_1356_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR
      (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_253);
  nor_1357_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (NOT
      (fsm_output(2))) OR (fsm_output(10)));
  nor_1358_nl <= NOT((fsm_output(7)) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9))) OR (fsm_output(2)) OR (fsm_output(10)));
  mux_1288_nl <= MUX_s_1_2_2(nor_1357_nl, nor_1358_nl, fsm_output(5));
  mux_1289_nl <= MUX_s_1_2_2(nor_1356_nl, mux_1288_nl, fsm_output(1));
  mux_1293_nl <= MUX_s_1_2_2(mux_1292_nl, mux_1289_nl, fsm_output(0));
  nor_1359_nl <= NOT((NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (NOT (fsm_output(5)))
      OR (fsm_output(7)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR not_tmp_253);
  nor_1360_nl <= NOT((NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (NOT (fsm_output(5)))
      OR (fsm_output(7)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(3)) OR (fsm_output(9)) OR (NOT (fsm_output(2))) OR (fsm_output(10)));
  mux_1286_nl <= MUX_s_1_2_2(nor_1359_nl, nor_1360_nl, fsm_output(1));
  nor_1361_nl <= NOT((fsm_output(1)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO
      0)/=STD_LOGIC_VECTOR'("10")) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR mux_1157_cse);
  mux_1287_nl <= MUX_s_1_2_2(mux_1286_nl, nor_1361_nl, fsm_output(0));
  mux_1294_nl <= MUX_s_1_2_2(mux_1293_nl, mux_1287_nl, fsm_output(6));
  mux_1299_nl <= MUX_s_1_2_2(and_615_nl, mux_1294_nl, fsm_output(8));
  nor_1362_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (fsm_output(2))
      OR (fsm_output(10)));
  nor_1363_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(7)) OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(2)))
      OR (fsm_output(10)));
  mux_1280_nl <= MUX_s_1_2_2(nor_1362_nl, nor_1363_nl, fsm_output(5));
  and_616_nl <= COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm AND mux_1280_nl;
  nor_1364_nl <= NOT((NOT (fsm_output(7))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0010")) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR not_tmp_253);
  nor_1365_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(7)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9))) OR (fsm_output(2))
      OR (NOT (fsm_output(10))));
  mux_1279_nl <= MUX_s_1_2_2(nor_1364_nl, nor_1365_nl, fsm_output(5));
  and_617_nl <= COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm AND mux_1279_nl;
  mux_1281_nl <= MUX_s_1_2_2(and_616_nl, and_617_nl, fsm_output(1));
  nor_1366_nl <= NOT((VEC_LOOP_j_sva_11_0(3)) OR (NOT (VEC_LOOP_j_sva_11_0(1))) OR
      (VEC_LOOP_j_sva_11_0(0)) OR (NOT (fsm_output(5))) OR (VEC_LOOP_j_sva_11_0(2))
      OR (fsm_output(7)) OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(2))
      OR (fsm_output(10)));
  nor_1367_nl <= NOT((VEC_LOOP_j_sva_11_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR mux_1277_cse);
  mux_1278_nl <= MUX_s_1_2_2(nor_1366_nl, nor_1367_nl, fsm_output(1));
  mux_1282_nl <= MUX_s_1_2_2(mux_1281_nl, mux_1278_nl, fsm_output(0));
  nor_1368_nl <= NOT((NOT (fsm_output(1))) OR (fsm_output(5)) OR (fsm_output(7))
      OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010")) OR (NOT
      (fsm_output(3))) OR (fsm_output(9)) OR (fsm_output(2)) OR (fsm_output(10)));
  nor_1369_nl <= NOT((fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(3)))
      OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010")) OR (NOT
      (fsm_output(9))) OR (NOT (fsm_output(2))) OR (fsm_output(10)));
  nor_1370_nl <= NOT((VEC_LOOP_j_sva_11_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (NOT
      (fsm_output(2))) OR (fsm_output(10)));
  mux_1275_nl <= MUX_s_1_2_2(nor_1369_nl, nor_1370_nl, fsm_output(1));
  mux_1276_nl <= MUX_s_1_2_2(nor_1368_nl, mux_1275_nl, fsm_output(0));
  mux_1283_nl <= MUX_s_1_2_2(mux_1282_nl, mux_1276_nl, fsm_output(6));
  nor_1371_nl <= NOT((NOT (fsm_output(1))) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(3)) OR (NOT (fsm_output(9)))
      OR (fsm_output(2)) OR (fsm_output(10)));
  nor_1372_nl <= NOT((fsm_output(1)) OR (fsm_output(5)) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0010")) OR (NOT (fsm_output(7))) OR (fsm_output(3))
      OR (fsm_output(9)) OR not_tmp_253);
  mux_1273_nl <= MUX_s_1_2_2(nor_1371_nl, nor_1372_nl, fsm_output(0));
  nor_1373_nl <= NOT((NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0010")) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR not_tmp_253);
  nor_1374_nl <= NOT((NOT (fsm_output(7))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0010")) OR (fsm_output(3)) OR (NOT (fsm_output(9)))
      OR (fsm_output(2)) OR (fsm_output(10)));
  nor_1375_nl <= NOT((NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR not_tmp_253);
  mux_1269_nl <= MUX_s_1_2_2(nor_1374_nl, nor_1375_nl, fsm_output(5));
  mux_1270_nl <= MUX_s_1_2_2(nor_1373_nl, mux_1269_nl, COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm);
  nor_1376_nl <= NOT((NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0010")) OR (fsm_output(3)) OR (fsm_output(9))
      OR (NOT (fsm_output(2))) OR (fsm_output(10)));
  mux_1271_nl <= MUX_s_1_2_2(mux_1270_nl, nor_1376_nl, fsm_output(1));
  nor_1377_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3)))
      OR (NOT (fsm_output(9))) OR (fsm_output(2)) OR (fsm_output(10)));
  nor_1378_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (VEC_LOOP_j_sva_11_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR
      (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(3)) OR (fsm_output(9))
      OR (fsm_output(2)) OR (NOT (fsm_output(10))));
  mux_1268_nl <= MUX_s_1_2_2(nor_1377_nl, nor_1378_nl, fsm_output(1));
  mux_1272_nl <= MUX_s_1_2_2(mux_1271_nl, mux_1268_nl, fsm_output(0));
  mux_1274_nl <= MUX_s_1_2_2(mux_1273_nl, mux_1272_nl, fsm_output(6));
  mux_1284_nl <= MUX_s_1_2_2(mux_1283_nl, mux_1274_nl, fsm_output(8));
  vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_1299_nl, mux_1284_nl,
      fsm_output(4));
  or_949_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11")) OR
      (NOT (fsm_output(9))) OR (NOT (fsm_output(5))) OR (fsm_output(10));
  nand_404_nl <= NOT((fsm_output(9)) AND (fsm_output(5)) AND CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)=STD_LOGIC_VECTOR'("0011")) AND (fsm_output(10)));
  mux_1326_nl <= MUX_s_1_2_2(or_949_nl, nand_404_nl, fsm_output(7));
  or_946_nl <= CONV_SL_1_1(VEC_LOOP_j_sva_11_0(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT (fsm_output(7))) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR (fsm_output(9)) OR (fsm_output(5)) OR (fsm_output(10));
  mux_1327_nl <= MUX_s_1_2_2(mux_1326_nl, or_946_nl, fsm_output(2));
  nor_1333_nl <= NOT((fsm_output(6)) OR (fsm_output(4)) OR mux_1327_nl);
  nor_1334_nl <= NOT((fsm_output(6)) OR (fsm_output(4)) OR (NOT (fsm_output(2)))
      OR (fsm_output(7)) OR (fsm_output(9)) OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0011")) OR (NOT (fsm_output(10))));
  mux_1328_nl <= MUX_s_1_2_2(nor_1333_nl, nor_1334_nl, fsm_output(8));
  nor_1335_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT (fsm_output(6))) OR (NOT (fsm_output(4))) OR (fsm_output(2)) OR (NOT
      (fsm_output(7))) OR (fsm_output(9)) OR not_tmp_248);
  nor_1336_nl <= NOT((fsm_output(4)) OR (fsm_output(2)) OR (fsm_output(7)) OR (NOT
      (fsm_output(9))) OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0011")) OR (fsm_output(10)));
  nor_1337_nl <= NOT((NOT (fsm_output(2))) OR (fsm_output(7)) OR (fsm_output(9))
      OR (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("0011")) OR (fsm_output(10)));
  nor_1338_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT (fsm_output(2))) OR (fsm_output(7)) OR (NOT (fsm_output(9))) OR (fsm_output(5))
      OR (fsm_output(10)));
  mux_1323_nl <= MUX_s_1_2_2(nor_1337_nl, nor_1338_nl, fsm_output(4));
  mux_1324_nl <= MUX_s_1_2_2(nor_1336_nl, mux_1323_nl, fsm_output(6));
  mux_1325_nl <= MUX_s_1_2_2(nor_1335_nl, mux_1324_nl, fsm_output(8));
  mux_1329_nl <= MUX_s_1_2_2(mux_1328_nl, mux_1325_nl, fsm_output(0));
  nand_327_nl <= NOT((NOT (COMP_LOOP_acc_16_psp_sva(0))) AND (fsm_output(4)) AND
      (fsm_output(2)) AND (NOT (VEC_LOOP_j_sva_11_0(2))) AND (fsm_output(7)) AND
      CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND (fsm_output(9))
      AND (fsm_output(5)) AND (NOT (fsm_output(10))));
  or_936_nl <= CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (fsm_output(2)) OR (fsm_output(7)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("11")) OR (fsm_output(9)) OR (fsm_output(5)) OR
      (NOT (fsm_output(10)));
  mux_1320_nl <= MUX_s_1_2_2(mux_tmp_1308, or_936_nl, fsm_output(4));
  mux_1321_nl <= MUX_s_1_2_2(nand_327_nl, mux_1320_nl, fsm_output(6));
  and_614_nl <= (fsm_output(8)) AND (NOT mux_1321_nl);
  or_933_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(7))) OR (NOT (fsm_output(9)))
      OR (fsm_output(5)) OR (NOT (fsm_output(10)));
  or_931_nl <= (fsm_output(7)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(5)))
      OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT (fsm_output(10)));
  mux_1317_nl <= MUX_s_1_2_2(or_931_nl, or_tmp_866, fsm_output(2));
  mux_1318_nl <= MUX_s_1_2_2(or_933_nl, mux_1317_nl, fsm_output(4));
  nor_1339_nl <= NOT((fsm_output(6)) OR mux_1318_nl);
  nor_1340_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(6)) OR (NOT (fsm_output(4))) OR (fsm_output(2)) OR (NOT (fsm_output(7)))
      OR (fsm_output(9)) OR (NOT (fsm_output(5))) OR (fsm_output(10)));
  mux_1319_nl <= MUX_s_1_2_2(nor_1339_nl, nor_1340_nl, fsm_output(8));
  mux_1322_nl <= MUX_s_1_2_2(and_614_nl, mux_1319_nl, fsm_output(0));
  mux_1330_nl <= MUX_s_1_2_2(mux_1329_nl, mux_1322_nl, fsm_output(3));
  or_927_nl <= CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (NOT (fsm_output(2))) OR (fsm_output(7)) OR nand_334_cse;
  or_925_nl <= (NOT (fsm_output(2))) OR (fsm_output(7)) OR (fsm_output(9)) OR (NOT
      (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT (fsm_output(10)));
  mux_1313_nl <= MUX_s_1_2_2(or_927_nl, or_925_nl, fsm_output(4));
  nor_1341_nl <= NOT((fsm_output(6)) OR mux_1313_nl);
  or_919_nl <= (fsm_output(9)) OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0011")) OR (NOT (fsm_output(10)));
  mux_1311_nl <= MUX_s_1_2_2(or_702_cse, or_919_nl, fsm_output(7));
  mux_1312_nl <= MUX_s_1_2_2(or_tmp_866, mux_1311_nl, nor_209_cse);
  nor_1342_nl <= NOT((NOT (fsm_output(6))) OR (NOT (fsm_output(4))) OR (fsm_output(2))
      OR mux_1312_nl);
  mux_1314_nl <= MUX_s_1_2_2(nor_1341_nl, nor_1342_nl, fsm_output(8));
  or_915_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(7)) OR (fsm_output(9)) OR not_tmp_248;
  or_913_nl <= (NOT (fsm_output(7))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("0011")) OR (NOT (fsm_output(9))) OR (fsm_output(5))
      OR (fsm_output(10));
  mux_1309_nl <= MUX_s_1_2_2(or_915_nl, or_913_nl, fsm_output(2));
  mux_1310_nl <= MUX_s_1_2_2(mux_1309_nl, mux_tmp_1308, fsm_output(4));
  nor_1343_nl <= NOT((fsm_output(8)) OR (fsm_output(6)) OR mux_1310_nl);
  mux_1315_nl <= MUX_s_1_2_2(mux_1314_nl, nor_1343_nl, fsm_output(0));
  or_908_nl <= CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (fsm_output(2)) OR (NOT (fsm_output(7))) OR (NOT (VEC_LOOP_j_sva_11_0(0)))
      OR (fsm_output(9)) OR (fsm_output(5)) OR (NOT (fsm_output(10)));
  or_906_nl <= (fsm_output(2)) OR (NOT (fsm_output(7))) OR (NOT (fsm_output(9)))
      OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("0011")) OR (fsm_output(10));
  mux_1305_nl <= MUX_s_1_2_2(or_908_nl, or_906_nl, fsm_output(4));
  or_905_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(7))) OR (NOT (VEC_LOOP_j_sva_11_0(0)))
      OR (NOT (fsm_output(9))) OR (NOT (fsm_output(5))) OR (fsm_output(10));
  or_904_nl <= (NOT (fsm_output(2))) OR (NOT (fsm_output(7))) OR (fsm_output(9))
      OR (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("0011")) OR (fsm_output(10));
  mux_1304_nl <= MUX_s_1_2_2(or_905_nl, or_904_nl, fsm_output(4));
  mux_1306_nl <= MUX_s_1_2_2(mux_1305_nl, mux_1304_nl, fsm_output(6));
  nor_1344_nl <= NOT((fsm_output(8)) OR mux_1306_nl);
  nor_1345_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT (fsm_output(6))) OR (fsm_output(4)) OR (fsm_output(2)) OR (NOT (fsm_output(7)))
      OR (fsm_output(9)) OR (NOT (fsm_output(5))) OR (fsm_output(10)));
  nor_1346_nl <= NOT((NOT (fsm_output(4))) OR (NOT (fsm_output(2))) OR (NOT (fsm_output(7)))
      OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(9)) OR not_tmp_248);
  or_899_nl <= (fsm_output(7)) OR (fsm_output(9)) OR (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0011")) OR (NOT (fsm_output(10)));
  or_897_nl <= (NOT (fsm_output(7))) OR (NOT (fsm_output(9))) OR (fsm_output(5))
      OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(10));
  mux_1301_nl <= MUX_s_1_2_2(or_899_nl, or_897_nl, fsm_output(2));
  nor_1347_nl <= NOT((fsm_output(4)) OR mux_1301_nl);
  mux_1302_nl <= MUX_s_1_2_2(nor_1346_nl, nor_1347_nl, fsm_output(6));
  mux_1303_nl <= MUX_s_1_2_2(nor_1345_nl, mux_1302_nl, fsm_output(8));
  mux_1307_nl <= MUX_s_1_2_2(nor_1344_nl, mux_1303_nl, fsm_output(0));
  mux_1316_nl <= MUX_s_1_2_2(mux_1315_nl, mux_1307_nl, fsm_output(3));
  vec_rsc_0_3_i_wea_d_pff <= MUX_s_1_2_2(mux_1330_nl, mux_1316_nl, fsm_output(1));
  or_1005_nl <= (NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(2))) OR (fsm_output(10));
  or_1004_nl <= (fsm_output(7)) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(2)) OR (NOT (fsm_output(10)));
  mux_1361_nl <= MUX_s_1_2_2(or_1005_nl, or_1004_nl, fsm_output(5));
  nor_1302_nl <= NOT((fsm_output(1)) OR mux_1361_nl);
  nor_1303_nl <= NOT((fsm_output(5)) OR (NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0011")) OR (fsm_output(3)) OR (fsm_output(9))
      OR (fsm_output(2)) OR (fsm_output(10)));
  nor_1304_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT (fsm_output(7))) OR (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_253);
  nor_1305_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(7)) OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (fsm_output(2))
      OR (NOT (fsm_output(10))));
  mux_1359_nl <= MUX_s_1_2_2(nor_1304_nl, nor_1305_nl, fsm_output(5));
  mux_1360_nl <= MUX_s_1_2_2(nor_1303_nl, mux_1359_nl, fsm_output(1));
  mux_1362_nl <= MUX_s_1_2_2(nor_1302_nl, mux_1360_nl, fsm_output(0));
  and_611_nl <= (fsm_output(6)) AND mux_1362_nl;
  nor_1306_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR (fsm_output(2)) OR (fsm_output(10)));
  nor_1308_nl <= NOT((fsm_output(7)) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR not_tmp_253);
  mux_1354_nl <= MUX_s_1_2_2(nor_1445_cse, nor_1308_nl, fsm_output(5));
  nor_1309_nl <= NOT((NOT (fsm_output(5))) OR (fsm_output(7)) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0011")) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR not_tmp_253);
  or_991_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm);
  mux_1355_nl <= MUX_s_1_2_2(mux_1354_nl, nor_1309_nl, or_991_nl);
  mux_1356_nl <= MUX_s_1_2_2(nor_1306_nl, mux_1355_nl, fsm_output(1));
  nor_1310_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11")) OR
      (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_253);
  nor_1311_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (NOT
      (fsm_output(2))) OR (fsm_output(10)));
  nor_1312_nl <= NOT((fsm_output(7)) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9))) OR (fsm_output(2)) OR (fsm_output(10)));
  mux_1352_nl <= MUX_s_1_2_2(nor_1311_nl, nor_1312_nl, fsm_output(5));
  mux_1353_nl <= MUX_s_1_2_2(nor_1310_nl, mux_1352_nl, fsm_output(1));
  mux_1357_nl <= MUX_s_1_2_2(mux_1356_nl, mux_1353_nl, fsm_output(0));
  nor_1313_nl <= NOT((NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (NOT (fsm_output(5)))
      OR (fsm_output(7)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR not_tmp_253);
  nor_1314_nl <= NOT((NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (NOT (fsm_output(5)))
      OR (fsm_output(7)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(3)) OR (fsm_output(9)) OR (NOT (fsm_output(2))) OR (fsm_output(10)));
  mux_1350_nl <= MUX_s_1_2_2(nor_1313_nl, nor_1314_nl, fsm_output(1));
  nor_1315_nl <= NOT(nand_324_cse OR mux_1157_cse);
  mux_1351_nl <= MUX_s_1_2_2(mux_1350_nl, nor_1315_nl, fsm_output(0));
  mux_1358_nl <= MUX_s_1_2_2(mux_1357_nl, mux_1351_nl, fsm_output(6));
  mux_1363_nl <= MUX_s_1_2_2(and_611_nl, mux_1358_nl, fsm_output(8));
  nor_1316_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (fsm_output(2))
      OR (fsm_output(10)));
  nor_1317_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(7)) OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(2)))
      OR (fsm_output(10)));
  mux_1344_nl <= MUX_s_1_2_2(nor_1316_nl, nor_1317_nl, fsm_output(5));
  and_612_nl <= COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm AND mux_1344_nl;
  nor_1318_nl <= NOT((NOT (fsm_output(7))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0011")) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR not_tmp_253);
  nor_1319_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(7)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9))) OR (fsm_output(2))
      OR (NOT (fsm_output(10))));
  mux_1343_nl <= MUX_s_1_2_2(nor_1318_nl, nor_1319_nl, fsm_output(5));
  and_613_nl <= COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm AND mux_1343_nl;
  mux_1345_nl <= MUX_s_1_2_2(and_612_nl, and_613_nl, fsm_output(1));
  nor_1320_nl <= NOT((VEC_LOOP_j_sva_11_0(3)) OR (NOT (VEC_LOOP_j_sva_11_0(1))) OR
      (NOT (VEC_LOOP_j_sva_11_0(0))) OR (NOT (fsm_output(5))) OR (VEC_LOOP_j_sva_11_0(2))
      OR (fsm_output(7)) OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(2))
      OR (fsm_output(10)));
  nor_1321_nl <= NOT(nand_332_cse OR mux_1277_cse);
  mux_1342_nl <= MUX_s_1_2_2(nor_1320_nl, nor_1321_nl, fsm_output(1));
  mux_1346_nl <= MUX_s_1_2_2(mux_1345_nl, mux_1342_nl, fsm_output(0));
  nor_1322_nl <= NOT((NOT (fsm_output(1))) OR (fsm_output(5)) OR (fsm_output(7))
      OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011")) OR (NOT
      (fsm_output(3))) OR (fsm_output(9)) OR (fsm_output(2)) OR (fsm_output(10)));
  nor_1323_nl <= NOT((fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(3)))
      OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011")) OR (NOT
      (fsm_output(9))) OR (NOT (fsm_output(2))) OR (fsm_output(10)));
  nor_1324_nl <= NOT((NOT (VEC_LOOP_j_sva_11_0(0))) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (NOT
      (fsm_output(2))) OR (fsm_output(10)));
  mux_1339_nl <= MUX_s_1_2_2(nor_1323_nl, nor_1324_nl, fsm_output(1));
  mux_1340_nl <= MUX_s_1_2_2(nor_1322_nl, mux_1339_nl, fsm_output(0));
  mux_1347_nl <= MUX_s_1_2_2(mux_1346_nl, mux_1340_nl, fsm_output(6));
  nor_1325_nl <= NOT((NOT (fsm_output(1))) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(3)) OR (NOT (fsm_output(9)))
      OR (fsm_output(2)) OR (fsm_output(10)));
  nor_1326_nl <= NOT((fsm_output(1)) OR (fsm_output(5)) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0011")) OR (NOT (fsm_output(7))) OR (fsm_output(3))
      OR (fsm_output(9)) OR not_tmp_253);
  mux_1337_nl <= MUX_s_1_2_2(nor_1325_nl, nor_1326_nl, fsm_output(0));
  nor_1327_nl <= NOT((NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0011")) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR not_tmp_253);
  nor_1328_nl <= NOT((NOT (fsm_output(7))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0011")) OR (fsm_output(3)) OR (NOT (fsm_output(9)))
      OR (fsm_output(2)) OR (fsm_output(10)));
  nor_1329_nl <= NOT((NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR not_tmp_253);
  mux_1333_nl <= MUX_s_1_2_2(nor_1328_nl, nor_1329_nl, fsm_output(5));
  mux_1334_nl <= MUX_s_1_2_2(nor_1327_nl, mux_1333_nl, COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm);
  nor_1330_nl <= NOT((NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0011")) OR (fsm_output(3)) OR (fsm_output(9))
      OR (NOT (fsm_output(2))) OR (fsm_output(10)));
  mux_1335_nl <= MUX_s_1_2_2(mux_1334_nl, nor_1330_nl, fsm_output(1));
  nor_1331_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3)))
      OR (NOT (fsm_output(9))) OR (fsm_output(2)) OR (fsm_output(10)));
  nor_1332_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(3)) OR (fsm_output(9))
      OR (fsm_output(2)) OR (NOT (fsm_output(10))));
  mux_1332_nl <= MUX_s_1_2_2(nor_1331_nl, nor_1332_nl, fsm_output(1));
  mux_1336_nl <= MUX_s_1_2_2(mux_1335_nl, mux_1332_nl, fsm_output(0));
  mux_1338_nl <= MUX_s_1_2_2(mux_1337_nl, mux_1336_nl, fsm_output(6));
  mux_1348_nl <= MUX_s_1_2_2(mux_1347_nl, mux_1338_nl, fsm_output(8));
  vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_1363_nl, mux_1348_nl,
      fsm_output(4));
  or_1060_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR
      (NOT (fsm_output(9))) OR (NOT (fsm_output(5))) OR (fsm_output(10));
  or_1059_nl <= (NOT (fsm_output(9))) OR (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0100")) OR (NOT (fsm_output(10)));
  mux_1390_nl <= MUX_s_1_2_2(or_1060_nl, or_1059_nl, fsm_output(7));
  or_1057_nl <= CONV_SL_1_1(VEC_LOOP_j_sva_11_0(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01"))
      OR (NOT (fsm_output(7))) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (fsm_output(9)) OR (fsm_output(5)) OR (fsm_output(10));
  mux_1391_nl <= MUX_s_1_2_2(mux_1390_nl, or_1057_nl, fsm_output(2));
  nor_1287_nl <= NOT((fsm_output(6)) OR (fsm_output(4)) OR mux_1391_nl);
  nor_1288_nl <= NOT((fsm_output(6)) OR (fsm_output(4)) OR (NOT (fsm_output(2)))
      OR (fsm_output(7)) OR (fsm_output(9)) OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0100")) OR (NOT (fsm_output(10))));
  mux_1392_nl <= MUX_s_1_2_2(nor_1287_nl, nor_1288_nl, fsm_output(8));
  nor_1289_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT (fsm_output(6))) OR (NOT (fsm_output(4))) OR (fsm_output(2)) OR (NOT
      (fsm_output(7))) OR (fsm_output(9)) OR not_tmp_248);
  nor_1290_nl <= NOT((fsm_output(4)) OR (fsm_output(2)) OR (fsm_output(7)) OR (NOT
      (fsm_output(9))) OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0100")) OR (fsm_output(10)));
  nor_1291_nl <= NOT((NOT (fsm_output(2))) OR (fsm_output(7)) OR (fsm_output(9))
      OR (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("0100")) OR (fsm_output(10)));
  nor_1292_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT (fsm_output(2))) OR (fsm_output(7)) OR (NOT (fsm_output(9))) OR (fsm_output(5))
      OR (fsm_output(10)));
  mux_1387_nl <= MUX_s_1_2_2(nor_1291_nl, nor_1292_nl, fsm_output(4));
  mux_1388_nl <= MUX_s_1_2_2(nor_1290_nl, mux_1387_nl, fsm_output(6));
  mux_1389_nl <= MUX_s_1_2_2(nor_1289_nl, mux_1388_nl, fsm_output(8));
  mux_1393_nl <= MUX_s_1_2_2(mux_1392_nl, mux_1389_nl, fsm_output(0));
  or_1048_nl <= (COMP_LOOP_acc_16_psp_sva(0)) OR (NOT (fsm_output(4))) OR (NOT (fsm_output(2)))
      OR (NOT (VEC_LOOP_j_sva_11_0(2))) OR (NOT (fsm_output(7))) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(5)))
      OR (fsm_output(10));
  or_1047_nl <= CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR (fsm_output(2)) OR (fsm_output(7)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR (fsm_output(9)) OR (fsm_output(5)) OR
      (NOT (fsm_output(10)));
  mux_1384_nl <= MUX_s_1_2_2(mux_tmp_1372, or_1047_nl, fsm_output(4));
  mux_1385_nl <= MUX_s_1_2_2(or_1048_nl, mux_1384_nl, fsm_output(6));
  and_610_nl <= (fsm_output(8)) AND (NOT mux_1385_nl);
  or_1044_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(7))) OR (NOT (fsm_output(9)))
      OR (fsm_output(5)) OR (NOT (fsm_output(10)));
  or_1042_nl <= (fsm_output(7)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(5)))
      OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT (fsm_output(10)));
  mux_1381_nl <= MUX_s_1_2_2(or_1042_nl, or_tmp_974, fsm_output(2));
  mux_1382_nl <= MUX_s_1_2_2(or_1044_nl, mux_1381_nl, fsm_output(4));
  nor_1293_nl <= NOT((fsm_output(6)) OR mux_1382_nl);
  nor_1294_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(6)) OR (NOT (fsm_output(4))) OR (fsm_output(2)) OR (NOT (fsm_output(7)))
      OR (fsm_output(9)) OR (NOT (fsm_output(5))) OR (fsm_output(10)));
  mux_1383_nl <= MUX_s_1_2_2(nor_1293_nl, nor_1294_nl, fsm_output(8));
  mux_1386_nl <= MUX_s_1_2_2(and_610_nl, mux_1383_nl, fsm_output(0));
  mux_1394_nl <= MUX_s_1_2_2(mux_1393_nl, mux_1386_nl, fsm_output(3));
  or_1038_nl <= CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (NOT (fsm_output(2))) OR (fsm_output(7)) OR (VEC_LOOP_j_sva_11_0(0)) OR
      nand_337_cse;
  or_1036_nl <= (NOT (fsm_output(2))) OR (fsm_output(7)) OR (fsm_output(9)) OR (NOT
      (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT (fsm_output(10)));
  mux_1377_nl <= MUX_s_1_2_2(or_1038_nl, or_1036_nl, fsm_output(4));
  nor_1295_nl <= NOT((fsm_output(6)) OR mux_1377_nl);
  or_1032_nl <= (fsm_output(9)) OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0100")) OR (NOT (fsm_output(10)));
  mux_1375_nl <= MUX_s_1_2_2(or_591_cse, or_1032_nl, fsm_output(7));
  mux_1376_nl <= MUX_s_1_2_2(mux_1375_nl, or_tmp_974, or_1028_cse);
  nor_1296_nl <= NOT((NOT (fsm_output(6))) OR (NOT (fsm_output(4))) OR (fsm_output(2))
      OR mux_1376_nl);
  mux_1378_nl <= MUX_s_1_2_2(nor_1295_nl, nor_1296_nl, fsm_output(8));
  or_1025_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(7)) OR (fsm_output(9)) OR not_tmp_248;
  or_1023_nl <= (NOT (fsm_output(7))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0100")) OR (NOT (fsm_output(9))) OR (fsm_output(5))
      OR (fsm_output(10));
  mux_1373_nl <= MUX_s_1_2_2(or_1025_nl, or_1023_nl, fsm_output(2));
  mux_1374_nl <= MUX_s_1_2_2(mux_1373_nl, mux_tmp_1372, fsm_output(4));
  nor_1297_nl <= NOT((fsm_output(8)) OR (fsm_output(6)) OR mux_1374_nl);
  mux_1379_nl <= MUX_s_1_2_2(mux_1378_nl, nor_1297_nl, fsm_output(0));
  or_1018_nl <= CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (fsm_output(2)) OR (NOT (fsm_output(7))) OR (VEC_LOOP_j_sva_11_0(0)) OR
      (fsm_output(9)) OR (fsm_output(5)) OR (NOT (fsm_output(10)));
  or_1016_nl <= (fsm_output(2)) OR (NOT (fsm_output(7))) OR (NOT (fsm_output(9)))
      OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("0100")) OR (fsm_output(10));
  mux_1369_nl <= MUX_s_1_2_2(or_1018_nl, or_1016_nl, fsm_output(4));
  or_1015_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(7))) OR (VEC_LOOP_j_sva_11_0(0))
      OR (NOT (fsm_output(9))) OR (NOT (fsm_output(5))) OR (fsm_output(10));
  or_1014_nl <= (NOT (fsm_output(2))) OR (NOT (fsm_output(7))) OR (fsm_output(9))
      OR (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("0100")) OR (fsm_output(10));
  mux_1368_nl <= MUX_s_1_2_2(or_1015_nl, or_1014_nl, fsm_output(4));
  mux_1370_nl <= MUX_s_1_2_2(mux_1369_nl, mux_1368_nl, fsm_output(6));
  nor_1298_nl <= NOT((fsm_output(8)) OR mux_1370_nl);
  nor_1299_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT (fsm_output(6))) OR (fsm_output(4)) OR (fsm_output(2)) OR (NOT (fsm_output(7)))
      OR (fsm_output(9)) OR (NOT (fsm_output(5))) OR (fsm_output(10)));
  nor_1300_nl <= NOT((NOT (fsm_output(4))) OR (NOT (fsm_output(2))) OR (NOT (fsm_output(7)))
      OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(9)) OR not_tmp_248);
  or_1009_nl <= (fsm_output(7)) OR (fsm_output(9)) OR (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0100")) OR (NOT (fsm_output(10)));
  or_1007_nl <= (NOT (fsm_output(7))) OR (NOT (fsm_output(9))) OR (fsm_output(5))
      OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(10));
  mux_1365_nl <= MUX_s_1_2_2(or_1009_nl, or_1007_nl, fsm_output(2));
  nor_1301_nl <= NOT((fsm_output(4)) OR mux_1365_nl);
  mux_1366_nl <= MUX_s_1_2_2(nor_1300_nl, nor_1301_nl, fsm_output(6));
  mux_1367_nl <= MUX_s_1_2_2(nor_1299_nl, mux_1366_nl, fsm_output(8));
  mux_1371_nl <= MUX_s_1_2_2(nor_1298_nl, mux_1367_nl, fsm_output(0));
  mux_1380_nl <= MUX_s_1_2_2(mux_1379_nl, mux_1371_nl, fsm_output(3));
  vec_rsc_0_4_i_wea_d_pff <= MUX_s_1_2_2(mux_1394_nl, mux_1380_nl, fsm_output(1));
  or_1116_nl <= (NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(2))) OR (fsm_output(10));
  or_1115_nl <= (fsm_output(7)) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(2)) OR (NOT (fsm_output(10)));
  mux_1425_nl <= MUX_s_1_2_2(or_1116_nl, or_1115_nl, fsm_output(5));
  nor_1256_nl <= NOT((fsm_output(1)) OR mux_1425_nl);
  nor_1257_nl <= NOT((fsm_output(5)) OR (NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0100")) OR (fsm_output(3)) OR (fsm_output(9))
      OR (fsm_output(2)) OR (fsm_output(10)));
  nor_1258_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT (fsm_output(7))) OR (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_253);
  nor_1259_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(7)) OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (fsm_output(2))
      OR (NOT (fsm_output(10))));
  mux_1423_nl <= MUX_s_1_2_2(nor_1258_nl, nor_1259_nl, fsm_output(5));
  mux_1424_nl <= MUX_s_1_2_2(nor_1257_nl, mux_1423_nl, fsm_output(1));
  mux_1426_nl <= MUX_s_1_2_2(nor_1256_nl, mux_1424_nl, fsm_output(0));
  and_607_nl <= (fsm_output(6)) AND mux_1426_nl;
  nor_1260_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR (fsm_output(2)) OR (fsm_output(10)));
  nor_1262_nl <= NOT((fsm_output(7)) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR not_tmp_253);
  mux_1418_nl <= MUX_s_1_2_2(nor_1445_cse, nor_1262_nl, fsm_output(5));
  nor_1263_nl <= NOT((NOT (fsm_output(5))) OR (fsm_output(7)) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0100")) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR not_tmp_253);
  or_1102_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm);
  mux_1419_nl <= MUX_s_1_2_2(mux_1418_nl, nor_1263_nl, or_1102_nl);
  mux_1420_nl <= MUX_s_1_2_2(nor_1260_nl, mux_1419_nl, fsm_output(1));
  nor_1264_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR
      (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_253);
  nor_1265_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (NOT
      (fsm_output(2))) OR (fsm_output(10)));
  nor_1266_nl <= NOT((fsm_output(7)) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9))) OR (fsm_output(2)) OR (fsm_output(10)));
  mux_1416_nl <= MUX_s_1_2_2(nor_1265_nl, nor_1266_nl, fsm_output(5));
  mux_1417_nl <= MUX_s_1_2_2(nor_1264_nl, mux_1416_nl, fsm_output(1));
  mux_1421_nl <= MUX_s_1_2_2(mux_1420_nl, mux_1417_nl, fsm_output(0));
  nor_1267_nl <= NOT((NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (NOT (fsm_output(5)))
      OR (fsm_output(7)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR not_tmp_253);
  nor_1268_nl <= NOT((NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (NOT (fsm_output(5)))
      OR (fsm_output(7)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(3)) OR (fsm_output(9)) OR (NOT (fsm_output(2))) OR (fsm_output(10)));
  mux_1414_nl <= MUX_s_1_2_2(nor_1267_nl, nor_1268_nl, fsm_output(1));
  nor_1269_nl <= NOT((fsm_output(1)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO
      0)/=STD_LOGIC_VECTOR'("00")) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR mux_1413_cse);
  mux_1415_nl <= MUX_s_1_2_2(mux_1414_nl, nor_1269_nl, fsm_output(0));
  mux_1422_nl <= MUX_s_1_2_2(mux_1421_nl, mux_1415_nl, fsm_output(6));
  mux_1427_nl <= MUX_s_1_2_2(and_607_nl, mux_1422_nl, fsm_output(8));
  nor_1270_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (fsm_output(2))
      OR (fsm_output(10)));
  nor_1271_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(7)) OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(2)))
      OR (fsm_output(10)));
  mux_1408_nl <= MUX_s_1_2_2(nor_1270_nl, nor_1271_nl, fsm_output(5));
  and_608_nl <= COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm AND mux_1408_nl;
  nor_1272_nl <= NOT((NOT (fsm_output(7))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0100")) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR not_tmp_253);
  nor_1273_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(7)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9))) OR (fsm_output(2))
      OR (NOT (fsm_output(10))));
  mux_1407_nl <= MUX_s_1_2_2(nor_1272_nl, nor_1273_nl, fsm_output(5));
  and_609_nl <= COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm AND mux_1407_nl;
  mux_1409_nl <= MUX_s_1_2_2(and_608_nl, and_609_nl, fsm_output(1));
  nor_1274_nl <= NOT((VEC_LOOP_j_sva_11_0(3)) OR (VEC_LOOP_j_sva_11_0(1)) OR (VEC_LOOP_j_sva_11_0(0))
      OR (NOT (fsm_output(5))) OR (NOT (VEC_LOOP_j_sva_11_0(2))) OR (fsm_output(7))
      OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(2)) OR (fsm_output(10)));
  nor_1275_nl <= NOT((VEC_LOOP_j_sva_11_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR mux_1405_cse);
  mux_1406_nl <= MUX_s_1_2_2(nor_1274_nl, nor_1275_nl, fsm_output(1));
  mux_1410_nl <= MUX_s_1_2_2(mux_1409_nl, mux_1406_nl, fsm_output(0));
  nor_1276_nl <= NOT((NOT (fsm_output(1))) OR (fsm_output(5)) OR (fsm_output(7))
      OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100")) OR (NOT
      (fsm_output(3))) OR (fsm_output(9)) OR (fsm_output(2)) OR (fsm_output(10)));
  nor_1277_nl <= NOT((fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(3)))
      OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100")) OR (NOT
      (fsm_output(9))) OR (NOT (fsm_output(2))) OR (fsm_output(10)));
  nor_1278_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (VEC_LOOP_j_sva_11_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR
      (NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3))) OR
      (fsm_output(9)) OR (NOT (fsm_output(2))) OR (fsm_output(10)));
  mux_1403_nl <= MUX_s_1_2_2(nor_1277_nl, nor_1278_nl, fsm_output(1));
  mux_1404_nl <= MUX_s_1_2_2(nor_1276_nl, mux_1403_nl, fsm_output(0));
  mux_1411_nl <= MUX_s_1_2_2(mux_1410_nl, mux_1404_nl, fsm_output(6));
  nor_1279_nl <= NOT((NOT (fsm_output(1))) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(3)) OR (NOT (fsm_output(9)))
      OR (fsm_output(2)) OR (fsm_output(10)));
  nor_1280_nl <= NOT((fsm_output(1)) OR (fsm_output(5)) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0100")) OR (NOT (fsm_output(7))) OR (fsm_output(3))
      OR (fsm_output(9)) OR not_tmp_253);
  mux_1401_nl <= MUX_s_1_2_2(nor_1279_nl, nor_1280_nl, fsm_output(0));
  nor_1281_nl <= NOT((NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0100")) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR not_tmp_253);
  nor_1282_nl <= NOT((NOT (fsm_output(7))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0100")) OR (fsm_output(3)) OR (NOT (fsm_output(9)))
      OR (fsm_output(2)) OR (fsm_output(10)));
  nor_1283_nl <= NOT((NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR not_tmp_253);
  mux_1397_nl <= MUX_s_1_2_2(nor_1282_nl, nor_1283_nl, fsm_output(5));
  mux_1398_nl <= MUX_s_1_2_2(nor_1281_nl, mux_1397_nl, COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm);
  nor_1284_nl <= NOT((NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0100")) OR (fsm_output(3)) OR (fsm_output(9))
      OR (NOT (fsm_output(2))) OR (fsm_output(10)));
  mux_1399_nl <= MUX_s_1_2_2(mux_1398_nl, nor_1284_nl, fsm_output(1));
  nor_1285_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3)))
      OR (NOT (fsm_output(9))) OR (fsm_output(2)) OR (fsm_output(10)));
  nor_1286_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (VEC_LOOP_j_sva_11_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR
      (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(3)) OR (fsm_output(9))
      OR (fsm_output(2)) OR (NOT (fsm_output(10))));
  mux_1396_nl <= MUX_s_1_2_2(nor_1285_nl, nor_1286_nl, fsm_output(1));
  mux_1400_nl <= MUX_s_1_2_2(mux_1399_nl, mux_1396_nl, fsm_output(0));
  mux_1402_nl <= MUX_s_1_2_2(mux_1401_nl, mux_1400_nl, fsm_output(6));
  mux_1412_nl <= MUX_s_1_2_2(mux_1411_nl, mux_1402_nl, fsm_output(8));
  vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_1427_nl, mux_1412_nl,
      fsm_output(4));
  or_1171_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR
      (NOT (fsm_output(9))) OR (NOT (fsm_output(5))) OR (fsm_output(10));
  nand_403_nl <= NOT((fsm_output(9)) AND (fsm_output(5)) AND CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)=STD_LOGIC_VECTOR'("0101")) AND (fsm_output(10)));
  mux_1454_nl <= MUX_s_1_2_2(or_1171_nl, nand_403_nl, fsm_output(7));
  or_1168_nl <= CONV_SL_1_1(VEC_LOOP_j_sva_11_0(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01"))
      OR (NOT (fsm_output(7))) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR (fsm_output(9)) OR (fsm_output(5)) OR (fsm_output(10));
  mux_1455_nl <= MUX_s_1_2_2(mux_1454_nl, or_1168_nl, fsm_output(2));
  nor_1241_nl <= NOT((fsm_output(6)) OR (fsm_output(4)) OR mux_1455_nl);
  nor_1242_nl <= NOT((fsm_output(6)) OR (fsm_output(4)) OR (NOT (fsm_output(2)))
      OR (fsm_output(7)) OR (fsm_output(9)) OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0101")) OR (NOT (fsm_output(10))));
  mux_1456_nl <= MUX_s_1_2_2(nor_1241_nl, nor_1242_nl, fsm_output(8));
  nor_1243_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT (fsm_output(6))) OR (NOT (fsm_output(4))) OR (fsm_output(2)) OR (NOT
      (fsm_output(7))) OR (fsm_output(9)) OR not_tmp_248);
  nor_1244_nl <= NOT((fsm_output(4)) OR (fsm_output(2)) OR (fsm_output(7)) OR (NOT
      (fsm_output(9))) OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0101")) OR (fsm_output(10)));
  nor_1245_nl <= NOT((NOT (fsm_output(2))) OR (fsm_output(7)) OR (fsm_output(9))
      OR (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("0101")) OR (fsm_output(10)));
  nor_1246_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT (fsm_output(2))) OR (fsm_output(7)) OR (NOT (fsm_output(9))) OR (fsm_output(5))
      OR (fsm_output(10)));
  mux_1451_nl <= MUX_s_1_2_2(nor_1245_nl, nor_1246_nl, fsm_output(4));
  mux_1452_nl <= MUX_s_1_2_2(nor_1244_nl, mux_1451_nl, fsm_output(6));
  mux_1453_nl <= MUX_s_1_2_2(nor_1243_nl, mux_1452_nl, fsm_output(8));
  mux_1457_nl <= MUX_s_1_2_2(mux_1456_nl, mux_1453_nl, fsm_output(0));
  nand_318_nl <= NOT((NOT (COMP_LOOP_acc_16_psp_sva(0))) AND (fsm_output(4)) AND
      (fsm_output(2)) AND (VEC_LOOP_j_sva_11_0(2)) AND (fsm_output(7)) AND CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1
      DOWNTO 0)=STD_LOGIC_VECTOR'("01")) AND (fsm_output(9)) AND (fsm_output(5))
      AND (NOT (fsm_output(10))));
  or_1158_nl <= CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR (fsm_output(2)) OR (fsm_output(7)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR (fsm_output(9)) OR (fsm_output(5)) OR
      (NOT (fsm_output(10)));
  mux_1448_nl <= MUX_s_1_2_2(mux_tmp_1436, or_1158_nl, fsm_output(4));
  mux_1449_nl <= MUX_s_1_2_2(nand_318_nl, mux_1448_nl, fsm_output(6));
  and_606_nl <= (fsm_output(8)) AND (NOT mux_1449_nl);
  or_1155_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(7))) OR (NOT (fsm_output(9)))
      OR (fsm_output(5)) OR (NOT (fsm_output(10)));
  or_1153_nl <= (fsm_output(7)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(5)))
      OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT (fsm_output(10)));
  mux_1445_nl <= MUX_s_1_2_2(or_1153_nl, or_tmp_1085, fsm_output(2));
  mux_1446_nl <= MUX_s_1_2_2(or_1155_nl, mux_1445_nl, fsm_output(4));
  nor_1247_nl <= NOT((fsm_output(6)) OR mux_1446_nl);
  nor_1248_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(6)) OR (NOT (fsm_output(4))) OR (fsm_output(2)) OR (NOT (fsm_output(7)))
      OR (fsm_output(9)) OR (NOT (fsm_output(5))) OR (fsm_output(10)));
  mux_1447_nl <= MUX_s_1_2_2(nor_1247_nl, nor_1248_nl, fsm_output(8));
  mux_1450_nl <= MUX_s_1_2_2(and_606_nl, mux_1447_nl, fsm_output(0));
  mux_1458_nl <= MUX_s_1_2_2(mux_1457_nl, mux_1450_nl, fsm_output(3));
  or_1149_nl <= CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (NOT (fsm_output(2))) OR (fsm_output(7)) OR nand_334_cse;
  or_1147_nl <= (NOT (fsm_output(2))) OR (fsm_output(7)) OR (fsm_output(9)) OR (NOT
      (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT (fsm_output(10)));
  mux_1441_nl <= MUX_s_1_2_2(or_1149_nl, or_1147_nl, fsm_output(4));
  nor_1249_nl <= NOT((fsm_output(6)) OR mux_1441_nl);
  or_1143_nl <= (fsm_output(9)) OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0101")) OR (NOT (fsm_output(10)));
  mux_1439_nl <= MUX_s_1_2_2(or_702_cse, or_1143_nl, fsm_output(7));
  mux_1440_nl <= MUX_s_1_2_2(mux_1439_nl, or_tmp_1085, or_1028_cse);
  nor_1250_nl <= NOT((NOT (fsm_output(6))) OR (NOT (fsm_output(4))) OR (fsm_output(2))
      OR mux_1440_nl);
  mux_1442_nl <= MUX_s_1_2_2(nor_1249_nl, nor_1250_nl, fsm_output(8));
  or_1136_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(7)) OR (fsm_output(9)) OR not_tmp_248;
  or_1134_nl <= (NOT (fsm_output(7))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0101")) OR (NOT (fsm_output(9))) OR (fsm_output(5))
      OR (fsm_output(10));
  mux_1437_nl <= MUX_s_1_2_2(or_1136_nl, or_1134_nl, fsm_output(2));
  mux_1438_nl <= MUX_s_1_2_2(mux_1437_nl, mux_tmp_1436, fsm_output(4));
  nor_1251_nl <= NOT((fsm_output(8)) OR (fsm_output(6)) OR mux_1438_nl);
  mux_1443_nl <= MUX_s_1_2_2(mux_1442_nl, nor_1251_nl, fsm_output(0));
  or_1129_nl <= CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (fsm_output(2)) OR (NOT (fsm_output(7))) OR (NOT (VEC_LOOP_j_sva_11_0(0)))
      OR (fsm_output(9)) OR (fsm_output(5)) OR (NOT (fsm_output(10)));
  or_1127_nl <= (fsm_output(2)) OR (NOT (fsm_output(7))) OR (NOT (fsm_output(9)))
      OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("0101")) OR (fsm_output(10));
  mux_1433_nl <= MUX_s_1_2_2(or_1129_nl, or_1127_nl, fsm_output(4));
  or_1126_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(7))) OR (NOT (VEC_LOOP_j_sva_11_0(0)))
      OR (NOT (fsm_output(9))) OR (NOT (fsm_output(5))) OR (fsm_output(10));
  or_1125_nl <= (NOT (fsm_output(2))) OR (NOT (fsm_output(7))) OR (fsm_output(9))
      OR (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("0101")) OR (fsm_output(10));
  mux_1432_nl <= MUX_s_1_2_2(or_1126_nl, or_1125_nl, fsm_output(4));
  mux_1434_nl <= MUX_s_1_2_2(mux_1433_nl, mux_1432_nl, fsm_output(6));
  nor_1252_nl <= NOT((fsm_output(8)) OR mux_1434_nl);
  nor_1253_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT (fsm_output(6))) OR (fsm_output(4)) OR (fsm_output(2)) OR (NOT (fsm_output(7)))
      OR (fsm_output(9)) OR (NOT (fsm_output(5))) OR (fsm_output(10)));
  nor_1254_nl <= NOT((NOT (fsm_output(4))) OR (NOT (fsm_output(2))) OR (NOT (fsm_output(7)))
      OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(9)) OR not_tmp_248);
  or_1120_nl <= (fsm_output(7)) OR (fsm_output(9)) OR (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0101")) OR (NOT (fsm_output(10)));
  or_1118_nl <= (NOT (fsm_output(7))) OR (NOT (fsm_output(9))) OR (fsm_output(5))
      OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(10));
  mux_1429_nl <= MUX_s_1_2_2(or_1120_nl, or_1118_nl, fsm_output(2));
  nor_1255_nl <= NOT((fsm_output(4)) OR mux_1429_nl);
  mux_1430_nl <= MUX_s_1_2_2(nor_1254_nl, nor_1255_nl, fsm_output(6));
  mux_1431_nl <= MUX_s_1_2_2(nor_1253_nl, mux_1430_nl, fsm_output(8));
  mux_1435_nl <= MUX_s_1_2_2(nor_1252_nl, mux_1431_nl, fsm_output(0));
  mux_1444_nl <= MUX_s_1_2_2(mux_1443_nl, mux_1435_nl, fsm_output(3));
  vec_rsc_0_5_i_wea_d_pff <= MUX_s_1_2_2(mux_1458_nl, mux_1444_nl, fsm_output(1));
  or_1227_nl <= (NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(2))) OR (fsm_output(10));
  or_1226_nl <= (fsm_output(7)) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(2)) OR (NOT (fsm_output(10)));
  mux_1489_nl <= MUX_s_1_2_2(or_1227_nl, or_1226_nl, fsm_output(5));
  nor_1210_nl <= NOT((fsm_output(1)) OR mux_1489_nl);
  nor_1211_nl <= NOT((fsm_output(5)) OR (NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0101")) OR (fsm_output(3)) OR (fsm_output(9))
      OR (fsm_output(2)) OR (fsm_output(10)));
  nor_1212_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT (fsm_output(7))) OR (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_253);
  nor_1213_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(7)) OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (fsm_output(2))
      OR (NOT (fsm_output(10))));
  mux_1487_nl <= MUX_s_1_2_2(nor_1212_nl, nor_1213_nl, fsm_output(5));
  mux_1488_nl <= MUX_s_1_2_2(nor_1211_nl, mux_1487_nl, fsm_output(1));
  mux_1490_nl <= MUX_s_1_2_2(nor_1210_nl, mux_1488_nl, fsm_output(0));
  and_603_nl <= (fsm_output(6)) AND mux_1490_nl;
  nor_1214_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR (fsm_output(2)) OR (fsm_output(10)));
  nor_1216_nl <= NOT((fsm_output(7)) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR not_tmp_253);
  mux_1482_nl <= MUX_s_1_2_2(nor_1445_cse, nor_1216_nl, fsm_output(5));
  nor_1217_nl <= NOT((NOT (fsm_output(5))) OR (fsm_output(7)) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0101")) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR not_tmp_253);
  or_1213_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm);
  mux_1483_nl <= MUX_s_1_2_2(mux_1482_nl, nor_1217_nl, or_1213_nl);
  mux_1484_nl <= MUX_s_1_2_2(nor_1214_nl, mux_1483_nl, fsm_output(1));
  nor_1218_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR
      (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_253);
  nor_1219_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (NOT
      (fsm_output(2))) OR (fsm_output(10)));
  nor_1220_nl <= NOT((fsm_output(7)) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9))) OR (fsm_output(2)) OR (fsm_output(10)));
  mux_1480_nl <= MUX_s_1_2_2(nor_1219_nl, nor_1220_nl, fsm_output(5));
  mux_1481_nl <= MUX_s_1_2_2(nor_1218_nl, mux_1480_nl, fsm_output(1));
  mux_1485_nl <= MUX_s_1_2_2(mux_1484_nl, mux_1481_nl, fsm_output(0));
  nor_1221_nl <= NOT((NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (NOT (fsm_output(5)))
      OR (fsm_output(7)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR not_tmp_253);
  nor_1222_nl <= NOT((NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (NOT (fsm_output(5)))
      OR (fsm_output(7)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(3)) OR (fsm_output(9)) OR (NOT (fsm_output(2))) OR (fsm_output(10)));
  mux_1478_nl <= MUX_s_1_2_2(nor_1221_nl, nor_1222_nl, fsm_output(1));
  nor_1223_nl <= NOT((fsm_output(1)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO
      0)/=STD_LOGIC_VECTOR'("01")) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR mux_1413_cse);
  mux_1479_nl <= MUX_s_1_2_2(mux_1478_nl, nor_1223_nl, fsm_output(0));
  mux_1486_nl <= MUX_s_1_2_2(mux_1485_nl, mux_1479_nl, fsm_output(6));
  mux_1491_nl <= MUX_s_1_2_2(and_603_nl, mux_1486_nl, fsm_output(8));
  nor_1224_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (fsm_output(2))
      OR (fsm_output(10)));
  nor_1225_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(7)) OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(2)))
      OR (fsm_output(10)));
  mux_1472_nl <= MUX_s_1_2_2(nor_1224_nl, nor_1225_nl, fsm_output(5));
  and_604_nl <= COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm AND mux_1472_nl;
  nor_1226_nl <= NOT((NOT (fsm_output(7))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0101")) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR not_tmp_253);
  nor_1227_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(7)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9))) OR (fsm_output(2))
      OR (NOT (fsm_output(10))));
  mux_1471_nl <= MUX_s_1_2_2(nor_1226_nl, nor_1227_nl, fsm_output(5));
  and_605_nl <= COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm AND mux_1471_nl;
  mux_1473_nl <= MUX_s_1_2_2(and_604_nl, and_605_nl, fsm_output(1));
  nor_1228_nl <= NOT((VEC_LOOP_j_sva_11_0(3)) OR (VEC_LOOP_j_sva_11_0(1)) OR (NOT
      (VEC_LOOP_j_sva_11_0(0))) OR (NOT (fsm_output(5))) OR (NOT (VEC_LOOP_j_sva_11_0(2)))
      OR (fsm_output(7)) OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(2))
      OR (fsm_output(10)));
  nor_1229_nl <= NOT(nand_332_cse OR mux_1405_cse);
  mux_1470_nl <= MUX_s_1_2_2(nor_1228_nl, nor_1229_nl, fsm_output(1));
  mux_1474_nl <= MUX_s_1_2_2(mux_1473_nl, mux_1470_nl, fsm_output(0));
  nor_1230_nl <= NOT((NOT (fsm_output(1))) OR (fsm_output(5)) OR (fsm_output(7))
      OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101")) OR (NOT
      (fsm_output(3))) OR (fsm_output(9)) OR (fsm_output(2)) OR (fsm_output(10)));
  nor_1231_nl <= NOT((fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(3)))
      OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101")) OR (NOT
      (fsm_output(9))) OR (NOT (fsm_output(2))) OR (fsm_output(10)));
  nor_1232_nl <= NOT((NOT (VEC_LOOP_j_sva_11_0(0))) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (NOT
      (fsm_output(2))) OR (fsm_output(10)));
  mux_1467_nl <= MUX_s_1_2_2(nor_1231_nl, nor_1232_nl, fsm_output(1));
  mux_1468_nl <= MUX_s_1_2_2(nor_1230_nl, mux_1467_nl, fsm_output(0));
  mux_1475_nl <= MUX_s_1_2_2(mux_1474_nl, mux_1468_nl, fsm_output(6));
  nor_1233_nl <= NOT((NOT (fsm_output(1))) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(3)) OR (NOT (fsm_output(9)))
      OR (fsm_output(2)) OR (fsm_output(10)));
  nor_1234_nl <= NOT((fsm_output(1)) OR (fsm_output(5)) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0101")) OR (NOT (fsm_output(7))) OR (fsm_output(3))
      OR (fsm_output(9)) OR not_tmp_253);
  mux_1465_nl <= MUX_s_1_2_2(nor_1233_nl, nor_1234_nl, fsm_output(0));
  nor_1235_nl <= NOT((NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0101")) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR not_tmp_253);
  nor_1236_nl <= NOT((NOT (fsm_output(7))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0101")) OR (fsm_output(3)) OR (NOT (fsm_output(9)))
      OR (fsm_output(2)) OR (fsm_output(10)));
  nor_1237_nl <= NOT((NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR not_tmp_253);
  mux_1461_nl <= MUX_s_1_2_2(nor_1236_nl, nor_1237_nl, fsm_output(5));
  mux_1462_nl <= MUX_s_1_2_2(nor_1235_nl, mux_1461_nl, COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm);
  nor_1238_nl <= NOT((NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0101")) OR (fsm_output(3)) OR (fsm_output(9))
      OR (NOT (fsm_output(2))) OR (fsm_output(10)));
  mux_1463_nl <= MUX_s_1_2_2(mux_1462_nl, nor_1238_nl, fsm_output(1));
  nor_1239_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3)))
      OR (NOT (fsm_output(9))) OR (fsm_output(2)) OR (fsm_output(10)));
  nor_1240_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(3)) OR (fsm_output(9))
      OR (fsm_output(2)) OR (NOT (fsm_output(10))));
  mux_1460_nl <= MUX_s_1_2_2(nor_1239_nl, nor_1240_nl, fsm_output(1));
  mux_1464_nl <= MUX_s_1_2_2(mux_1463_nl, mux_1460_nl, fsm_output(0));
  mux_1466_nl <= MUX_s_1_2_2(mux_1465_nl, mux_1464_nl, fsm_output(6));
  mux_1476_nl <= MUX_s_1_2_2(mux_1475_nl, mux_1466_nl, fsm_output(8));
  vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_1491_nl, mux_1476_nl,
      fsm_output(4));
  or_1281_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR
      (NOT (fsm_output(9))) OR (NOT (fsm_output(5))) OR (fsm_output(10));
  nand_402_nl <= NOT((fsm_output(9)) AND (fsm_output(5)) AND CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)=STD_LOGIC_VECTOR'("0110")) AND (fsm_output(10)));
  mux_1518_nl <= MUX_s_1_2_2(or_1281_nl, nand_402_nl, fsm_output(7));
  or_1278_nl <= CONV_SL_1_1(VEC_LOOP_j_sva_11_0(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01"))
      OR (NOT (fsm_output(7))) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (fsm_output(9)) OR (fsm_output(5)) OR (fsm_output(10));
  mux_1519_nl <= MUX_s_1_2_2(mux_1518_nl, or_1278_nl, fsm_output(2));
  nor_1195_nl <= NOT((fsm_output(6)) OR (fsm_output(4)) OR mux_1519_nl);
  nor_1196_nl <= NOT((fsm_output(6)) OR (fsm_output(4)) OR (NOT (fsm_output(2)))
      OR (fsm_output(7)) OR (fsm_output(9)) OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0110")) OR (NOT (fsm_output(10))));
  mux_1520_nl <= MUX_s_1_2_2(nor_1195_nl, nor_1196_nl, fsm_output(8));
  nor_1197_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT (fsm_output(6))) OR (NOT (fsm_output(4))) OR (fsm_output(2)) OR (NOT
      (fsm_output(7))) OR (fsm_output(9)) OR not_tmp_248);
  nor_1198_nl <= NOT((fsm_output(4)) OR (fsm_output(2)) OR (fsm_output(7)) OR (NOT
      (fsm_output(9))) OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0110")) OR (fsm_output(10)));
  nor_1199_nl <= NOT((NOT (fsm_output(2))) OR (fsm_output(7)) OR (fsm_output(9))
      OR (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("0110")) OR (fsm_output(10)));
  nor_1200_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT (fsm_output(2))) OR (fsm_output(7)) OR (NOT (fsm_output(9))) OR (fsm_output(5))
      OR (fsm_output(10)));
  mux_1515_nl <= MUX_s_1_2_2(nor_1199_nl, nor_1200_nl, fsm_output(4));
  mux_1516_nl <= MUX_s_1_2_2(nor_1198_nl, mux_1515_nl, fsm_output(6));
  mux_1517_nl <= MUX_s_1_2_2(nor_1197_nl, mux_1516_nl, fsm_output(8));
  mux_1521_nl <= MUX_s_1_2_2(mux_1520_nl, mux_1517_nl, fsm_output(0));
  nand_313_nl <= NOT((NOT (COMP_LOOP_acc_16_psp_sva(0))) AND (fsm_output(4)) AND
      (fsm_output(2)) AND (VEC_LOOP_j_sva_11_0(2)) AND (fsm_output(7)) AND CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1
      DOWNTO 0)=STD_LOGIC_VECTOR'("10")) AND (fsm_output(9)) AND (fsm_output(5))
      AND (NOT (fsm_output(10))));
  or_1268_nl <= CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR (fsm_output(2)) OR (fsm_output(7)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR (fsm_output(9)) OR (fsm_output(5)) OR
      (NOT (fsm_output(10)));
  mux_1512_nl <= MUX_s_1_2_2(mux_tmp_1500, or_1268_nl, fsm_output(4));
  mux_1513_nl <= MUX_s_1_2_2(nand_313_nl, mux_1512_nl, fsm_output(6));
  and_602_nl <= (fsm_output(8)) AND (NOT mux_1513_nl);
  or_1265_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(7))) OR (NOT (fsm_output(9)))
      OR (fsm_output(5)) OR (NOT (fsm_output(10)));
  or_1263_nl <= (fsm_output(7)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(5)))
      OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT (fsm_output(10)));
  mux_1509_nl <= MUX_s_1_2_2(or_1263_nl, or_tmp_1198, fsm_output(2));
  mux_1510_nl <= MUX_s_1_2_2(or_1265_nl, mux_1509_nl, fsm_output(4));
  nor_1201_nl <= NOT((fsm_output(6)) OR mux_1510_nl);
  nor_1202_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(6)) OR (NOT (fsm_output(4))) OR (fsm_output(2)) OR (NOT (fsm_output(7)))
      OR (fsm_output(9)) OR (NOT (fsm_output(5))) OR (fsm_output(10)));
  mux_1511_nl <= MUX_s_1_2_2(nor_1201_nl, nor_1202_nl, fsm_output(8));
  mux_1514_nl <= MUX_s_1_2_2(and_602_nl, mux_1511_nl, fsm_output(0));
  mux_1522_nl <= MUX_s_1_2_2(mux_1521_nl, mux_1514_nl, fsm_output(3));
  or_1259_nl <= CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (NOT (fsm_output(2))) OR (fsm_output(7)) OR (VEC_LOOP_j_sva_11_0(0)) OR
      nand_337_cse;
  or_1257_nl <= (NOT (fsm_output(2))) OR (fsm_output(7)) OR (fsm_output(9)) OR (NOT
      (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT (fsm_output(10)));
  mux_1505_nl <= MUX_s_1_2_2(or_1259_nl, or_1257_nl, fsm_output(4));
  nor_1203_nl <= NOT((fsm_output(6)) OR mux_1505_nl);
  or_1251_nl <= (fsm_output(9)) OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0110")) OR (NOT (fsm_output(10)));
  mux_1503_nl <= MUX_s_1_2_2(or_591_cse, or_1251_nl, fsm_output(7));
  mux_1504_nl <= MUX_s_1_2_2(or_tmp_1198, mux_1503_nl, nor_223_cse);
  nor_1204_nl <= NOT((NOT (fsm_output(6))) OR (NOT (fsm_output(4))) OR (fsm_output(2))
      OR mux_1504_nl);
  mux_1506_nl <= MUX_s_1_2_2(nor_1203_nl, nor_1204_nl, fsm_output(8));
  or_1247_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(7)) OR (fsm_output(9)) OR not_tmp_248;
  or_1245_nl <= (NOT (fsm_output(7))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0110")) OR (NOT (fsm_output(9))) OR (fsm_output(5))
      OR (fsm_output(10));
  mux_1501_nl <= MUX_s_1_2_2(or_1247_nl, or_1245_nl, fsm_output(2));
  mux_1502_nl <= MUX_s_1_2_2(mux_1501_nl, mux_tmp_1500, fsm_output(4));
  nor_1205_nl <= NOT((fsm_output(8)) OR (fsm_output(6)) OR mux_1502_nl);
  mux_1507_nl <= MUX_s_1_2_2(mux_1506_nl, nor_1205_nl, fsm_output(0));
  or_1240_nl <= CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (fsm_output(2)) OR (NOT (fsm_output(7))) OR (VEC_LOOP_j_sva_11_0(0)) OR
      (fsm_output(9)) OR (fsm_output(5)) OR (NOT (fsm_output(10)));
  or_1238_nl <= (fsm_output(2)) OR (NOT (fsm_output(7))) OR (NOT (fsm_output(9)))
      OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("0110")) OR (fsm_output(10));
  mux_1497_nl <= MUX_s_1_2_2(or_1240_nl, or_1238_nl, fsm_output(4));
  or_1237_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(7))) OR (VEC_LOOP_j_sva_11_0(0))
      OR (NOT (fsm_output(9))) OR (NOT (fsm_output(5))) OR (fsm_output(10));
  or_1236_nl <= (NOT (fsm_output(2))) OR (NOT (fsm_output(7))) OR (fsm_output(9))
      OR (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("0110")) OR (fsm_output(10));
  mux_1496_nl <= MUX_s_1_2_2(or_1237_nl, or_1236_nl, fsm_output(4));
  mux_1498_nl <= MUX_s_1_2_2(mux_1497_nl, mux_1496_nl, fsm_output(6));
  nor_1206_nl <= NOT((fsm_output(8)) OR mux_1498_nl);
  nor_1207_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT (fsm_output(6))) OR (fsm_output(4)) OR (fsm_output(2)) OR (NOT (fsm_output(7)))
      OR (fsm_output(9)) OR (NOT (fsm_output(5))) OR (fsm_output(10)));
  nor_1208_nl <= NOT((NOT (fsm_output(4))) OR (NOT (fsm_output(2))) OR (NOT (fsm_output(7)))
      OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(9)) OR not_tmp_248);
  or_1231_nl <= (fsm_output(7)) OR (fsm_output(9)) OR (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0110")) OR (NOT (fsm_output(10)));
  or_1229_nl <= (NOT (fsm_output(7))) OR (NOT (fsm_output(9))) OR (fsm_output(5))
      OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(10));
  mux_1493_nl <= MUX_s_1_2_2(or_1231_nl, or_1229_nl, fsm_output(2));
  nor_1209_nl <= NOT((fsm_output(4)) OR mux_1493_nl);
  mux_1494_nl <= MUX_s_1_2_2(nor_1208_nl, nor_1209_nl, fsm_output(6));
  mux_1495_nl <= MUX_s_1_2_2(nor_1207_nl, mux_1494_nl, fsm_output(8));
  mux_1499_nl <= MUX_s_1_2_2(nor_1206_nl, mux_1495_nl, fsm_output(0));
  mux_1508_nl <= MUX_s_1_2_2(mux_1507_nl, mux_1499_nl, fsm_output(3));
  vec_rsc_0_6_i_wea_d_pff <= MUX_s_1_2_2(mux_1522_nl, mux_1508_nl, fsm_output(1));
  or_1337_nl <= (NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(2))) OR (fsm_output(10));
  or_1336_nl <= (fsm_output(7)) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(2)) OR (NOT (fsm_output(10)));
  mux_1553_nl <= MUX_s_1_2_2(or_1337_nl, or_1336_nl, fsm_output(5));
  nor_1164_nl <= NOT((fsm_output(1)) OR mux_1553_nl);
  nor_1165_nl <= NOT((fsm_output(5)) OR (NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0110")) OR (fsm_output(3)) OR (fsm_output(9))
      OR (fsm_output(2)) OR (fsm_output(10)));
  nor_1166_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT (fsm_output(7))) OR (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_253);
  nor_1167_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(7)) OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (fsm_output(2))
      OR (NOT (fsm_output(10))));
  mux_1551_nl <= MUX_s_1_2_2(nor_1166_nl, nor_1167_nl, fsm_output(5));
  mux_1552_nl <= MUX_s_1_2_2(nor_1165_nl, mux_1551_nl, fsm_output(1));
  mux_1554_nl <= MUX_s_1_2_2(nor_1164_nl, mux_1552_nl, fsm_output(0));
  and_599_nl <= (fsm_output(6)) AND mux_1554_nl;
  nor_1168_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR (fsm_output(2)) OR (fsm_output(10)));
  nor_1170_nl <= NOT((fsm_output(7)) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR not_tmp_253);
  mux_1546_nl <= MUX_s_1_2_2(nor_1445_cse, nor_1170_nl, fsm_output(5));
  nor_1171_nl <= NOT((NOT (fsm_output(5))) OR (fsm_output(7)) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0110")) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR not_tmp_253);
  or_1323_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm);
  mux_1547_nl <= MUX_s_1_2_2(mux_1546_nl, nor_1171_nl, or_1323_nl);
  mux_1548_nl <= MUX_s_1_2_2(nor_1168_nl, mux_1547_nl, fsm_output(1));
  nor_1172_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR
      (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_253);
  nor_1173_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (NOT
      (fsm_output(2))) OR (fsm_output(10)));
  nor_1174_nl <= NOT((fsm_output(7)) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9))) OR (fsm_output(2)) OR (fsm_output(10)));
  mux_1544_nl <= MUX_s_1_2_2(nor_1173_nl, nor_1174_nl, fsm_output(5));
  mux_1545_nl <= MUX_s_1_2_2(nor_1172_nl, mux_1544_nl, fsm_output(1));
  mux_1549_nl <= MUX_s_1_2_2(mux_1548_nl, mux_1545_nl, fsm_output(0));
  nor_1175_nl <= NOT((NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (NOT (fsm_output(5)))
      OR (fsm_output(7)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR not_tmp_253);
  nor_1176_nl <= NOT((NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (NOT (fsm_output(5)))
      OR (fsm_output(7)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(3)) OR (fsm_output(9)) OR (NOT (fsm_output(2))) OR (fsm_output(10)));
  mux_1542_nl <= MUX_s_1_2_2(nor_1175_nl, nor_1176_nl, fsm_output(1));
  nor_1177_nl <= NOT((fsm_output(1)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO
      0)/=STD_LOGIC_VECTOR'("10")) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR mux_1413_cse);
  mux_1543_nl <= MUX_s_1_2_2(mux_1542_nl, nor_1177_nl, fsm_output(0));
  mux_1550_nl <= MUX_s_1_2_2(mux_1549_nl, mux_1543_nl, fsm_output(6));
  mux_1555_nl <= MUX_s_1_2_2(and_599_nl, mux_1550_nl, fsm_output(8));
  nor_1178_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (fsm_output(2))
      OR (fsm_output(10)));
  nor_1179_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(7)) OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(2)))
      OR (fsm_output(10)));
  mux_1536_nl <= MUX_s_1_2_2(nor_1178_nl, nor_1179_nl, fsm_output(5));
  and_600_nl <= COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm AND mux_1536_nl;
  nor_1180_nl <= NOT((NOT (fsm_output(7))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0110")) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR not_tmp_253);
  nor_1181_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(7)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9))) OR (fsm_output(2))
      OR (NOT (fsm_output(10))));
  mux_1535_nl <= MUX_s_1_2_2(nor_1180_nl, nor_1181_nl, fsm_output(5));
  and_601_nl <= COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm AND mux_1535_nl;
  mux_1537_nl <= MUX_s_1_2_2(and_600_nl, and_601_nl, fsm_output(1));
  nor_1182_nl <= NOT((VEC_LOOP_j_sva_11_0(3)) OR (NOT (VEC_LOOP_j_sva_11_0(1))) OR
      (VEC_LOOP_j_sva_11_0(0)) OR (NOT (fsm_output(5))) OR (NOT (VEC_LOOP_j_sva_11_0(2)))
      OR (fsm_output(7)) OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(2))
      OR (fsm_output(10)));
  nor_1183_nl <= NOT((VEC_LOOP_j_sva_11_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR mux_1533_cse);
  mux_1534_nl <= MUX_s_1_2_2(nor_1182_nl, nor_1183_nl, fsm_output(1));
  mux_1538_nl <= MUX_s_1_2_2(mux_1537_nl, mux_1534_nl, fsm_output(0));
  nor_1184_nl <= NOT((NOT (fsm_output(1))) OR (fsm_output(5)) OR (fsm_output(7))
      OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110")) OR (NOT
      (fsm_output(3))) OR (fsm_output(9)) OR (fsm_output(2)) OR (fsm_output(10)));
  nor_1185_nl <= NOT((fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(3)))
      OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110")) OR (NOT
      (fsm_output(9))) OR (NOT (fsm_output(2))) OR (fsm_output(10)));
  nor_1186_nl <= NOT((VEC_LOOP_j_sva_11_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (NOT
      (fsm_output(2))) OR (fsm_output(10)));
  mux_1531_nl <= MUX_s_1_2_2(nor_1185_nl, nor_1186_nl, fsm_output(1));
  mux_1532_nl <= MUX_s_1_2_2(nor_1184_nl, mux_1531_nl, fsm_output(0));
  mux_1539_nl <= MUX_s_1_2_2(mux_1538_nl, mux_1532_nl, fsm_output(6));
  nor_1187_nl <= NOT((NOT (fsm_output(1))) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(3)) OR (NOT (fsm_output(9)))
      OR (fsm_output(2)) OR (fsm_output(10)));
  nor_1188_nl <= NOT((fsm_output(1)) OR (fsm_output(5)) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0110")) OR (NOT (fsm_output(7))) OR (fsm_output(3))
      OR (fsm_output(9)) OR not_tmp_253);
  mux_1529_nl <= MUX_s_1_2_2(nor_1187_nl, nor_1188_nl, fsm_output(0));
  nor_1189_nl <= NOT((NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0110")) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR not_tmp_253);
  nor_1190_nl <= NOT((NOT (fsm_output(7))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0110")) OR (fsm_output(3)) OR (NOT (fsm_output(9)))
      OR (fsm_output(2)) OR (fsm_output(10)));
  nor_1191_nl <= NOT((NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR not_tmp_253);
  mux_1525_nl <= MUX_s_1_2_2(nor_1190_nl, nor_1191_nl, fsm_output(5));
  mux_1526_nl <= MUX_s_1_2_2(nor_1189_nl, mux_1525_nl, COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm);
  nor_1192_nl <= NOT((NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0110")) OR (fsm_output(3)) OR (fsm_output(9))
      OR (NOT (fsm_output(2))) OR (fsm_output(10)));
  mux_1527_nl <= MUX_s_1_2_2(mux_1526_nl, nor_1192_nl, fsm_output(1));
  nor_1193_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3)))
      OR (NOT (fsm_output(9))) OR (fsm_output(2)) OR (fsm_output(10)));
  nor_1194_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (VEC_LOOP_j_sva_11_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR
      (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(3)) OR (fsm_output(9))
      OR (fsm_output(2)) OR (NOT (fsm_output(10))));
  mux_1524_nl <= MUX_s_1_2_2(nor_1193_nl, nor_1194_nl, fsm_output(1));
  mux_1528_nl <= MUX_s_1_2_2(mux_1527_nl, mux_1524_nl, fsm_output(0));
  mux_1530_nl <= MUX_s_1_2_2(mux_1529_nl, mux_1528_nl, fsm_output(6));
  mux_1540_nl <= MUX_s_1_2_2(mux_1539_nl, mux_1530_nl, fsm_output(8));
  vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_1555_nl, mux_1540_nl,
      fsm_output(4));
  nand_302_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("01"))
      AND (VEC_LOOP_j_sva_11_0(1)) AND (fsm_output(5)) AND (VEC_LOOP_j_sva_11_0(0))
      AND CONV_SL_1_1(fsm_output(10 DOWNTO 9)=STD_LOGIC_VECTOR'("01")));
  nand_401_nl <= NOT((fsm_output(5)) AND (fsm_output(9)) AND CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)=STD_LOGIC_VECTOR'("0111")) AND (fsm_output(10)));
  mux_1582_nl <= MUX_s_1_2_2(nand_302_nl, nand_401_nl, fsm_output(7));
  or_1388_nl <= CONV_SL_1_1(VEC_LOOP_j_sva_11_0(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01"))
      OR (NOT (fsm_output(7))) OR (NOT (VEC_LOOP_j_sva_11_0(1))) OR (fsm_output(5))
      OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR CONV_SL_1_1(fsm_output(10 DOWNTO 9)/=STD_LOGIC_VECTOR'("00"));
  mux_1583_nl <= MUX_s_1_2_2(mux_1582_nl, or_1388_nl, fsm_output(2));
  nor_1149_nl <= NOT((fsm_output(6)) OR (fsm_output(4)) OR mux_1583_nl);
  nor_1150_nl <= NOT((fsm_output(6)) OR (fsm_output(4)) OR (NOT (fsm_output(2)))
      OR (fsm_output(7)) OR (fsm_output(5)) OR (fsm_output(9)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0111")) OR (NOT (fsm_output(10))));
  mux_1584_nl <= MUX_s_1_2_2(nor_1149_nl, nor_1150_nl, fsm_output(8));
  and_762_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0111"))
      AND (fsm_output(6)) AND (fsm_output(4)) AND (NOT (fsm_output(2))) AND (fsm_output(7))
      AND (fsm_output(5)) AND (NOT (fsm_output(9))) AND (fsm_output(10));
  nor_1152_nl <= NOT((fsm_output(4)) OR (fsm_output(2)) OR (fsm_output(7)) OR (fsm_output(5))
      OR (NOT (fsm_output(9))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("0111")) OR (fsm_output(10)));
  nor_1153_nl <= NOT((NOT (fsm_output(2))) OR (fsm_output(7)) OR (NOT (fsm_output(5)))
      OR (fsm_output(9)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("0111")) OR (fsm_output(10)));
  nor_1154_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (NOT (fsm_output(2))) OR (fsm_output(7)) OR (fsm_output(5)) OR (NOT (fsm_output(9)))
      OR (fsm_output(10)));
  mux_1579_nl <= MUX_s_1_2_2(nor_1153_nl, nor_1154_nl, fsm_output(4));
  mux_1580_nl <= MUX_s_1_2_2(nor_1152_nl, mux_1579_nl, fsm_output(6));
  mux_1581_nl <= MUX_s_1_2_2(and_762_nl, mux_1580_nl, fsm_output(8));
  mux_1585_nl <= MUX_s_1_2_2(mux_1584_nl, mux_1581_nl, fsm_output(0));
  nand_305_nl <= NOT((NOT (COMP_LOOP_acc_16_psp_sva(0))) AND (fsm_output(4)) AND
      (fsm_output(2)) AND (VEC_LOOP_j_sva_11_0(2)) AND (fsm_output(7)) AND (VEC_LOOP_j_sva_11_0(1))
      AND (fsm_output(5)) AND (VEC_LOOP_j_sva_11_0(0)) AND CONV_SL_1_1(fsm_output(10
      DOWNTO 9)=STD_LOGIC_VECTOR'("01")));
  or_1378_nl <= CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR (fsm_output(2)) OR (fsm_output(7)) OR (NOT (VEC_LOOP_j_sva_11_0(1))) OR
      (fsm_output(5)) OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR CONV_SL_1_1(fsm_output(10
      DOWNTO 9)/=STD_LOGIC_VECTOR'("10"));
  mux_1576_nl <= MUX_s_1_2_2(mux_tmp_1564, or_1378_nl, fsm_output(4));
  mux_1577_nl <= MUX_s_1_2_2(nand_305_nl, mux_1576_nl, fsm_output(6));
  and_598_nl <= (fsm_output(8)) AND (NOT mux_1577_nl);
  or_1375_nl <= (NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0111"))
      AND (fsm_output(2)) AND (fsm_output(7)) AND (NOT (fsm_output(5))))) OR nand_358_cse;
  nand_400_nl <= NOT((NOT (fsm_output(7))) AND (fsm_output(5)) AND (fsm_output(9))
      AND CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0111"))
      AND (fsm_output(10)));
  mux_1573_nl <= MUX_s_1_2_2(nand_400_nl, or_tmp_1308, fsm_output(2));
  mux_1574_nl <= MUX_s_1_2_2(or_1375_nl, mux_1573_nl, fsm_output(4));
  nor_1155_nl <= NOT((fsm_output(6)) OR mux_1574_nl);
  nor_1156_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(6)) OR (NOT (fsm_output(4))) OR (fsm_output(2)) OR (NOT (fsm_output(7)))
      OR (NOT (fsm_output(5))) OR (fsm_output(9)) OR (fsm_output(10)));
  mux_1575_nl <= MUX_s_1_2_2(nor_1155_nl, nor_1156_nl, fsm_output(8));
  mux_1578_nl <= MUX_s_1_2_2(and_598_nl, mux_1575_nl, fsm_output(0));
  mux_1586_nl <= MUX_s_1_2_2(mux_1585_nl, mux_1578_nl, fsm_output(3));
  or_1369_nl <= CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (NOT (fsm_output(2))) OR (fsm_output(7)) OR nand_334_cse;
  or_1367_nl <= (NOT (fsm_output(2))) OR (fsm_output(7)) OR (NOT (fsm_output(5)))
      OR (fsm_output(9)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("0111")) OR (NOT (fsm_output(10)));
  mux_1569_nl <= MUX_s_1_2_2(or_1369_nl, or_1367_nl, fsm_output(4));
  nor_1157_nl <= NOT((fsm_output(6)) OR mux_1569_nl);
  or_1361_nl <= (fsm_output(5)) OR (fsm_output(9)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0111")) OR (NOT (fsm_output(10)));
  mux_1567_nl <= MUX_s_1_2_2(or_702_cse, or_1361_nl, fsm_output(7));
  mux_1568_nl <= MUX_s_1_2_2(or_tmp_1308, mux_1567_nl, nor_223_cse);
  nor_1158_nl <= NOT((NOT (fsm_output(6))) OR (NOT (fsm_output(4))) OR (fsm_output(2))
      OR mux_1568_nl);
  mux_1570_nl <= MUX_s_1_2_2(nor_1157_nl, nor_1158_nl, fsm_output(8));
  or_1357_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(7)) OR (NOT (fsm_output(5))) OR (fsm_output(9)) OR (NOT (fsm_output(10)));
  or_1355_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (NOT (fsm_output(7))) OR (fsm_output(5)) OR (NOT (fsm_output(9))) OR (fsm_output(10));
  mux_1565_nl <= MUX_s_1_2_2(or_1357_nl, or_1355_nl, fsm_output(2));
  mux_1566_nl <= MUX_s_1_2_2(mux_1565_nl, mux_tmp_1564, fsm_output(4));
  nor_1159_nl <= NOT((fsm_output(8)) OR (fsm_output(6)) OR mux_1566_nl);
  mux_1571_nl <= MUX_s_1_2_2(mux_1570_nl, nor_1159_nl, fsm_output(0));
  or_1350_nl <= CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (fsm_output(2)) OR (NOT (fsm_output(7))) OR (fsm_output(5)) OR (NOT (VEC_LOOP_j_sva_11_0(0)))
      OR CONV_SL_1_1(fsm_output(10 DOWNTO 9)/=STD_LOGIC_VECTOR'("10"));
  or_1348_nl <= (fsm_output(2)) OR (NOT (fsm_output(7))) OR (fsm_output(5)) OR (NOT
      (fsm_output(9))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(10));
  mux_1561_nl <= MUX_s_1_2_2(or_1350_nl, or_1348_nl, fsm_output(4));
  nand_310_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("011"))
      AND (fsm_output(2)) AND (fsm_output(7)) AND (fsm_output(5)) AND (VEC_LOOP_j_sva_11_0(0))
      AND CONV_SL_1_1(fsm_output(10 DOWNTO 9)=STD_LOGIC_VECTOR'("01")));
  or_1346_nl <= (NOT (fsm_output(2))) OR (NOT (fsm_output(7))) OR (NOT (fsm_output(5)))
      OR (fsm_output(9)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("0111")) OR (fsm_output(10));
  mux_1560_nl <= MUX_s_1_2_2(nand_310_nl, or_1346_nl, fsm_output(4));
  mux_1562_nl <= MUX_s_1_2_2(mux_1561_nl, mux_1560_nl, fsm_output(6));
  nor_1160_nl <= NOT((fsm_output(8)) OR mux_1562_nl);
  nor_1161_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (NOT (fsm_output(6))) OR (fsm_output(4)) OR (fsm_output(2)) OR (NOT (fsm_output(7)))
      OR (NOT (fsm_output(5))) OR (fsm_output(9)) OR (fsm_output(10)));
  and_763_nl <= (fsm_output(4)) AND (fsm_output(2)) AND (fsm_output(7)) AND CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3
      DOWNTO 0)=STD_LOGIC_VECTOR'("0111")) AND (fsm_output(5)) AND (NOT (fsm_output(9)))
      AND (fsm_output(10));
  or_1341_nl <= (fsm_output(7)) OR (NOT (fsm_output(5))) OR (fsm_output(9)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0111")) OR (NOT (fsm_output(10)));
  or_1339_nl <= (NOT (fsm_output(7))) OR (fsm_output(5)) OR (NOT (fsm_output(9)))
      OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(10));
  mux_1557_nl <= MUX_s_1_2_2(or_1341_nl, or_1339_nl, fsm_output(2));
  nor_1163_nl <= NOT((fsm_output(4)) OR mux_1557_nl);
  mux_1558_nl <= MUX_s_1_2_2(and_763_nl, nor_1163_nl, fsm_output(6));
  mux_1559_nl <= MUX_s_1_2_2(nor_1161_nl, mux_1558_nl, fsm_output(8));
  mux_1563_nl <= MUX_s_1_2_2(nor_1160_nl, mux_1559_nl, fsm_output(0));
  mux_1572_nl <= MUX_s_1_2_2(mux_1571_nl, mux_1563_nl, fsm_output(3));
  vec_rsc_0_7_i_wea_d_pff <= MUX_s_1_2_2(mux_1586_nl, mux_1572_nl, fsm_output(1));
  or_1447_nl <= (NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(2))) OR (fsm_output(10));
  or_1446_nl <= (fsm_output(7)) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(2)) OR (NOT (fsm_output(10)));
  mux_1617_nl <= MUX_s_1_2_2(or_1447_nl, or_1446_nl, fsm_output(5));
  nor_1120_nl <= NOT((fsm_output(1)) OR mux_1617_nl);
  nor_1121_nl <= NOT((fsm_output(5)) OR (NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0111")) OR (fsm_output(3)) OR (fsm_output(9))
      OR (fsm_output(2)) OR (fsm_output(10)));
  nor_1122_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (NOT (fsm_output(7))) OR (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_253);
  nor_1123_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(7)) OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (fsm_output(2))
      OR (NOT (fsm_output(10))));
  mux_1615_nl <= MUX_s_1_2_2(nor_1122_nl, nor_1123_nl, fsm_output(5));
  mux_1616_nl <= MUX_s_1_2_2(nor_1121_nl, mux_1615_nl, fsm_output(1));
  mux_1618_nl <= MUX_s_1_2_2(nor_1120_nl, mux_1616_nl, fsm_output(0));
  and_593_nl <= (fsm_output(6)) AND mux_1618_nl;
  nor_1124_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR (fsm_output(2)) OR (fsm_output(10)));
  nor_1126_nl <= NOT((fsm_output(7)) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR not_tmp_253);
  mux_1610_nl <= MUX_s_1_2_2(nor_1445_cse, nor_1126_nl, fsm_output(5));
  nor_1127_nl <= NOT((NOT (fsm_output(5))) OR (fsm_output(7)) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0111")) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR not_tmp_253);
  nand_295_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0111"))
      AND COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm);
  mux_1611_nl <= MUX_s_1_2_2(mux_1610_nl, nor_1127_nl, nand_295_nl);
  mux_1612_nl <= MUX_s_1_2_2(nor_1124_nl, mux_1611_nl, fsm_output(1));
  nor_1128_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11")) OR
      (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_253);
  nor_1129_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (NOT
      (fsm_output(2))) OR (fsm_output(10)));
  nor_1130_nl <= NOT((fsm_output(7)) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9))) OR (fsm_output(2)) OR (fsm_output(10)));
  mux_1608_nl <= MUX_s_1_2_2(nor_1129_nl, nor_1130_nl, fsm_output(5));
  mux_1609_nl <= MUX_s_1_2_2(nor_1128_nl, mux_1608_nl, fsm_output(1));
  mux_1613_nl <= MUX_s_1_2_2(mux_1612_nl, mux_1609_nl, fsm_output(0));
  nor_1131_nl <= NOT((NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (NOT (fsm_output(5)))
      OR (fsm_output(7)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR not_tmp_253);
  nor_1132_nl <= NOT((NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (NOT (fsm_output(5)))
      OR (fsm_output(7)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(3)) OR (fsm_output(9)) OR (NOT (fsm_output(2))) OR (fsm_output(10)));
  mux_1606_nl <= MUX_s_1_2_2(nor_1131_nl, nor_1132_nl, fsm_output(1));
  nor_1133_nl <= NOT(nand_324_cse OR mux_1413_cse);
  mux_1607_nl <= MUX_s_1_2_2(mux_1606_nl, nor_1133_nl, fsm_output(0));
  mux_1614_nl <= MUX_s_1_2_2(mux_1613_nl, mux_1607_nl, fsm_output(6));
  mux_1619_nl <= MUX_s_1_2_2(and_593_nl, mux_1614_nl, fsm_output(8));
  nor_1134_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (fsm_output(2))
      OR (fsm_output(10)));
  nor_1135_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(7)) OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(2)))
      OR (fsm_output(10)));
  mux_1600_nl <= MUX_s_1_2_2(nor_1134_nl, nor_1135_nl, fsm_output(5));
  and_594_nl <= COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm AND mux_1600_nl;
  nor_1136_nl <= NOT((NOT((fsm_output(7)) AND CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3
      DOWNTO 0)=STD_LOGIC_VECTOR'("0111")) AND (fsm_output(3)) AND (NOT (fsm_output(9)))))
      OR not_tmp_253);
  nor_1137_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(7)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9))) OR (fsm_output(2))
      OR (NOT (fsm_output(10))));
  mux_1599_nl <= MUX_s_1_2_2(nor_1136_nl, nor_1137_nl, fsm_output(5));
  and_595_nl <= COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm AND mux_1599_nl;
  mux_1601_nl <= MUX_s_1_2_2(and_594_nl, and_595_nl, fsm_output(1));
  nor_1138_nl <= NOT((VEC_LOOP_j_sva_11_0(3)) OR (NOT (VEC_LOOP_j_sva_11_0(1))) OR
      (NOT (VEC_LOOP_j_sva_11_0(0))) OR (NOT (fsm_output(5))) OR (NOT (VEC_LOOP_j_sva_11_0(2)))
      OR (fsm_output(7)) OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(2))
      OR (fsm_output(10)));
  nor_1139_nl <= NOT(nand_332_cse OR mux_1533_cse);
  mux_1598_nl <= MUX_s_1_2_2(nor_1138_nl, nor_1139_nl, fsm_output(1));
  mux_1602_nl <= MUX_s_1_2_2(mux_1601_nl, mux_1598_nl, fsm_output(0));
  nor_1140_nl <= NOT((NOT (fsm_output(1))) OR (fsm_output(5)) OR (fsm_output(7))
      OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111")) OR (NOT
      (fsm_output(3))) OR (fsm_output(9)) OR (fsm_output(2)) OR (fsm_output(10)));
  nor_1141_nl <= NOT((fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(3)))
      OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111")) OR (NOT
      (fsm_output(9))) OR (NOT (fsm_output(2))) OR (fsm_output(10)));
  and_596_nl <= (VEC_LOOP_j_sva_11_0(0)) AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm
      AND (fsm_output(5)) AND CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("011"))
      AND (fsm_output(7)) AND (fsm_output(3)) AND (NOT (fsm_output(9))) AND (fsm_output(2))
      AND (NOT (fsm_output(10)));
  mux_1595_nl <= MUX_s_1_2_2(nor_1141_nl, and_596_nl, fsm_output(1));
  mux_1596_nl <= MUX_s_1_2_2(nor_1140_nl, mux_1595_nl, fsm_output(0));
  mux_1603_nl <= MUX_s_1_2_2(mux_1602_nl, mux_1596_nl, fsm_output(6));
  nor_1142_nl <= NOT((NOT (fsm_output(1))) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(3)) OR (NOT (fsm_output(9)))
      OR (fsm_output(2)) OR (fsm_output(10)));
  nor_1143_nl <= NOT((fsm_output(1)) OR (fsm_output(5)) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0111")) OR (NOT (fsm_output(7))) OR (fsm_output(3))
      OR (fsm_output(9)) OR not_tmp_253);
  mux_1593_nl <= MUX_s_1_2_2(nor_1142_nl, nor_1143_nl, fsm_output(0));
  nor_1144_nl <= NOT((NOT((fsm_output(5)) AND (fsm_output(7)) AND CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)=STD_LOGIC_VECTOR'("0111")) AND (fsm_output(3)) AND (NOT (fsm_output(9)))))
      OR not_tmp_253);
  nor_1145_nl <= NOT((NOT (fsm_output(7))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0111")) OR (fsm_output(3)) OR (NOT (fsm_output(9)))
      OR (fsm_output(2)) OR (fsm_output(10)));
  nor_1146_nl <= NOT((NOT((fsm_output(7)) AND CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0111"))
      AND (fsm_output(3)) AND (NOT (fsm_output(9))))) OR not_tmp_253);
  mux_1589_nl <= MUX_s_1_2_2(nor_1145_nl, nor_1146_nl, fsm_output(5));
  mux_1590_nl <= MUX_s_1_2_2(nor_1144_nl, mux_1589_nl, COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm);
  nor_1147_nl <= NOT((NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0111")) OR (fsm_output(3)) OR (fsm_output(9))
      OR (NOT (fsm_output(2))) OR (fsm_output(10)));
  mux_1591_nl <= MUX_s_1_2_2(mux_1590_nl, nor_1147_nl, fsm_output(1));
  and_597_nl <= CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0111")) AND
      (fsm_output(5)) AND (fsm_output(7)) AND (fsm_output(3)) AND (fsm_output(9))
      AND (NOT (fsm_output(2))) AND (NOT (fsm_output(10)));
  nor_1148_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(3)) OR (fsm_output(9))
      OR (fsm_output(2)) OR (NOT (fsm_output(10))));
  mux_1588_nl <= MUX_s_1_2_2(and_597_nl, nor_1148_nl, fsm_output(1));
  mux_1592_nl <= MUX_s_1_2_2(mux_1591_nl, mux_1588_nl, fsm_output(0));
  mux_1594_nl <= MUX_s_1_2_2(mux_1593_nl, mux_1592_nl, fsm_output(6));
  mux_1604_nl <= MUX_s_1_2_2(mux_1603_nl, mux_1594_nl, fsm_output(8));
  vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_1619_nl, mux_1604_nl,
      fsm_output(4));
  or_1502_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR
      (NOT (fsm_output(9))) OR (NOT (fsm_output(5))) OR (fsm_output(10));
  or_1501_nl <= (NOT (fsm_output(9))) OR (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000")) OR not_tmp_318;
  mux_1646_nl <= MUX_s_1_2_2(or_1502_nl, or_1501_nl, fsm_output(7));
  or_1499_nl <= CONV_SL_1_1(VEC_LOOP_j_sva_11_0(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("10"))
      OR (NOT (fsm_output(7))) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (fsm_output(9)) OR (fsm_output(5)) OR (fsm_output(10));
  mux_1647_nl <= MUX_s_1_2_2(mux_1646_nl, or_1499_nl, fsm_output(2));
  nor_1105_nl <= NOT((fsm_output(6)) OR (fsm_output(4)) OR mux_1647_nl);
  nor_1106_nl <= NOT((fsm_output(6)) OR (fsm_output(4)) OR (NOT (fsm_output(2)))
      OR (fsm_output(7)) OR (fsm_output(9)) OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000")) OR not_tmp_318);
  mux_1648_nl <= MUX_s_1_2_2(nor_1105_nl, nor_1106_nl, fsm_output(8));
  nor_1107_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT (fsm_output(6))) OR (NOT (fsm_output(4))) OR (fsm_output(2)) OR (NOT
      (fsm_output(7))) OR (fsm_output(9)) OR not_tmp_248);
  nor_1108_nl <= NOT((fsm_output(4)) OR (fsm_output(2)) OR (fsm_output(7)) OR (NOT
      (fsm_output(9))) OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1000")) OR (fsm_output(10)));
  nor_1109_nl <= NOT((NOT (fsm_output(2))) OR (fsm_output(7)) OR (fsm_output(9))
      OR (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("1000")) OR (fsm_output(10)));
  nor_1110_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT (fsm_output(2))) OR (fsm_output(7)) OR (NOT (fsm_output(9))) OR (fsm_output(5))
      OR (fsm_output(10)));
  mux_1643_nl <= MUX_s_1_2_2(nor_1109_nl, nor_1110_nl, fsm_output(4));
  mux_1644_nl <= MUX_s_1_2_2(nor_1108_nl, mux_1643_nl, fsm_output(6));
  mux_1645_nl <= MUX_s_1_2_2(nor_1107_nl, mux_1644_nl, fsm_output(8));
  mux_1649_nl <= MUX_s_1_2_2(mux_1648_nl, mux_1645_nl, fsm_output(0));
  or_1490_nl <= (NOT (COMP_LOOP_acc_16_psp_sva(0))) OR (NOT (fsm_output(4))) OR (NOT
      (fsm_output(2))) OR (VEC_LOOP_j_sva_11_0(2)) OR (NOT (fsm_output(7))) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(5)))
      OR (fsm_output(10));
  or_1489_nl <= CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (fsm_output(2)) OR (fsm_output(7)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR (fsm_output(9)) OR (fsm_output(5)) OR
      (NOT (fsm_output(10)));
  mux_1640_nl <= MUX_s_1_2_2(mux_tmp_1628, or_1489_nl, fsm_output(4));
  mux_1641_nl <= MUX_s_1_2_2(or_1490_nl, mux_1640_nl, fsm_output(6));
  and_592_nl <= (fsm_output(8)) AND (NOT mux_1641_nl);
  or_1486_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(7))) OR (NOT (fsm_output(9)))
      OR (fsm_output(5)) OR (NOT (fsm_output(10)));
  or_1484_nl <= (fsm_output(7)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(5)))
      OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR not_tmp_318;
  mux_1637_nl <= MUX_s_1_2_2(or_1484_nl, or_tmp_1416, fsm_output(2));
  mux_1638_nl <= MUX_s_1_2_2(or_1486_nl, mux_1637_nl, fsm_output(4));
  nor_1111_nl <= NOT((fsm_output(6)) OR mux_1638_nl);
  nor_1112_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(6)) OR (NOT (fsm_output(4))) OR (fsm_output(2)) OR (NOT (fsm_output(7)))
      OR (fsm_output(9)) OR (NOT (fsm_output(5))) OR (fsm_output(10)));
  mux_1639_nl <= MUX_s_1_2_2(nor_1111_nl, nor_1112_nl, fsm_output(8));
  mux_1642_nl <= MUX_s_1_2_2(and_592_nl, mux_1639_nl, fsm_output(0));
  mux_1650_nl <= MUX_s_1_2_2(mux_1649_nl, mux_1642_nl, fsm_output(3));
  or_1480_nl <= CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (NOT (fsm_output(2))) OR (fsm_output(7)) OR (VEC_LOOP_j_sva_11_0(0)) OR
      nand_337_cse;
  or_1478_nl <= (NOT (fsm_output(2))) OR (fsm_output(7)) OR (fsm_output(9)) OR (NOT
      (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR not_tmp_318;
  mux_1633_nl <= MUX_s_1_2_2(or_1480_nl, or_1478_nl, fsm_output(4));
  nor_1113_nl <= NOT((fsm_output(6)) OR mux_1633_nl);
  or_1474_nl <= (fsm_output(9)) OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000")) OR not_tmp_318;
  mux_1631_nl <= MUX_s_1_2_2(or_591_cse, or_1474_nl, fsm_output(7));
  mux_1632_nl <= MUX_s_1_2_2(mux_1631_nl, or_tmp_1416, or_1470_cse);
  nor_1114_nl <= NOT((NOT (fsm_output(6))) OR (NOT (fsm_output(4))) OR (fsm_output(2))
      OR mux_1632_nl);
  mux_1634_nl <= MUX_s_1_2_2(nor_1113_nl, nor_1114_nl, fsm_output(8));
  or_1467_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(7)) OR (fsm_output(9)) OR not_tmp_248;
  or_1465_nl <= (NOT (fsm_output(7))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1000")) OR (NOT (fsm_output(9))) OR (fsm_output(5))
      OR (fsm_output(10));
  mux_1629_nl <= MUX_s_1_2_2(or_1467_nl, or_1465_nl, fsm_output(2));
  mux_1630_nl <= MUX_s_1_2_2(mux_1629_nl, mux_tmp_1628, fsm_output(4));
  nor_1115_nl <= NOT((fsm_output(8)) OR (fsm_output(6)) OR mux_1630_nl);
  mux_1635_nl <= MUX_s_1_2_2(mux_1634_nl, nor_1115_nl, fsm_output(0));
  or_1460_nl <= CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (fsm_output(2)) OR (NOT (fsm_output(7))) OR (VEC_LOOP_j_sva_11_0(0)) OR
      (fsm_output(9)) OR (fsm_output(5)) OR (NOT (fsm_output(10)));
  or_1458_nl <= (fsm_output(2)) OR (NOT (fsm_output(7))) OR (NOT (fsm_output(9)))
      OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("1000")) OR (fsm_output(10));
  mux_1625_nl <= MUX_s_1_2_2(or_1460_nl, or_1458_nl, fsm_output(4));
  or_1457_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(7))) OR (VEC_LOOP_j_sva_11_0(0))
      OR (NOT (fsm_output(9))) OR (NOT (fsm_output(5))) OR (fsm_output(10));
  or_1456_nl <= (NOT (fsm_output(2))) OR (NOT (fsm_output(7))) OR (fsm_output(9))
      OR (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("1000")) OR (fsm_output(10));
  mux_1624_nl <= MUX_s_1_2_2(or_1457_nl, or_1456_nl, fsm_output(4));
  mux_1626_nl <= MUX_s_1_2_2(mux_1625_nl, mux_1624_nl, fsm_output(6));
  nor_1116_nl <= NOT((fsm_output(8)) OR mux_1626_nl);
  nor_1117_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT (fsm_output(6))) OR (fsm_output(4)) OR (fsm_output(2)) OR (NOT (fsm_output(7)))
      OR (fsm_output(9)) OR (NOT (fsm_output(5))) OR (fsm_output(10)));
  nor_1118_nl <= NOT((NOT (fsm_output(4))) OR (NOT (fsm_output(2))) OR (NOT (fsm_output(7)))
      OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(9)) OR not_tmp_248);
  or_1451_nl <= (fsm_output(7)) OR (fsm_output(9)) OR (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000")) OR not_tmp_318;
  or_1449_nl <= (NOT (fsm_output(7))) OR (NOT (fsm_output(9))) OR (fsm_output(5))
      OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(10));
  mux_1621_nl <= MUX_s_1_2_2(or_1451_nl, or_1449_nl, fsm_output(2));
  nor_1119_nl <= NOT((fsm_output(4)) OR mux_1621_nl);
  mux_1622_nl <= MUX_s_1_2_2(nor_1118_nl, nor_1119_nl, fsm_output(6));
  mux_1623_nl <= MUX_s_1_2_2(nor_1117_nl, mux_1622_nl, fsm_output(8));
  mux_1627_nl <= MUX_s_1_2_2(nor_1116_nl, mux_1623_nl, fsm_output(0));
  mux_1636_nl <= MUX_s_1_2_2(mux_1635_nl, mux_1627_nl, fsm_output(3));
  vec_rsc_0_8_i_wea_d_pff <= MUX_s_1_2_2(mux_1650_nl, mux_1636_nl, fsm_output(1));
  or_1558_nl <= (NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(2))) OR (fsm_output(10));
  or_1557_nl <= (fsm_output(7)) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(2)) OR (NOT (fsm_output(10)));
  mux_1681_nl <= MUX_s_1_2_2(or_1558_nl, or_1557_nl, fsm_output(5));
  nor_1074_nl <= NOT((fsm_output(1)) OR mux_1681_nl);
  nor_1075_nl <= NOT((fsm_output(5)) OR (NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1000")) OR (fsm_output(3)) OR (fsm_output(9))
      OR (fsm_output(2)) OR (fsm_output(10)));
  nor_1076_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT (fsm_output(7))) OR (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_253);
  nor_1077_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(7)) OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (fsm_output(2))
      OR (NOT (fsm_output(10))));
  mux_1679_nl <= MUX_s_1_2_2(nor_1076_nl, nor_1077_nl, fsm_output(5));
  mux_1680_nl <= MUX_s_1_2_2(nor_1075_nl, mux_1679_nl, fsm_output(1));
  mux_1682_nl <= MUX_s_1_2_2(nor_1074_nl, mux_1680_nl, fsm_output(0));
  and_589_nl <= (fsm_output(6)) AND mux_1682_nl;
  nor_1078_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR (fsm_output(2)) OR (fsm_output(10)));
  nor_1080_nl <= NOT((fsm_output(7)) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR not_tmp_253);
  mux_1674_nl <= MUX_s_1_2_2(nor_1445_cse, nor_1080_nl, fsm_output(5));
  nor_1081_nl <= NOT((NOT (fsm_output(5))) OR (fsm_output(7)) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1000")) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR not_tmp_253);
  or_1544_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm);
  mux_1675_nl <= MUX_s_1_2_2(mux_1674_nl, nor_1081_nl, or_1544_nl);
  mux_1676_nl <= MUX_s_1_2_2(nor_1078_nl, mux_1675_nl, fsm_output(1));
  nor_1082_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR
      (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_253);
  nor_1083_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (NOT
      (fsm_output(2))) OR (fsm_output(10)));
  nor_1084_nl <= NOT((fsm_output(7)) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9))) OR (fsm_output(2)) OR (fsm_output(10)));
  mux_1672_nl <= MUX_s_1_2_2(nor_1083_nl, nor_1084_nl, fsm_output(5));
  mux_1673_nl <= MUX_s_1_2_2(nor_1082_nl, mux_1672_nl, fsm_output(1));
  mux_1677_nl <= MUX_s_1_2_2(mux_1676_nl, mux_1673_nl, fsm_output(0));
  nor_1085_nl <= NOT((NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (NOT (fsm_output(5)))
      OR (fsm_output(7)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR not_tmp_253);
  nor_1086_nl <= NOT((NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (NOT (fsm_output(5)))
      OR (fsm_output(7)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(3)) OR (fsm_output(9)) OR (NOT (fsm_output(2))) OR (fsm_output(10)));
  mux_1670_nl <= MUX_s_1_2_2(nor_1085_nl, nor_1086_nl, fsm_output(1));
  nor_1087_nl <= NOT((fsm_output(1)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO
      0)/=STD_LOGIC_VECTOR'("00")) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR mux_1669_cse);
  mux_1671_nl <= MUX_s_1_2_2(mux_1670_nl, nor_1087_nl, fsm_output(0));
  mux_1678_nl <= MUX_s_1_2_2(mux_1677_nl, mux_1671_nl, fsm_output(6));
  mux_1683_nl <= MUX_s_1_2_2(and_589_nl, mux_1678_nl, fsm_output(8));
  nor_1088_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (fsm_output(2))
      OR (fsm_output(10)));
  nor_1089_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(7)) OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(2)))
      OR (fsm_output(10)));
  mux_1664_nl <= MUX_s_1_2_2(nor_1088_nl, nor_1089_nl, fsm_output(5));
  and_590_nl <= COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm AND mux_1664_nl;
  nor_1090_nl <= NOT((NOT (fsm_output(7))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1000")) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR not_tmp_253);
  nor_1091_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(7)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9))) OR (fsm_output(2))
      OR (NOT (fsm_output(10))));
  mux_1663_nl <= MUX_s_1_2_2(nor_1090_nl, nor_1091_nl, fsm_output(5));
  and_591_nl <= COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm AND mux_1663_nl;
  mux_1665_nl <= MUX_s_1_2_2(and_590_nl, and_591_nl, fsm_output(1));
  nor_1092_nl <= NOT((NOT (VEC_LOOP_j_sva_11_0(3))) OR (VEC_LOOP_j_sva_11_0(1)) OR
      (VEC_LOOP_j_sva_11_0(0)) OR (NOT (fsm_output(5))) OR (VEC_LOOP_j_sva_11_0(2))
      OR (fsm_output(7)) OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(2))
      OR (fsm_output(10)));
  nor_1093_nl <= NOT((VEC_LOOP_j_sva_11_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR mux_1661_cse);
  mux_1662_nl <= MUX_s_1_2_2(nor_1092_nl, nor_1093_nl, fsm_output(1));
  mux_1666_nl <= MUX_s_1_2_2(mux_1665_nl, mux_1662_nl, fsm_output(0));
  nor_1094_nl <= NOT((NOT (fsm_output(1))) OR (fsm_output(5)) OR (fsm_output(7))
      OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000")) OR (NOT
      (fsm_output(3))) OR (fsm_output(9)) OR (fsm_output(2)) OR (fsm_output(10)));
  nor_1095_nl <= NOT((fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(3)))
      OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000")) OR (NOT
      (fsm_output(9))) OR (NOT (fsm_output(2))) OR (fsm_output(10)));
  nor_1096_nl <= NOT((VEC_LOOP_j_sva_11_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (NOT
      (fsm_output(2))) OR (fsm_output(10)));
  mux_1659_nl <= MUX_s_1_2_2(nor_1095_nl, nor_1096_nl, fsm_output(1));
  mux_1660_nl <= MUX_s_1_2_2(nor_1094_nl, mux_1659_nl, fsm_output(0));
  mux_1667_nl <= MUX_s_1_2_2(mux_1666_nl, mux_1660_nl, fsm_output(6));
  nor_1097_nl <= NOT((NOT (fsm_output(1))) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(3)) OR (NOT (fsm_output(9)))
      OR (fsm_output(2)) OR (fsm_output(10)));
  nor_1098_nl <= NOT((fsm_output(1)) OR (fsm_output(5)) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1000")) OR (NOT (fsm_output(7))) OR (fsm_output(3))
      OR (fsm_output(9)) OR not_tmp_253);
  mux_1657_nl <= MUX_s_1_2_2(nor_1097_nl, nor_1098_nl, fsm_output(0));
  nor_1099_nl <= NOT((NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1000")) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR not_tmp_253);
  nor_1100_nl <= NOT((NOT (fsm_output(7))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1000")) OR (fsm_output(3)) OR (NOT (fsm_output(9)))
      OR (fsm_output(2)) OR (fsm_output(10)));
  nor_1101_nl <= NOT((NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR not_tmp_253);
  mux_1653_nl <= MUX_s_1_2_2(nor_1100_nl, nor_1101_nl, fsm_output(5));
  mux_1654_nl <= MUX_s_1_2_2(nor_1099_nl, mux_1653_nl, COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm);
  nor_1102_nl <= NOT((NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1000")) OR (fsm_output(3)) OR (fsm_output(9))
      OR (NOT (fsm_output(2))) OR (fsm_output(10)));
  mux_1655_nl <= MUX_s_1_2_2(mux_1654_nl, nor_1102_nl, fsm_output(1));
  nor_1103_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3)))
      OR (NOT (fsm_output(9))) OR (fsm_output(2)) OR (fsm_output(10)));
  nor_1104_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (VEC_LOOP_j_sva_11_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR
      (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(3)) OR (fsm_output(9))
      OR (fsm_output(2)) OR (NOT (fsm_output(10))));
  mux_1652_nl <= MUX_s_1_2_2(nor_1103_nl, nor_1104_nl, fsm_output(1));
  mux_1656_nl <= MUX_s_1_2_2(mux_1655_nl, mux_1652_nl, fsm_output(0));
  mux_1658_nl <= MUX_s_1_2_2(mux_1657_nl, mux_1656_nl, fsm_output(6));
  mux_1668_nl <= MUX_s_1_2_2(mux_1667_nl, mux_1658_nl, fsm_output(8));
  vec_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_1683_nl, mux_1668_nl,
      fsm_output(4));
  or_1613_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR
      (NOT (fsm_output(9))) OR (NOT (fsm_output(5))) OR (fsm_output(10));
  or_1612_nl <= (NOT (fsm_output(9))) OR (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001")) OR not_tmp_318;
  mux_1710_nl <= MUX_s_1_2_2(or_1613_nl, or_1612_nl, fsm_output(7));
  or_1610_nl <= CONV_SL_1_1(VEC_LOOP_j_sva_11_0(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("10"))
      OR (NOT (fsm_output(7))) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR (fsm_output(9)) OR (fsm_output(5)) OR (fsm_output(10));
  mux_1711_nl <= MUX_s_1_2_2(mux_1710_nl, or_1610_nl, fsm_output(2));
  nor_1059_nl <= NOT((fsm_output(6)) OR (fsm_output(4)) OR mux_1711_nl);
  nor_1060_nl <= NOT((fsm_output(6)) OR (fsm_output(4)) OR (NOT (fsm_output(2)))
      OR (fsm_output(7)) OR (fsm_output(9)) OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001")) OR not_tmp_318);
  mux_1712_nl <= MUX_s_1_2_2(nor_1059_nl, nor_1060_nl, fsm_output(8));
  nor_1061_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT (fsm_output(6))) OR (NOT (fsm_output(4))) OR (fsm_output(2)) OR (NOT
      (fsm_output(7))) OR (fsm_output(9)) OR not_tmp_248);
  nor_1062_nl <= NOT((fsm_output(4)) OR (fsm_output(2)) OR (fsm_output(7)) OR (NOT
      (fsm_output(9))) OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1001")) OR (fsm_output(10)));
  nor_1063_nl <= NOT((NOT (fsm_output(2))) OR (fsm_output(7)) OR (fsm_output(9))
      OR (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("1001")) OR (fsm_output(10)));
  nor_1064_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT (fsm_output(2))) OR (fsm_output(7)) OR (NOT (fsm_output(9))) OR (fsm_output(5))
      OR (fsm_output(10)));
  mux_1707_nl <= MUX_s_1_2_2(nor_1063_nl, nor_1064_nl, fsm_output(4));
  mux_1708_nl <= MUX_s_1_2_2(nor_1062_nl, mux_1707_nl, fsm_output(6));
  mux_1709_nl <= MUX_s_1_2_2(nor_1061_nl, mux_1708_nl, fsm_output(8));
  mux_1713_nl <= MUX_s_1_2_2(mux_1712_nl, mux_1709_nl, fsm_output(0));
  nand_287_nl <= NOT((COMP_LOOP_acc_16_psp_sva(0)) AND (fsm_output(4)) AND (fsm_output(2))
      AND (NOT (VEC_LOOP_j_sva_11_0(2))) AND (fsm_output(7)) AND CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1
      DOWNTO 0)=STD_LOGIC_VECTOR'("01")) AND (fsm_output(9)) AND (fsm_output(5))
      AND (NOT (fsm_output(10))));
  or_1600_nl <= CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (fsm_output(2)) OR (fsm_output(7)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR (fsm_output(9)) OR (fsm_output(5)) OR
      (NOT (fsm_output(10)));
  mux_1704_nl <= MUX_s_1_2_2(mux_tmp_1692, or_1600_nl, fsm_output(4));
  mux_1705_nl <= MUX_s_1_2_2(nand_287_nl, mux_1704_nl, fsm_output(6));
  and_588_nl <= (fsm_output(8)) AND (NOT mux_1705_nl);
  or_1597_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(7))) OR (NOT (fsm_output(9)))
      OR (fsm_output(5)) OR (NOT (fsm_output(10)));
  or_1595_nl <= (fsm_output(7)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(5)))
      OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR not_tmp_318;
  mux_1701_nl <= MUX_s_1_2_2(or_1595_nl, or_tmp_1527, fsm_output(2));
  mux_1702_nl <= MUX_s_1_2_2(or_1597_nl, mux_1701_nl, fsm_output(4));
  nor_1065_nl <= NOT((fsm_output(6)) OR mux_1702_nl);
  nor_1066_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(6)) OR (NOT (fsm_output(4))) OR (fsm_output(2)) OR (NOT (fsm_output(7)))
      OR (fsm_output(9)) OR (NOT (fsm_output(5))) OR (fsm_output(10)));
  mux_1703_nl <= MUX_s_1_2_2(nor_1065_nl, nor_1066_nl, fsm_output(8));
  mux_1706_nl <= MUX_s_1_2_2(and_588_nl, mux_1703_nl, fsm_output(0));
  mux_1714_nl <= MUX_s_1_2_2(mux_1713_nl, mux_1706_nl, fsm_output(3));
  or_1591_nl <= CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (NOT (fsm_output(2))) OR (fsm_output(7)) OR nand_334_cse;
  or_1589_nl <= (NOT (fsm_output(2))) OR (fsm_output(7)) OR (fsm_output(9)) OR (NOT
      (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR not_tmp_318;
  mux_1697_nl <= MUX_s_1_2_2(or_1591_nl, or_1589_nl, fsm_output(4));
  nor_1067_nl <= NOT((fsm_output(6)) OR mux_1697_nl);
  or_1585_nl <= (fsm_output(9)) OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001")) OR not_tmp_318;
  mux_1695_nl <= MUX_s_1_2_2(or_702_cse, or_1585_nl, fsm_output(7));
  mux_1696_nl <= MUX_s_1_2_2(mux_1695_nl, or_tmp_1527, or_1470_cse);
  nor_1068_nl <= NOT((NOT (fsm_output(6))) OR (NOT (fsm_output(4))) OR (fsm_output(2))
      OR mux_1696_nl);
  mux_1698_nl <= MUX_s_1_2_2(nor_1067_nl, nor_1068_nl, fsm_output(8));
  or_1578_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(7)) OR (fsm_output(9)) OR not_tmp_248;
  or_1576_nl <= (NOT (fsm_output(7))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1001")) OR (NOT (fsm_output(9))) OR (fsm_output(5))
      OR (fsm_output(10));
  mux_1693_nl <= MUX_s_1_2_2(or_1578_nl, or_1576_nl, fsm_output(2));
  mux_1694_nl <= MUX_s_1_2_2(mux_1693_nl, mux_tmp_1692, fsm_output(4));
  nor_1069_nl <= NOT((fsm_output(8)) OR (fsm_output(6)) OR mux_1694_nl);
  mux_1699_nl <= MUX_s_1_2_2(mux_1698_nl, nor_1069_nl, fsm_output(0));
  or_1571_nl <= CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (fsm_output(2)) OR (NOT (fsm_output(7))) OR (NOT (VEC_LOOP_j_sva_11_0(0)))
      OR (fsm_output(9)) OR (fsm_output(5)) OR (NOT (fsm_output(10)));
  or_1569_nl <= (fsm_output(2)) OR (NOT (fsm_output(7))) OR (NOT (fsm_output(9)))
      OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("1001")) OR (fsm_output(10));
  mux_1689_nl <= MUX_s_1_2_2(or_1571_nl, or_1569_nl, fsm_output(4));
  or_1568_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(7))) OR (NOT (VEC_LOOP_j_sva_11_0(0)))
      OR (NOT (fsm_output(9))) OR (NOT (fsm_output(5))) OR (fsm_output(10));
  or_1567_nl <= (NOT (fsm_output(2))) OR (NOT (fsm_output(7))) OR (fsm_output(9))
      OR (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("1001")) OR (fsm_output(10));
  mux_1688_nl <= MUX_s_1_2_2(or_1568_nl, or_1567_nl, fsm_output(4));
  mux_1690_nl <= MUX_s_1_2_2(mux_1689_nl, mux_1688_nl, fsm_output(6));
  nor_1070_nl <= NOT((fsm_output(8)) OR mux_1690_nl);
  nor_1071_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT (fsm_output(6))) OR (fsm_output(4)) OR (fsm_output(2)) OR (NOT (fsm_output(7)))
      OR (fsm_output(9)) OR (NOT (fsm_output(5))) OR (fsm_output(10)));
  nor_1072_nl <= NOT((NOT (fsm_output(4))) OR (NOT (fsm_output(2))) OR (NOT (fsm_output(7)))
      OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(9)) OR not_tmp_248);
  or_1562_nl <= (fsm_output(7)) OR (fsm_output(9)) OR (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001")) OR not_tmp_318;
  or_1560_nl <= (NOT (fsm_output(7))) OR (NOT (fsm_output(9))) OR (fsm_output(5))
      OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(10));
  mux_1685_nl <= MUX_s_1_2_2(or_1562_nl, or_1560_nl, fsm_output(2));
  nor_1073_nl <= NOT((fsm_output(4)) OR mux_1685_nl);
  mux_1686_nl <= MUX_s_1_2_2(nor_1072_nl, nor_1073_nl, fsm_output(6));
  mux_1687_nl <= MUX_s_1_2_2(nor_1071_nl, mux_1686_nl, fsm_output(8));
  mux_1691_nl <= MUX_s_1_2_2(nor_1070_nl, mux_1687_nl, fsm_output(0));
  mux_1700_nl <= MUX_s_1_2_2(mux_1699_nl, mux_1691_nl, fsm_output(3));
  vec_rsc_0_9_i_wea_d_pff <= MUX_s_1_2_2(mux_1714_nl, mux_1700_nl, fsm_output(1));
  or_1669_nl <= (NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(2))) OR (fsm_output(10));
  or_1668_nl <= (fsm_output(7)) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(2)) OR (NOT (fsm_output(10)));
  mux_1745_nl <= MUX_s_1_2_2(or_1669_nl, or_1668_nl, fsm_output(5));
  nor_1028_nl <= NOT((fsm_output(1)) OR mux_1745_nl);
  nor_1029_nl <= NOT((fsm_output(5)) OR (NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1001")) OR (fsm_output(3)) OR (fsm_output(9))
      OR (fsm_output(2)) OR (fsm_output(10)));
  nor_1030_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT (fsm_output(7))) OR (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_253);
  nor_1031_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(7)) OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (fsm_output(2))
      OR (NOT (fsm_output(10))));
  mux_1743_nl <= MUX_s_1_2_2(nor_1030_nl, nor_1031_nl, fsm_output(5));
  mux_1744_nl <= MUX_s_1_2_2(nor_1029_nl, mux_1743_nl, fsm_output(1));
  mux_1746_nl <= MUX_s_1_2_2(nor_1028_nl, mux_1744_nl, fsm_output(0));
  and_585_nl <= (fsm_output(6)) AND mux_1746_nl;
  nor_1032_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR (fsm_output(2)) OR (fsm_output(10)));
  nor_1034_nl <= NOT((fsm_output(7)) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR not_tmp_253);
  mux_1738_nl <= MUX_s_1_2_2(nor_1445_cse, nor_1034_nl, fsm_output(5));
  nor_1035_nl <= NOT((NOT (fsm_output(5))) OR (fsm_output(7)) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1001")) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR not_tmp_253);
  or_1655_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm);
  mux_1739_nl <= MUX_s_1_2_2(mux_1738_nl, nor_1035_nl, or_1655_nl);
  mux_1740_nl <= MUX_s_1_2_2(nor_1032_nl, mux_1739_nl, fsm_output(1));
  nor_1036_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR
      (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_253);
  nor_1037_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (NOT
      (fsm_output(2))) OR (fsm_output(10)));
  nor_1038_nl <= NOT((fsm_output(7)) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9))) OR (fsm_output(2)) OR (fsm_output(10)));
  mux_1736_nl <= MUX_s_1_2_2(nor_1037_nl, nor_1038_nl, fsm_output(5));
  mux_1737_nl <= MUX_s_1_2_2(nor_1036_nl, mux_1736_nl, fsm_output(1));
  mux_1741_nl <= MUX_s_1_2_2(mux_1740_nl, mux_1737_nl, fsm_output(0));
  nor_1039_nl <= NOT((NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (NOT (fsm_output(5)))
      OR (fsm_output(7)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR not_tmp_253);
  nor_1040_nl <= NOT((NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (NOT (fsm_output(5)))
      OR (fsm_output(7)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(3)) OR (fsm_output(9)) OR (NOT (fsm_output(2))) OR (fsm_output(10)));
  mux_1734_nl <= MUX_s_1_2_2(nor_1039_nl, nor_1040_nl, fsm_output(1));
  nor_1041_nl <= NOT((fsm_output(1)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO
      0)/=STD_LOGIC_VECTOR'("01")) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR mux_1669_cse);
  mux_1735_nl <= MUX_s_1_2_2(mux_1734_nl, nor_1041_nl, fsm_output(0));
  mux_1742_nl <= MUX_s_1_2_2(mux_1741_nl, mux_1735_nl, fsm_output(6));
  mux_1747_nl <= MUX_s_1_2_2(and_585_nl, mux_1742_nl, fsm_output(8));
  nor_1042_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (fsm_output(2))
      OR (fsm_output(10)));
  nor_1043_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(7)) OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(2)))
      OR (fsm_output(10)));
  mux_1728_nl <= MUX_s_1_2_2(nor_1042_nl, nor_1043_nl, fsm_output(5));
  and_586_nl <= COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm AND mux_1728_nl;
  nor_1044_nl <= NOT((NOT (fsm_output(7))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1001")) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR not_tmp_253);
  nor_1045_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(7)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9))) OR (fsm_output(2))
      OR (NOT (fsm_output(10))));
  mux_1727_nl <= MUX_s_1_2_2(nor_1044_nl, nor_1045_nl, fsm_output(5));
  and_587_nl <= COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm AND mux_1727_nl;
  mux_1729_nl <= MUX_s_1_2_2(and_586_nl, and_587_nl, fsm_output(1));
  nor_1046_nl <= NOT((NOT (VEC_LOOP_j_sva_11_0(3))) OR (VEC_LOOP_j_sva_11_0(1)) OR
      (NOT (VEC_LOOP_j_sva_11_0(0))) OR (NOT (fsm_output(5))) OR (VEC_LOOP_j_sva_11_0(2))
      OR (fsm_output(7)) OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(2))
      OR (fsm_output(10)));
  nor_1047_nl <= NOT(nand_332_cse OR mux_1661_cse);
  mux_1726_nl <= MUX_s_1_2_2(nor_1046_nl, nor_1047_nl, fsm_output(1));
  mux_1730_nl <= MUX_s_1_2_2(mux_1729_nl, mux_1726_nl, fsm_output(0));
  nor_1048_nl <= NOT((NOT (fsm_output(1))) OR (fsm_output(5)) OR (fsm_output(7))
      OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001")) OR (NOT
      (fsm_output(3))) OR (fsm_output(9)) OR (fsm_output(2)) OR (fsm_output(10)));
  nor_1049_nl <= NOT((fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(3)))
      OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001")) OR (NOT
      (fsm_output(9))) OR (NOT (fsm_output(2))) OR (fsm_output(10)));
  nor_1050_nl <= NOT((NOT (VEC_LOOP_j_sva_11_0(0))) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (NOT
      (fsm_output(2))) OR (fsm_output(10)));
  mux_1723_nl <= MUX_s_1_2_2(nor_1049_nl, nor_1050_nl, fsm_output(1));
  mux_1724_nl <= MUX_s_1_2_2(nor_1048_nl, mux_1723_nl, fsm_output(0));
  mux_1731_nl <= MUX_s_1_2_2(mux_1730_nl, mux_1724_nl, fsm_output(6));
  nor_1051_nl <= NOT((NOT (fsm_output(1))) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(3)) OR (NOT (fsm_output(9)))
      OR (fsm_output(2)) OR (fsm_output(10)));
  nor_1052_nl <= NOT((fsm_output(1)) OR (fsm_output(5)) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1001")) OR (NOT (fsm_output(7))) OR (fsm_output(3))
      OR (fsm_output(9)) OR not_tmp_253);
  mux_1721_nl <= MUX_s_1_2_2(nor_1051_nl, nor_1052_nl, fsm_output(0));
  nor_1053_nl <= NOT((NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1001")) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR not_tmp_253);
  nor_1054_nl <= NOT((NOT (fsm_output(7))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1001")) OR (fsm_output(3)) OR (NOT (fsm_output(9)))
      OR (fsm_output(2)) OR (fsm_output(10)));
  nor_1055_nl <= NOT((NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR not_tmp_253);
  mux_1717_nl <= MUX_s_1_2_2(nor_1054_nl, nor_1055_nl, fsm_output(5));
  mux_1718_nl <= MUX_s_1_2_2(nor_1053_nl, mux_1717_nl, COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm);
  nor_1056_nl <= NOT((NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1001")) OR (fsm_output(3)) OR (fsm_output(9))
      OR (NOT (fsm_output(2))) OR (fsm_output(10)));
  mux_1719_nl <= MUX_s_1_2_2(mux_1718_nl, nor_1056_nl, fsm_output(1));
  nor_1057_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3)))
      OR (NOT (fsm_output(9))) OR (fsm_output(2)) OR (fsm_output(10)));
  nor_1058_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(3)) OR (fsm_output(9))
      OR (fsm_output(2)) OR (NOT (fsm_output(10))));
  mux_1716_nl <= MUX_s_1_2_2(nor_1057_nl, nor_1058_nl, fsm_output(1));
  mux_1720_nl <= MUX_s_1_2_2(mux_1719_nl, mux_1716_nl, fsm_output(0));
  mux_1722_nl <= MUX_s_1_2_2(mux_1721_nl, mux_1720_nl, fsm_output(6));
  mux_1732_nl <= MUX_s_1_2_2(mux_1731_nl, mux_1722_nl, fsm_output(8));
  vec_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_1747_nl, mux_1732_nl,
      fsm_output(4));
  or_1723_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (NOT (VEC_LOOP_j_sva_11_0(1))) OR (NOT (fsm_output(5))) OR (VEC_LOOP_j_sva_11_0(0))
      OR CONV_SL_1_1(fsm_output(10 DOWNTO 9)/=STD_LOGIC_VECTOR'("01"));
  or_1722_nl <= (NOT (fsm_output(5))) OR (NOT (fsm_output(9))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010")) OR not_tmp_318;
  mux_1774_nl <= MUX_s_1_2_2(or_1723_nl, or_1722_nl, fsm_output(7));
  or_1720_nl <= CONV_SL_1_1(VEC_LOOP_j_sva_11_0(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("10"))
      OR (NOT (fsm_output(7))) OR (NOT (VEC_LOOP_j_sva_11_0(1))) OR (fsm_output(5))
      OR (VEC_LOOP_j_sva_11_0(0)) OR CONV_SL_1_1(fsm_output(10 DOWNTO 9)/=STD_LOGIC_VECTOR'("00"));
  mux_1775_nl <= MUX_s_1_2_2(mux_1774_nl, or_1720_nl, fsm_output(2));
  nor_1013_nl <= NOT((fsm_output(6)) OR (fsm_output(4)) OR mux_1775_nl);
  nor_1014_nl <= NOT((fsm_output(6)) OR (fsm_output(4)) OR (NOT (fsm_output(2)))
      OR (fsm_output(7)) OR (fsm_output(5)) OR (fsm_output(9)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010")) OR not_tmp_318);
  mux_1776_nl <= MUX_s_1_2_2(nor_1013_nl, nor_1014_nl, fsm_output(8));
  nor_1015_nl <= NOT((NOT (fsm_output(6))) OR (NOT (fsm_output(4))) OR (fsm_output(2))
      OR (NOT (fsm_output(7))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("1010")) OR (NOT (fsm_output(5))) OR (fsm_output(9))
      OR (NOT (fsm_output(10))));
  nor_1016_nl <= NOT((fsm_output(4)) OR (fsm_output(2)) OR (fsm_output(7)) OR (fsm_output(5))
      OR (NOT (fsm_output(9))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("1010")) OR (fsm_output(10)));
  nor_1017_nl <= NOT((NOT (fsm_output(2))) OR (fsm_output(7)) OR (NOT (fsm_output(5)))
      OR (fsm_output(9)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("1010")) OR (fsm_output(10)));
  nor_1018_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT (fsm_output(2))) OR (fsm_output(7)) OR (fsm_output(5)) OR (NOT (fsm_output(9)))
      OR (fsm_output(10)));
  mux_1771_nl <= MUX_s_1_2_2(nor_1017_nl, nor_1018_nl, fsm_output(4));
  mux_1772_nl <= MUX_s_1_2_2(nor_1016_nl, mux_1771_nl, fsm_output(6));
  mux_1773_nl <= MUX_s_1_2_2(nor_1015_nl, mux_1772_nl, fsm_output(8));
  mux_1777_nl <= MUX_s_1_2_2(mux_1776_nl, mux_1773_nl, fsm_output(0));
  nand_282_nl <= NOT((COMP_LOOP_acc_16_psp_sva(0)) AND (fsm_output(4)) AND (fsm_output(2))
      AND (NOT (VEC_LOOP_j_sva_11_0(2))) AND (fsm_output(7)) AND (VEC_LOOP_j_sva_11_0(1))
      AND (fsm_output(5)) AND (NOT (VEC_LOOP_j_sva_11_0(0))) AND CONV_SL_1_1(fsm_output(10
      DOWNTO 9)=STD_LOGIC_VECTOR'("01")));
  or_1710_nl <= CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (fsm_output(2)) OR (fsm_output(7)) OR (NOT (VEC_LOOP_j_sva_11_0(1))) OR
      (fsm_output(5)) OR (VEC_LOOP_j_sva_11_0(0)) OR CONV_SL_1_1(fsm_output(10 DOWNTO
      9)/=STD_LOGIC_VECTOR'("10"));
  mux_1768_nl <= MUX_s_1_2_2(mux_tmp_1756, or_1710_nl, fsm_output(4));
  mux_1769_nl <= MUX_s_1_2_2(nand_282_nl, mux_1768_nl, fsm_output(6));
  and_584_nl <= (fsm_output(8)) AND (NOT mux_1769_nl);
  or_1707_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(7))) OR (fsm_output(5)) OR nand_358_cse;
  or_1705_nl <= (fsm_output(7)) OR (NOT (fsm_output(5))) OR (NOT (fsm_output(9)))
      OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR not_tmp_318;
  mux_1765_nl <= MUX_s_1_2_2(or_1705_nl, or_tmp_1640, fsm_output(2));
  mux_1766_nl <= MUX_s_1_2_2(or_1707_nl, mux_1765_nl, fsm_output(4));
  nor_1019_nl <= NOT((fsm_output(6)) OR mux_1766_nl);
  nor_1020_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(6)) OR (NOT (fsm_output(4))) OR (fsm_output(2)) OR (NOT (fsm_output(7)))
      OR (NOT (fsm_output(5))) OR (fsm_output(9)) OR (fsm_output(10)));
  mux_1767_nl <= MUX_s_1_2_2(nor_1019_nl, nor_1020_nl, fsm_output(8));
  mux_1770_nl <= MUX_s_1_2_2(and_584_nl, mux_1767_nl, fsm_output(0));
  mux_1778_nl <= MUX_s_1_2_2(mux_1777_nl, mux_1770_nl, fsm_output(3));
  or_1701_nl <= CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (NOT (fsm_output(2))) OR (fsm_output(7)) OR (NOT (fsm_output(5))) OR (VEC_LOOP_j_sva_11_0(0))
      OR nand_358_cse;
  or_1699_nl <= (NOT (fsm_output(2))) OR (fsm_output(7)) OR (NOT (fsm_output(5)))
      OR (fsm_output(9)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(2 DOWNTO
      0)/=STD_LOGIC_VECTOR'("010")) OR not_tmp_318;
  mux_1761_nl <= MUX_s_1_2_2(or_1701_nl, or_1699_nl, fsm_output(4));
  nor_1021_nl <= NOT((fsm_output(6)) OR mux_1761_nl);
  or_1693_nl <= (fsm_output(5)) OR (fsm_output(9)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010")) OR not_tmp_318;
  mux_1759_nl <= MUX_s_1_2_2(or_591_cse, or_1693_nl, fsm_output(7));
  mux_1760_nl <= MUX_s_1_2_2(or_tmp_1640, mux_1759_nl, nor_239_cse);
  nor_1022_nl <= NOT((NOT (fsm_output(6))) OR (NOT (fsm_output(4))) OR (fsm_output(2))
      OR mux_1760_nl);
  mux_1762_nl <= MUX_s_1_2_2(nor_1021_nl, nor_1022_nl, fsm_output(8));
  or_1689_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(7)) OR (NOT (fsm_output(5))) OR (fsm_output(9)) OR (NOT (fsm_output(10)));
  or_1687_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT (fsm_output(7))) OR (fsm_output(5)) OR (NOT (fsm_output(9))) OR (fsm_output(10));
  mux_1757_nl <= MUX_s_1_2_2(or_1689_nl, or_1687_nl, fsm_output(2));
  mux_1758_nl <= MUX_s_1_2_2(mux_1757_nl, mux_tmp_1756, fsm_output(4));
  nor_1023_nl <= NOT((fsm_output(8)) OR (fsm_output(6)) OR mux_1758_nl);
  mux_1763_nl <= MUX_s_1_2_2(mux_1762_nl, nor_1023_nl, fsm_output(0));
  or_1682_nl <= CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (fsm_output(2)) OR (NOT (fsm_output(7))) OR (fsm_output(5)) OR (VEC_LOOP_j_sva_11_0(0))
      OR CONV_SL_1_1(fsm_output(10 DOWNTO 9)/=STD_LOGIC_VECTOR'("10"));
  or_1680_nl <= (fsm_output(2)) OR (NOT (fsm_output(7))) OR (fsm_output(5)) OR (NOT
      (fsm_output(9))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(10));
  mux_1753_nl <= MUX_s_1_2_2(or_1682_nl, or_1680_nl, fsm_output(4));
  or_1679_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(7))) OR (NOT (fsm_output(5)))
      OR (VEC_LOOP_j_sva_11_0(0)) OR CONV_SL_1_1(fsm_output(10 DOWNTO 9)/=STD_LOGIC_VECTOR'("01"));
  or_1678_nl <= (NOT (fsm_output(2))) OR (NOT (fsm_output(7))) OR (NOT (fsm_output(5)))
      OR (fsm_output(9)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("1010")) OR (fsm_output(10));
  mux_1752_nl <= MUX_s_1_2_2(or_1679_nl, or_1678_nl, fsm_output(4));
  mux_1754_nl <= MUX_s_1_2_2(mux_1753_nl, mux_1752_nl, fsm_output(6));
  nor_1024_nl <= NOT((fsm_output(8)) OR mux_1754_nl);
  nor_1025_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT (fsm_output(6))) OR (fsm_output(4)) OR (fsm_output(2)) OR (NOT (fsm_output(7)))
      OR (NOT (fsm_output(5))) OR (fsm_output(9)) OR (fsm_output(10)));
  and_761_nl <= (fsm_output(4)) AND (fsm_output(2)) AND (fsm_output(7)) AND CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3
      DOWNTO 0)=STD_LOGIC_VECTOR'("1010")) AND (fsm_output(5)) AND (NOT (fsm_output(9)))
      AND (fsm_output(10));
  or_1673_nl <= (fsm_output(7)) OR (NOT (fsm_output(5))) OR (fsm_output(9)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010")) OR not_tmp_318;
  or_1671_nl <= (NOT (fsm_output(7))) OR (fsm_output(5)) OR (NOT (fsm_output(9)))
      OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(10));
  mux_1749_nl <= MUX_s_1_2_2(or_1673_nl, or_1671_nl, fsm_output(2));
  nor_1027_nl <= NOT((fsm_output(4)) OR mux_1749_nl);
  mux_1750_nl <= MUX_s_1_2_2(and_761_nl, nor_1027_nl, fsm_output(6));
  mux_1751_nl <= MUX_s_1_2_2(nor_1025_nl, mux_1750_nl, fsm_output(8));
  mux_1755_nl <= MUX_s_1_2_2(nor_1024_nl, mux_1751_nl, fsm_output(0));
  mux_1764_nl <= MUX_s_1_2_2(mux_1763_nl, mux_1755_nl, fsm_output(3));
  vec_rsc_0_10_i_wea_d_pff <= MUX_s_1_2_2(mux_1778_nl, mux_1764_nl, fsm_output(1));
  or_1779_nl <= (NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(2))) OR (fsm_output(10));
  or_1778_nl <= (fsm_output(7)) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(2)) OR (NOT (fsm_output(10)));
  mux_1809_nl <= MUX_s_1_2_2(or_1779_nl, or_1778_nl, fsm_output(5));
  nor_982_nl <= NOT((fsm_output(1)) OR mux_1809_nl);
  nor_983_nl <= NOT((fsm_output(5)) OR (NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1010")) OR (fsm_output(3)) OR (fsm_output(9))
      OR (fsm_output(2)) OR (fsm_output(10)));
  nor_984_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT (fsm_output(7))) OR (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_253);
  nor_985_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(7)) OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (fsm_output(2))
      OR (NOT (fsm_output(10))));
  mux_1807_nl <= MUX_s_1_2_2(nor_984_nl, nor_985_nl, fsm_output(5));
  mux_1808_nl <= MUX_s_1_2_2(nor_983_nl, mux_1807_nl, fsm_output(1));
  mux_1810_nl <= MUX_s_1_2_2(nor_982_nl, mux_1808_nl, fsm_output(0));
  and_581_nl <= (fsm_output(6)) AND mux_1810_nl;
  nor_986_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR (fsm_output(2)) OR (fsm_output(10)));
  nor_988_nl <= NOT((fsm_output(7)) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR not_tmp_253);
  mux_1802_nl <= MUX_s_1_2_2(nor_1445_cse, nor_988_nl, fsm_output(5));
  nor_989_nl <= NOT((NOT (fsm_output(5))) OR (fsm_output(7)) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1010")) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR not_tmp_253);
  or_1765_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm);
  mux_1803_nl <= MUX_s_1_2_2(mux_1802_nl, nor_989_nl, or_1765_nl);
  mux_1804_nl <= MUX_s_1_2_2(nor_986_nl, mux_1803_nl, fsm_output(1));
  nor_990_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR
      (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_253);
  nor_991_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (NOT
      (fsm_output(2))) OR (fsm_output(10)));
  nor_992_nl <= NOT((fsm_output(7)) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9))) OR (fsm_output(2)) OR (fsm_output(10)));
  mux_1800_nl <= MUX_s_1_2_2(nor_991_nl, nor_992_nl, fsm_output(5));
  mux_1801_nl <= MUX_s_1_2_2(nor_990_nl, mux_1800_nl, fsm_output(1));
  mux_1805_nl <= MUX_s_1_2_2(mux_1804_nl, mux_1801_nl, fsm_output(0));
  nor_993_nl <= NOT((NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (NOT (fsm_output(5)))
      OR (fsm_output(7)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR not_tmp_253);
  nor_994_nl <= NOT((NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (NOT (fsm_output(5)))
      OR (fsm_output(7)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(3)) OR (fsm_output(9)) OR (NOT (fsm_output(2))) OR (fsm_output(10)));
  mux_1798_nl <= MUX_s_1_2_2(nor_993_nl, nor_994_nl, fsm_output(1));
  nor_995_nl <= NOT((fsm_output(1)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR mux_1669_cse);
  mux_1799_nl <= MUX_s_1_2_2(mux_1798_nl, nor_995_nl, fsm_output(0));
  mux_1806_nl <= MUX_s_1_2_2(mux_1805_nl, mux_1799_nl, fsm_output(6));
  mux_1811_nl <= MUX_s_1_2_2(and_581_nl, mux_1806_nl, fsm_output(8));
  nor_996_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (fsm_output(2))
      OR (fsm_output(10)));
  nor_997_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(7)) OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(2)))
      OR (fsm_output(10)));
  mux_1792_nl <= MUX_s_1_2_2(nor_996_nl, nor_997_nl, fsm_output(5));
  and_582_nl <= COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm AND mux_1792_nl;
  nor_998_nl <= NOT((NOT (fsm_output(7))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1010")) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR not_tmp_253);
  nor_999_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(7)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9))) OR (fsm_output(2))
      OR (NOT (fsm_output(10))));
  mux_1791_nl <= MUX_s_1_2_2(nor_998_nl, nor_999_nl, fsm_output(5));
  and_583_nl <= COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm AND mux_1791_nl;
  mux_1793_nl <= MUX_s_1_2_2(and_582_nl, and_583_nl, fsm_output(1));
  nor_1000_nl <= NOT((NOT (VEC_LOOP_j_sva_11_0(3))) OR (NOT (VEC_LOOP_j_sva_11_0(1)))
      OR (VEC_LOOP_j_sva_11_0(0)) OR (NOT (fsm_output(5))) OR (VEC_LOOP_j_sva_11_0(2))
      OR (fsm_output(7)) OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(2))
      OR (fsm_output(10)));
  nor_1001_nl <= NOT((VEC_LOOP_j_sva_11_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR mux_1789_cse);
  mux_1790_nl <= MUX_s_1_2_2(nor_1000_nl, nor_1001_nl, fsm_output(1));
  mux_1794_nl <= MUX_s_1_2_2(mux_1793_nl, mux_1790_nl, fsm_output(0));
  nor_1002_nl <= NOT((NOT (fsm_output(1))) OR (fsm_output(5)) OR (fsm_output(7))
      OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010")) OR (NOT
      (fsm_output(3))) OR (fsm_output(9)) OR (fsm_output(2)) OR (fsm_output(10)));
  nor_1003_nl <= NOT((fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(3)))
      OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010")) OR (NOT
      (fsm_output(9))) OR (NOT (fsm_output(2))) OR (fsm_output(10)));
  nor_1004_nl <= NOT((VEC_LOOP_j_sva_11_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (NOT
      (fsm_output(2))) OR (fsm_output(10)));
  mux_1787_nl <= MUX_s_1_2_2(nor_1003_nl, nor_1004_nl, fsm_output(1));
  mux_1788_nl <= MUX_s_1_2_2(nor_1002_nl, mux_1787_nl, fsm_output(0));
  mux_1795_nl <= MUX_s_1_2_2(mux_1794_nl, mux_1788_nl, fsm_output(6));
  nor_1005_nl <= NOT((NOT (fsm_output(1))) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(3)) OR (NOT (fsm_output(9)))
      OR (fsm_output(2)) OR (fsm_output(10)));
  nor_1006_nl <= NOT((fsm_output(1)) OR (fsm_output(5)) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1010")) OR (NOT (fsm_output(7))) OR (fsm_output(3))
      OR (fsm_output(9)) OR not_tmp_253);
  mux_1785_nl <= MUX_s_1_2_2(nor_1005_nl, nor_1006_nl, fsm_output(0));
  nor_1007_nl <= NOT((NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1010")) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR not_tmp_253);
  nor_1008_nl <= NOT((NOT (fsm_output(7))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1010")) OR (fsm_output(3)) OR (NOT (fsm_output(9)))
      OR (fsm_output(2)) OR (fsm_output(10)));
  nor_1009_nl <= NOT((NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR not_tmp_253);
  mux_1781_nl <= MUX_s_1_2_2(nor_1008_nl, nor_1009_nl, fsm_output(5));
  mux_1782_nl <= MUX_s_1_2_2(nor_1007_nl, mux_1781_nl, COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm);
  nor_1010_nl <= NOT((NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1010")) OR (fsm_output(3)) OR (fsm_output(9))
      OR (NOT (fsm_output(2))) OR (fsm_output(10)));
  mux_1783_nl <= MUX_s_1_2_2(mux_1782_nl, nor_1010_nl, fsm_output(1));
  nor_1011_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3)))
      OR (NOT (fsm_output(9))) OR (fsm_output(2)) OR (fsm_output(10)));
  nor_1012_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (VEC_LOOP_j_sva_11_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR
      (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(3)) OR (fsm_output(9))
      OR (fsm_output(2)) OR (NOT (fsm_output(10))));
  mux_1780_nl <= MUX_s_1_2_2(nor_1011_nl, nor_1012_nl, fsm_output(1));
  mux_1784_nl <= MUX_s_1_2_2(mux_1783_nl, mux_1780_nl, fsm_output(0));
  mux_1786_nl <= MUX_s_1_2_2(mux_1785_nl, mux_1784_nl, fsm_output(6));
  mux_1796_nl <= MUX_s_1_2_2(mux_1795_nl, mux_1786_nl, fsm_output(8));
  vec_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_1811_nl, mux_1796_nl,
      fsm_output(4));
  nand_272_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("10"))
      AND CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND
      (fsm_output(9)) AND (fsm_output(5)) AND (NOT (fsm_output(10))));
  or_1832_nl <= (NOT((fsm_output(9)) AND (fsm_output(5)) AND CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(2
      DOWNTO 0)=STD_LOGIC_VECTOR'("011")))) OR not_tmp_318;
  mux_1838_nl <= MUX_s_1_2_2(nand_272_nl, or_1832_nl, fsm_output(7));
  or_1830_nl <= CONV_SL_1_1(VEC_LOOP_j_sva_11_0(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("10"))
      OR (NOT (fsm_output(7))) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR (fsm_output(9)) OR (fsm_output(5)) OR (fsm_output(10));
  mux_1839_nl <= MUX_s_1_2_2(mux_1838_nl, or_1830_nl, fsm_output(2));
  nor_967_nl <= NOT((fsm_output(6)) OR (fsm_output(4)) OR mux_1839_nl);
  nor_968_nl <= NOT((fsm_output(6)) OR (fsm_output(4)) OR (NOT (fsm_output(2))) OR
      (fsm_output(7)) OR (fsm_output(9)) OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("011")) OR not_tmp_318);
  mux_1840_nl <= MUX_s_1_2_2(nor_967_nl, nor_968_nl, fsm_output(8));
  nor_969_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (NOT (fsm_output(6))) OR (NOT (fsm_output(4))) OR (fsm_output(2)) OR (NOT
      (fsm_output(7))) OR (fsm_output(9)) OR not_tmp_248);
  nor_970_nl <= NOT((fsm_output(4)) OR (fsm_output(2)) OR (fsm_output(7)) OR (NOT
      (fsm_output(9))) OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1011")) OR (fsm_output(10)));
  nor_971_nl <= NOT((NOT (fsm_output(2))) OR (fsm_output(7)) OR (fsm_output(9)) OR
      (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("1011")) OR (fsm_output(10)));
  nor_972_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (NOT (fsm_output(2))) OR (fsm_output(7)) OR (NOT (fsm_output(9))) OR (fsm_output(5))
      OR (fsm_output(10)));
  mux_1835_nl <= MUX_s_1_2_2(nor_971_nl, nor_972_nl, fsm_output(4));
  mux_1836_nl <= MUX_s_1_2_2(nor_970_nl, mux_1835_nl, fsm_output(6));
  mux_1837_nl <= MUX_s_1_2_2(nor_969_nl, mux_1836_nl, fsm_output(8));
  mux_1841_nl <= MUX_s_1_2_2(mux_1840_nl, mux_1837_nl, fsm_output(0));
  nand_274_nl <= NOT((COMP_LOOP_acc_16_psp_sva(0)) AND (fsm_output(4)) AND (fsm_output(2))
      AND (NOT (VEC_LOOP_j_sva_11_0(2))) AND (fsm_output(7)) AND CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1
      DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND (fsm_output(9)) AND (fsm_output(5))
      AND (NOT (fsm_output(10))));
  or_1820_nl <= CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (fsm_output(2)) OR (fsm_output(7)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("11")) OR (fsm_output(9)) OR (fsm_output(5)) OR
      (NOT (fsm_output(10)));
  mux_1832_nl <= MUX_s_1_2_2(mux_tmp_1820, or_1820_nl, fsm_output(4));
  mux_1833_nl <= MUX_s_1_2_2(nand_274_nl, mux_1832_nl, fsm_output(6));
  and_580_nl <= (fsm_output(8)) AND (NOT mux_1833_nl);
  nand_398_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1011"))
      AND (fsm_output(2)) AND (fsm_output(7)) AND (fsm_output(9)) AND (NOT (fsm_output(5)))
      AND (fsm_output(10)));
  or_1815_nl <= (fsm_output(7)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(5)))
      OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR not_tmp_318;
  mux_1829_nl <= MUX_s_1_2_2(or_1815_nl, or_tmp_1750, fsm_output(2));
  mux_1830_nl <= MUX_s_1_2_2(nand_398_nl, mux_1829_nl, fsm_output(4));
  nor_973_nl <= NOT((fsm_output(6)) OR mux_1830_nl);
  nor_974_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(6)) OR (NOT (fsm_output(4))) OR (fsm_output(2)) OR (NOT (fsm_output(7)))
      OR (fsm_output(9)) OR (NOT (fsm_output(5))) OR (fsm_output(10)));
  mux_1831_nl <= MUX_s_1_2_2(nor_973_nl, nor_974_nl, fsm_output(8));
  mux_1834_nl <= MUX_s_1_2_2(and_580_nl, mux_1831_nl, fsm_output(0));
  mux_1842_nl <= MUX_s_1_2_2(mux_1841_nl, mux_1834_nl, fsm_output(3));
  or_1811_nl <= CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (NOT (fsm_output(2))) OR (fsm_output(7)) OR nand_334_cse;
  or_1809_nl <= (NOT (fsm_output(2))) OR (fsm_output(7)) OR (fsm_output(9)) OR (NOT
      (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR not_tmp_318;
  mux_1825_nl <= MUX_s_1_2_2(or_1811_nl, or_1809_nl, fsm_output(4));
  nor_975_nl <= NOT((fsm_output(6)) OR mux_1825_nl);
  or_1803_nl <= (fsm_output(9)) OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("011")) OR not_tmp_318;
  mux_1823_nl <= MUX_s_1_2_2(or_702_cse, or_1803_nl, fsm_output(7));
  mux_1824_nl <= MUX_s_1_2_2(or_tmp_1750, mux_1823_nl, nor_239_cse);
  nor_976_nl <= NOT((NOT (fsm_output(6))) OR (NOT (fsm_output(4))) OR (fsm_output(2))
      OR mux_1824_nl);
  mux_1826_nl <= MUX_s_1_2_2(nor_975_nl, nor_976_nl, fsm_output(8));
  or_1799_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(7)) OR (fsm_output(9)) OR not_tmp_248;
  or_1797_nl <= (NOT (fsm_output(7))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1011")) OR (NOT (fsm_output(9))) OR (fsm_output(5))
      OR (fsm_output(10));
  mux_1821_nl <= MUX_s_1_2_2(or_1799_nl, or_1797_nl, fsm_output(2));
  mux_1822_nl <= MUX_s_1_2_2(mux_1821_nl, mux_tmp_1820, fsm_output(4));
  nor_977_nl <= NOT((fsm_output(8)) OR (fsm_output(6)) OR mux_1822_nl);
  mux_1827_nl <= MUX_s_1_2_2(mux_1826_nl, nor_977_nl, fsm_output(0));
  or_1792_nl <= CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (fsm_output(2)) OR (NOT (fsm_output(7))) OR (NOT (VEC_LOOP_j_sva_11_0(0)))
      OR (fsm_output(9)) OR (fsm_output(5)) OR (NOT (fsm_output(10)));
  or_1790_nl <= (fsm_output(2)) OR (NOT (fsm_output(7))) OR (NOT (fsm_output(9)))
      OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("1011")) OR (fsm_output(10));
  mux_1817_nl <= MUX_s_1_2_2(or_1792_nl, or_1790_nl, fsm_output(4));
  nand_277_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("101"))
      AND (fsm_output(2)) AND (fsm_output(7)) AND (VEC_LOOP_j_sva_11_0(0)) AND (fsm_output(9))
      AND (fsm_output(5)) AND (NOT (fsm_output(10))));
  or_1788_nl <= (NOT (fsm_output(2))) OR (NOT (fsm_output(7))) OR (fsm_output(9))
      OR (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("1011")) OR (fsm_output(10));
  mux_1816_nl <= MUX_s_1_2_2(nand_277_nl, or_1788_nl, fsm_output(4));
  mux_1818_nl <= MUX_s_1_2_2(mux_1817_nl, mux_1816_nl, fsm_output(6));
  nor_978_nl <= NOT((fsm_output(8)) OR mux_1818_nl);
  nor_979_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (NOT (fsm_output(6))) OR (fsm_output(4)) OR (fsm_output(2)) OR (NOT (fsm_output(7)))
      OR (fsm_output(9)) OR (NOT (fsm_output(5))) OR (fsm_output(10)));
  nor_980_nl <= NOT((NOT((fsm_output(4)) AND (fsm_output(2)) AND (fsm_output(7))
      AND CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1011"))
      AND (NOT (fsm_output(9))))) OR not_tmp_248);
  or_1783_nl <= (fsm_output(7)) OR (fsm_output(9)) OR (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("011")) OR not_tmp_318;
  or_1781_nl <= (NOT (fsm_output(7))) OR (NOT (fsm_output(9))) OR (fsm_output(5))
      OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(10));
  mux_1813_nl <= MUX_s_1_2_2(or_1783_nl, or_1781_nl, fsm_output(2));
  nor_981_nl <= NOT((fsm_output(4)) OR mux_1813_nl);
  mux_1814_nl <= MUX_s_1_2_2(nor_980_nl, nor_981_nl, fsm_output(6));
  mux_1815_nl <= MUX_s_1_2_2(nor_979_nl, mux_1814_nl, fsm_output(8));
  mux_1819_nl <= MUX_s_1_2_2(nor_978_nl, mux_1815_nl, fsm_output(0));
  mux_1828_nl <= MUX_s_1_2_2(mux_1827_nl, mux_1819_nl, fsm_output(3));
  vec_rsc_0_11_i_wea_d_pff <= MUX_s_1_2_2(mux_1842_nl, mux_1828_nl, fsm_output(1));
  or_1889_nl <= (NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(2))) OR (fsm_output(10));
  or_1888_nl <= (fsm_output(7)) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(2)) OR (NOT (fsm_output(10)));
  mux_1873_nl <= MUX_s_1_2_2(or_1889_nl, or_1888_nl, fsm_output(5));
  nor_938_nl <= NOT((fsm_output(1)) OR mux_1873_nl);
  nor_939_nl <= NOT((fsm_output(5)) OR (NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1011")) OR (fsm_output(3)) OR (fsm_output(9))
      OR (fsm_output(2)) OR (fsm_output(10)));
  nor_940_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (NOT (fsm_output(7))) OR (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_253);
  nor_941_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(7)) OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (fsm_output(2))
      OR (NOT (fsm_output(10))));
  mux_1871_nl <= MUX_s_1_2_2(nor_940_nl, nor_941_nl, fsm_output(5));
  mux_1872_nl <= MUX_s_1_2_2(nor_939_nl, mux_1871_nl, fsm_output(1));
  mux_1874_nl <= MUX_s_1_2_2(nor_938_nl, mux_1872_nl, fsm_output(0));
  and_575_nl <= (fsm_output(6)) AND mux_1874_nl;
  nor_942_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR (fsm_output(2)) OR (fsm_output(10)));
  nor_944_nl <= NOT((fsm_output(7)) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR not_tmp_253);
  mux_1866_nl <= MUX_s_1_2_2(nor_1445_cse, nor_944_nl, fsm_output(5));
  nor_945_nl <= NOT((NOT (fsm_output(5))) OR (fsm_output(7)) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1011")) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR not_tmp_253);
  nand_265_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1011"))
      AND COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm);
  mux_1867_nl <= MUX_s_1_2_2(mux_1866_nl, nor_945_nl, nand_265_nl);
  mux_1868_nl <= MUX_s_1_2_2(nor_942_nl, mux_1867_nl, fsm_output(1));
  nor_946_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11")) OR
      (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_253);
  nor_947_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (NOT
      (fsm_output(2))) OR (fsm_output(10)));
  nor_948_nl <= NOT((fsm_output(7)) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9))) OR (fsm_output(2)) OR (fsm_output(10)));
  mux_1864_nl <= MUX_s_1_2_2(nor_947_nl, nor_948_nl, fsm_output(5));
  mux_1865_nl <= MUX_s_1_2_2(nor_946_nl, mux_1864_nl, fsm_output(1));
  mux_1869_nl <= MUX_s_1_2_2(mux_1868_nl, mux_1865_nl, fsm_output(0));
  nor_949_nl <= NOT((NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (NOT (fsm_output(5)))
      OR (fsm_output(7)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR not_tmp_253);
  nor_950_nl <= NOT((NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (NOT (fsm_output(5)))
      OR (fsm_output(7)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(3)) OR (fsm_output(9)) OR (NOT (fsm_output(2))) OR (fsm_output(10)));
  mux_1862_nl <= MUX_s_1_2_2(nor_949_nl, nor_950_nl, fsm_output(1));
  nor_951_nl <= NOT(nand_324_cse OR mux_1669_cse);
  mux_1863_nl <= MUX_s_1_2_2(mux_1862_nl, nor_951_nl, fsm_output(0));
  mux_1870_nl <= MUX_s_1_2_2(mux_1869_nl, mux_1863_nl, fsm_output(6));
  mux_1875_nl <= MUX_s_1_2_2(and_575_nl, mux_1870_nl, fsm_output(8));
  nor_952_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (fsm_output(2))
      OR (fsm_output(10)));
  nor_953_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(7)) OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(2)))
      OR (fsm_output(10)));
  mux_1856_nl <= MUX_s_1_2_2(nor_952_nl, nor_953_nl, fsm_output(5));
  and_576_nl <= COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm AND mux_1856_nl;
  nor_954_nl <= NOT((NOT((fsm_output(7)) AND CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3
      DOWNTO 0)=STD_LOGIC_VECTOR'("1011")) AND (fsm_output(3)) AND (NOT (fsm_output(9)))))
      OR not_tmp_253);
  nor_955_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(7)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9))) OR (fsm_output(2))
      OR (NOT (fsm_output(10))));
  mux_1855_nl <= MUX_s_1_2_2(nor_954_nl, nor_955_nl, fsm_output(5));
  and_577_nl <= COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm AND mux_1855_nl;
  mux_1857_nl <= MUX_s_1_2_2(and_576_nl, and_577_nl, fsm_output(1));
  nor_956_nl <= NOT((NOT (VEC_LOOP_j_sva_11_0(3))) OR (NOT (VEC_LOOP_j_sva_11_0(1)))
      OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR (NOT (fsm_output(5))) OR (VEC_LOOP_j_sva_11_0(2))
      OR (fsm_output(7)) OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(2))
      OR (fsm_output(10)));
  nor_957_nl <= NOT(nand_332_cse OR mux_1789_cse);
  mux_1854_nl <= MUX_s_1_2_2(nor_956_nl, nor_957_nl, fsm_output(1));
  mux_1858_nl <= MUX_s_1_2_2(mux_1857_nl, mux_1854_nl, fsm_output(0));
  nor_958_nl <= NOT((NOT (fsm_output(1))) OR (fsm_output(5)) OR (fsm_output(7)) OR
      CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011")) OR (NOT (fsm_output(3)))
      OR (fsm_output(9)) OR (fsm_output(2)) OR (fsm_output(10)));
  nor_959_nl <= NOT((fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(3))) OR
      CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011")) OR (NOT (fsm_output(9)))
      OR (NOT (fsm_output(2))) OR (fsm_output(10)));
  and_578_nl <= (VEC_LOOP_j_sva_11_0(0)) AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm
      AND (fsm_output(5)) AND CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("101"))
      AND (fsm_output(7)) AND (fsm_output(3)) AND (NOT (fsm_output(9))) AND (fsm_output(2))
      AND (NOT (fsm_output(10)));
  mux_1851_nl <= MUX_s_1_2_2(nor_959_nl, and_578_nl, fsm_output(1));
  mux_1852_nl <= MUX_s_1_2_2(nor_958_nl, mux_1851_nl, fsm_output(0));
  mux_1859_nl <= MUX_s_1_2_2(mux_1858_nl, mux_1852_nl, fsm_output(6));
  nor_960_nl <= NOT((NOT (fsm_output(1))) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(3)) OR (NOT (fsm_output(9)))
      OR (fsm_output(2)) OR (fsm_output(10)));
  nor_961_nl <= NOT((fsm_output(1)) OR (fsm_output(5)) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1011")) OR (NOT (fsm_output(7))) OR (fsm_output(3))
      OR (fsm_output(9)) OR not_tmp_253);
  mux_1849_nl <= MUX_s_1_2_2(nor_960_nl, nor_961_nl, fsm_output(0));
  nor_962_nl <= NOT((NOT((fsm_output(5)) AND (fsm_output(7)) AND CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)=STD_LOGIC_VECTOR'("1011")) AND (fsm_output(3)) AND (NOT (fsm_output(9)))))
      OR not_tmp_253);
  nor_963_nl <= NOT((NOT (fsm_output(7))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1011")) OR (fsm_output(3)) OR (NOT (fsm_output(9)))
      OR (fsm_output(2)) OR (fsm_output(10)));
  nor_964_nl <= NOT((NOT((fsm_output(7)) AND CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1011"))
      AND (fsm_output(3)) AND (NOT (fsm_output(9))))) OR not_tmp_253);
  mux_1845_nl <= MUX_s_1_2_2(nor_963_nl, nor_964_nl, fsm_output(5));
  mux_1846_nl <= MUX_s_1_2_2(nor_962_nl, mux_1845_nl, COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm);
  nor_965_nl <= NOT((NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1011")) OR (fsm_output(3)) OR (fsm_output(9))
      OR (NOT (fsm_output(2))) OR (fsm_output(10)));
  mux_1847_nl <= MUX_s_1_2_2(mux_1846_nl, nor_965_nl, fsm_output(1));
  and_579_nl <= CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1011")) AND
      (fsm_output(5)) AND (fsm_output(7)) AND (fsm_output(3)) AND (fsm_output(9))
      AND (NOT (fsm_output(2))) AND (NOT (fsm_output(10)));
  nor_966_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(3)) OR (fsm_output(9))
      OR (fsm_output(2)) OR (NOT (fsm_output(10))));
  mux_1844_nl <= MUX_s_1_2_2(and_579_nl, nor_966_nl, fsm_output(1));
  mux_1848_nl <= MUX_s_1_2_2(mux_1847_nl, mux_1844_nl, fsm_output(0));
  mux_1850_nl <= MUX_s_1_2_2(mux_1849_nl, mux_1848_nl, fsm_output(6));
  mux_1860_nl <= MUX_s_1_2_2(mux_1859_nl, mux_1850_nl, fsm_output(8));
  vec_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_1875_nl, mux_1860_nl,
      fsm_output(4));
  or_1944_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR
      (NOT (fsm_output(9))) OR (NOT (fsm_output(5))) OR (fsm_output(10));
  or_1943_nl <= (NOT (fsm_output(9))) OR (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR not_tmp_357;
  mux_1902_nl <= MUX_s_1_2_2(or_1944_nl, or_1943_nl, fsm_output(7));
  or_1941_nl <= CONV_SL_1_1(VEC_LOOP_j_sva_11_0(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("11"))
      OR (NOT (fsm_output(7))) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (fsm_output(9)) OR (fsm_output(5)) OR (fsm_output(10));
  mux_1903_nl <= MUX_s_1_2_2(mux_1902_nl, or_1941_nl, fsm_output(2));
  nor_923_nl <= NOT((fsm_output(6)) OR (fsm_output(4)) OR mux_1903_nl);
  nor_924_nl <= NOT((fsm_output(6)) OR (fsm_output(4)) OR (NOT (fsm_output(2))) OR
      (fsm_output(7)) OR (fsm_output(9)) OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR not_tmp_357);
  mux_1904_nl <= MUX_s_1_2_2(nor_923_nl, nor_924_nl, fsm_output(8));
  nor_925_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT (fsm_output(6))) OR (NOT (fsm_output(4))) OR (fsm_output(2)) OR (NOT
      (fsm_output(7))) OR (fsm_output(9)) OR not_tmp_248);
  nor_926_nl <= NOT((fsm_output(4)) OR (fsm_output(2)) OR (fsm_output(7)) OR (NOT
      (fsm_output(9))) OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1100")) OR (fsm_output(10)));
  nor_927_nl <= NOT((NOT (fsm_output(2))) OR (fsm_output(7)) OR (fsm_output(9)) OR
      (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("1100")) OR (fsm_output(10)));
  nor_928_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT (fsm_output(2))) OR (fsm_output(7)) OR (NOT (fsm_output(9))) OR (fsm_output(5))
      OR (fsm_output(10)));
  mux_1899_nl <= MUX_s_1_2_2(nor_927_nl, nor_928_nl, fsm_output(4));
  mux_1900_nl <= MUX_s_1_2_2(nor_926_nl, mux_1899_nl, fsm_output(6));
  mux_1901_nl <= MUX_s_1_2_2(nor_925_nl, mux_1900_nl, fsm_output(8));
  mux_1905_nl <= MUX_s_1_2_2(mux_1904_nl, mux_1901_nl, fsm_output(0));
  nand_261_nl <= NOT((COMP_LOOP_acc_16_psp_sva(0)) AND (fsm_output(4)) AND (fsm_output(2))
      AND (VEC_LOOP_j_sva_11_0(2)) AND (fsm_output(7)) AND CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1
      DOWNTO 0)=STD_LOGIC_VECTOR'("00")) AND (fsm_output(9)) AND (fsm_output(5))
      AND (NOT (fsm_output(10))));
  or_1931_nl <= CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR (fsm_output(2)) OR (fsm_output(7)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR (fsm_output(9)) OR (fsm_output(5)) OR
      (NOT (fsm_output(10)));
  mux_1896_nl <= MUX_s_1_2_2(mux_tmp_1884, or_1931_nl, fsm_output(4));
  mux_1897_nl <= MUX_s_1_2_2(nand_261_nl, mux_1896_nl, fsm_output(6));
  and_574_nl <= (fsm_output(8)) AND (NOT mux_1897_nl);
  or_1928_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(7))) OR (NOT (fsm_output(9)))
      OR (fsm_output(5)) OR (NOT (fsm_output(10)));
  or_1926_nl <= (fsm_output(7)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(5)))
      OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR not_tmp_357;
  mux_1893_nl <= MUX_s_1_2_2(or_1926_nl, or_tmp_1858, fsm_output(2));
  mux_1894_nl <= MUX_s_1_2_2(or_1928_nl, mux_1893_nl, fsm_output(4));
  nor_929_nl <= NOT((fsm_output(6)) OR mux_1894_nl);
  nor_930_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(6)) OR (NOT (fsm_output(4))) OR (fsm_output(2)) OR (NOT (fsm_output(7)))
      OR (fsm_output(9)) OR (NOT (fsm_output(5))) OR (fsm_output(10)));
  mux_1895_nl <= MUX_s_1_2_2(nor_929_nl, nor_930_nl, fsm_output(8));
  mux_1898_nl <= MUX_s_1_2_2(and_574_nl, mux_1895_nl, fsm_output(0));
  mux_1906_nl <= MUX_s_1_2_2(mux_1905_nl, mux_1898_nl, fsm_output(3));
  or_1922_nl <= CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (NOT (fsm_output(2))) OR (fsm_output(7)) OR (VEC_LOOP_j_sva_11_0(0)) OR
      nand_337_cse;
  or_1920_nl <= (NOT (fsm_output(2))) OR (fsm_output(7)) OR (fsm_output(9)) OR (NOT
      (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR not_tmp_357;
  mux_1889_nl <= MUX_s_1_2_2(or_1922_nl, or_1920_nl, fsm_output(4));
  nor_931_nl <= NOT((fsm_output(6)) OR mux_1889_nl);
  or_1916_nl <= (fsm_output(9)) OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR not_tmp_357;
  mux_1887_nl <= MUX_s_1_2_2(or_591_cse, or_1916_nl, fsm_output(7));
  mux_1888_nl <= MUX_s_1_2_2(mux_1887_nl, or_tmp_1858, or_1912_cse);
  nor_932_nl <= NOT((NOT (fsm_output(6))) OR (NOT (fsm_output(4))) OR (fsm_output(2))
      OR mux_1888_nl);
  mux_1890_nl <= MUX_s_1_2_2(nor_931_nl, nor_932_nl, fsm_output(8));
  or_1909_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(7)) OR (fsm_output(9)) OR not_tmp_248;
  or_1907_nl <= (NOT (fsm_output(7))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1100")) OR (NOT (fsm_output(9))) OR (fsm_output(5))
      OR (fsm_output(10));
  mux_1885_nl <= MUX_s_1_2_2(or_1909_nl, or_1907_nl, fsm_output(2));
  mux_1886_nl <= MUX_s_1_2_2(mux_1885_nl, mux_tmp_1884, fsm_output(4));
  nor_933_nl <= NOT((fsm_output(8)) OR (fsm_output(6)) OR mux_1886_nl);
  mux_1891_nl <= MUX_s_1_2_2(mux_1890_nl, nor_933_nl, fsm_output(0));
  or_1902_nl <= CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (fsm_output(2)) OR (NOT (fsm_output(7))) OR (VEC_LOOP_j_sva_11_0(0)) OR
      (fsm_output(9)) OR (fsm_output(5)) OR (NOT (fsm_output(10)));
  or_1900_nl <= (fsm_output(2)) OR (NOT (fsm_output(7))) OR (NOT (fsm_output(9)))
      OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("1100")) OR (fsm_output(10));
  mux_1881_nl <= MUX_s_1_2_2(or_1902_nl, or_1900_nl, fsm_output(4));
  or_1899_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(7))) OR (VEC_LOOP_j_sva_11_0(0))
      OR (NOT (fsm_output(9))) OR (NOT (fsm_output(5))) OR (fsm_output(10));
  or_1898_nl <= (NOT (fsm_output(2))) OR (NOT (fsm_output(7))) OR (fsm_output(9))
      OR (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("1100")) OR (fsm_output(10));
  mux_1880_nl <= MUX_s_1_2_2(or_1899_nl, or_1898_nl, fsm_output(4));
  mux_1882_nl <= MUX_s_1_2_2(mux_1881_nl, mux_1880_nl, fsm_output(6));
  nor_934_nl <= NOT((fsm_output(8)) OR mux_1882_nl);
  nor_935_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT (fsm_output(6))) OR (fsm_output(4)) OR (fsm_output(2)) OR (NOT (fsm_output(7)))
      OR (fsm_output(9)) OR (NOT (fsm_output(5))) OR (fsm_output(10)));
  nor_936_nl <= NOT((NOT (fsm_output(4))) OR (NOT (fsm_output(2))) OR (NOT (fsm_output(7)))
      OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(9)) OR not_tmp_248);
  or_1893_nl <= (fsm_output(7)) OR (fsm_output(9)) OR (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR not_tmp_357;
  or_1891_nl <= (NOT (fsm_output(7))) OR (NOT (fsm_output(9))) OR (fsm_output(5))
      OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(10));
  mux_1877_nl <= MUX_s_1_2_2(or_1893_nl, or_1891_nl, fsm_output(2));
  nor_937_nl <= NOT((fsm_output(4)) OR mux_1877_nl);
  mux_1878_nl <= MUX_s_1_2_2(nor_936_nl, nor_937_nl, fsm_output(6));
  mux_1879_nl <= MUX_s_1_2_2(nor_935_nl, mux_1878_nl, fsm_output(8));
  mux_1883_nl <= MUX_s_1_2_2(nor_934_nl, mux_1879_nl, fsm_output(0));
  mux_1892_nl <= MUX_s_1_2_2(mux_1891_nl, mux_1883_nl, fsm_output(3));
  vec_rsc_0_12_i_wea_d_pff <= MUX_s_1_2_2(mux_1906_nl, mux_1892_nl, fsm_output(1));
  or_2000_nl <= (NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(2))) OR (fsm_output(10));
  or_1999_nl <= (fsm_output(7)) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(2)) OR (NOT (fsm_output(10)));
  mux_1937_nl <= MUX_s_1_2_2(or_2000_nl, or_1999_nl, fsm_output(5));
  nor_892_nl <= NOT((fsm_output(1)) OR mux_1937_nl);
  nor_893_nl <= NOT((fsm_output(5)) OR (NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1100")) OR (fsm_output(3)) OR (fsm_output(9))
      OR (fsm_output(2)) OR (fsm_output(10)));
  nor_894_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT (fsm_output(7))) OR (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_253);
  nor_895_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(7)) OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (fsm_output(2))
      OR (NOT (fsm_output(10))));
  mux_1935_nl <= MUX_s_1_2_2(nor_894_nl, nor_895_nl, fsm_output(5));
  mux_1936_nl <= MUX_s_1_2_2(nor_893_nl, mux_1935_nl, fsm_output(1));
  mux_1938_nl <= MUX_s_1_2_2(nor_892_nl, mux_1936_nl, fsm_output(0));
  and_571_nl <= (fsm_output(6)) AND mux_1938_nl;
  nor_896_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR (fsm_output(2)) OR (fsm_output(10)));
  nor_898_nl <= NOT((fsm_output(7)) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR not_tmp_253);
  mux_1930_nl <= MUX_s_1_2_2(nor_1445_cse, nor_898_nl, fsm_output(5));
  nor_899_nl <= NOT((NOT (fsm_output(5))) OR (fsm_output(7)) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1100")) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR not_tmp_253);
  or_1986_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm);
  mux_1931_nl <= MUX_s_1_2_2(mux_1930_nl, nor_899_nl, or_1986_nl);
  mux_1932_nl <= MUX_s_1_2_2(nor_896_nl, mux_1931_nl, fsm_output(1));
  nor_900_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR
      (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_253);
  nor_901_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (NOT
      (fsm_output(2))) OR (fsm_output(10)));
  nor_902_nl <= NOT((fsm_output(7)) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9))) OR (fsm_output(2)) OR (fsm_output(10)));
  mux_1928_nl <= MUX_s_1_2_2(nor_901_nl, nor_902_nl, fsm_output(5));
  mux_1929_nl <= MUX_s_1_2_2(nor_900_nl, mux_1928_nl, fsm_output(1));
  mux_1933_nl <= MUX_s_1_2_2(mux_1932_nl, mux_1929_nl, fsm_output(0));
  nor_903_nl <= NOT((NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (NOT (fsm_output(5)))
      OR (fsm_output(7)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR not_tmp_253);
  nor_904_nl <= NOT((NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (NOT (fsm_output(5)))
      OR (fsm_output(7)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(3)) OR (fsm_output(9)) OR (NOT (fsm_output(2))) OR (fsm_output(10)));
  mux_1926_nl <= MUX_s_1_2_2(nor_903_nl, nor_904_nl, fsm_output(1));
  nor_905_nl <= NOT((fsm_output(1)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR mux_1925_cse);
  mux_1927_nl <= MUX_s_1_2_2(mux_1926_nl, nor_905_nl, fsm_output(0));
  mux_1934_nl <= MUX_s_1_2_2(mux_1933_nl, mux_1927_nl, fsm_output(6));
  mux_1939_nl <= MUX_s_1_2_2(and_571_nl, mux_1934_nl, fsm_output(8));
  nor_906_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (fsm_output(2))
      OR (fsm_output(10)));
  nor_907_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(7)) OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(2)))
      OR (fsm_output(10)));
  mux_1920_nl <= MUX_s_1_2_2(nor_906_nl, nor_907_nl, fsm_output(5));
  and_572_nl <= COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm AND mux_1920_nl;
  nor_908_nl <= NOT((NOT (fsm_output(7))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1100")) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR not_tmp_253);
  nor_909_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(7)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9))) OR (fsm_output(2))
      OR (NOT (fsm_output(10))));
  mux_1919_nl <= MUX_s_1_2_2(nor_908_nl, nor_909_nl, fsm_output(5));
  and_573_nl <= COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm AND mux_1919_nl;
  mux_1921_nl <= MUX_s_1_2_2(and_572_nl, and_573_nl, fsm_output(1));
  nor_910_nl <= NOT((NOT (VEC_LOOP_j_sva_11_0(3))) OR (VEC_LOOP_j_sva_11_0(1)) OR
      (VEC_LOOP_j_sva_11_0(0)) OR (NOT (fsm_output(5))) OR (NOT (VEC_LOOP_j_sva_11_0(2)))
      OR (fsm_output(7)) OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(2))
      OR (fsm_output(10)));
  nor_911_nl <= NOT((VEC_LOOP_j_sva_11_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR mux_1917_cse);
  mux_1918_nl <= MUX_s_1_2_2(nor_910_nl, nor_911_nl, fsm_output(1));
  mux_1922_nl <= MUX_s_1_2_2(mux_1921_nl, mux_1918_nl, fsm_output(0));
  nor_912_nl <= NOT((NOT (fsm_output(1))) OR (fsm_output(5)) OR (fsm_output(7)) OR
      CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100")) OR (NOT (fsm_output(3)))
      OR (fsm_output(9)) OR (fsm_output(2)) OR (fsm_output(10)));
  nor_913_nl <= NOT((fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(3))) OR
      CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100")) OR (NOT (fsm_output(9)))
      OR (NOT (fsm_output(2))) OR (fsm_output(10)));
  nor_914_nl <= NOT((VEC_LOOP_j_sva_11_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (NOT
      (fsm_output(2))) OR (fsm_output(10)));
  mux_1915_nl <= MUX_s_1_2_2(nor_913_nl, nor_914_nl, fsm_output(1));
  mux_1916_nl <= MUX_s_1_2_2(nor_912_nl, mux_1915_nl, fsm_output(0));
  mux_1923_nl <= MUX_s_1_2_2(mux_1922_nl, mux_1916_nl, fsm_output(6));
  nor_915_nl <= NOT((NOT (fsm_output(1))) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(3)) OR (NOT (fsm_output(9)))
      OR (fsm_output(2)) OR (fsm_output(10)));
  nor_916_nl <= NOT((fsm_output(1)) OR (fsm_output(5)) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1100")) OR (NOT (fsm_output(7))) OR (fsm_output(3))
      OR (fsm_output(9)) OR not_tmp_253);
  mux_1913_nl <= MUX_s_1_2_2(nor_915_nl, nor_916_nl, fsm_output(0));
  nor_917_nl <= NOT((NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1100")) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR not_tmp_253);
  nor_918_nl <= NOT((NOT (fsm_output(7))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1100")) OR (fsm_output(3)) OR (NOT (fsm_output(9)))
      OR (fsm_output(2)) OR (fsm_output(10)));
  nor_919_nl <= NOT((NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR not_tmp_253);
  mux_1909_nl <= MUX_s_1_2_2(nor_918_nl, nor_919_nl, fsm_output(5));
  mux_1910_nl <= MUX_s_1_2_2(nor_917_nl, mux_1909_nl, COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm);
  nor_920_nl <= NOT((NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1100")) OR (fsm_output(3)) OR (fsm_output(9))
      OR (NOT (fsm_output(2))) OR (fsm_output(10)));
  mux_1911_nl <= MUX_s_1_2_2(mux_1910_nl, nor_920_nl, fsm_output(1));
  nor_921_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3)))
      OR (NOT (fsm_output(9))) OR (fsm_output(2)) OR (fsm_output(10)));
  nor_922_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (VEC_LOOP_j_sva_11_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR
      (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(3)) OR (fsm_output(9))
      OR (fsm_output(2)) OR (NOT (fsm_output(10))));
  mux_1908_nl <= MUX_s_1_2_2(nor_921_nl, nor_922_nl, fsm_output(1));
  mux_1912_nl <= MUX_s_1_2_2(mux_1911_nl, mux_1908_nl, fsm_output(0));
  mux_1914_nl <= MUX_s_1_2_2(mux_1913_nl, mux_1912_nl, fsm_output(6));
  mux_1924_nl <= MUX_s_1_2_2(mux_1923_nl, mux_1914_nl, fsm_output(8));
  vec_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_1939_nl, mux_1924_nl,
      fsm_output(4));
  nand_250_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)=STD_LOGIC_VECTOR'("01")) AND
      (fsm_output(9)) AND (fsm_output(5)) AND (NOT (fsm_output(10))));
  or_2054_nl <= (NOT((fsm_output(9)) AND (fsm_output(5)) AND CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(1
      DOWNTO 0)=STD_LOGIC_VECTOR'("01")))) OR not_tmp_357;
  mux_1966_nl <= MUX_s_1_2_2(nand_250_nl, or_2054_nl, fsm_output(7));
  or_2052_nl <= CONV_SL_1_1(VEC_LOOP_j_sva_11_0(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("11"))
      OR (NOT (fsm_output(7))) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR (fsm_output(9)) OR (fsm_output(5)) OR (fsm_output(10));
  mux_1967_nl <= MUX_s_1_2_2(mux_1966_nl, or_2052_nl, fsm_output(2));
  nor_877_nl <= NOT((fsm_output(6)) OR (fsm_output(4)) OR mux_1967_nl);
  nor_878_nl <= NOT((fsm_output(6)) OR (fsm_output(4)) OR (NOT (fsm_output(2))) OR
      (fsm_output(7)) OR (fsm_output(9)) OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR not_tmp_357);
  mux_1968_nl <= MUX_s_1_2_2(nor_877_nl, nor_878_nl, fsm_output(8));
  nor_879_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (NOT (fsm_output(6))) OR (NOT (fsm_output(4))) OR (fsm_output(2)) OR (NOT
      (fsm_output(7))) OR (fsm_output(9)) OR not_tmp_248);
  nor_880_nl <= NOT((fsm_output(4)) OR (fsm_output(2)) OR (fsm_output(7)) OR (NOT
      (fsm_output(9))) OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1101")) OR (fsm_output(10)));
  nor_881_nl <= NOT((NOT (fsm_output(2))) OR (fsm_output(7)) OR (fsm_output(9)) OR
      (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("1101")) OR (fsm_output(10)));
  nor_882_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (NOT (fsm_output(2))) OR (fsm_output(7)) OR (NOT (fsm_output(9))) OR (fsm_output(5))
      OR (fsm_output(10)));
  mux_1963_nl <= MUX_s_1_2_2(nor_881_nl, nor_882_nl, fsm_output(4));
  mux_1964_nl <= MUX_s_1_2_2(nor_880_nl, mux_1963_nl, fsm_output(6));
  mux_1965_nl <= MUX_s_1_2_2(nor_879_nl, mux_1964_nl, fsm_output(8));
  mux_1969_nl <= MUX_s_1_2_2(mux_1968_nl, mux_1965_nl, fsm_output(0));
  nand_252_nl <= NOT((COMP_LOOP_acc_16_psp_sva(0)) AND (fsm_output(4)) AND (fsm_output(2))
      AND (VEC_LOOP_j_sva_11_0(2)) AND (fsm_output(7)) AND CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1
      DOWNTO 0)=STD_LOGIC_VECTOR'("01")) AND (fsm_output(9)) AND (fsm_output(5))
      AND (NOT (fsm_output(10))));
  or_2042_nl <= CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR (fsm_output(2)) OR (fsm_output(7)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR (fsm_output(9)) OR (fsm_output(5)) OR
      (NOT (fsm_output(10)));
  mux_1960_nl <= MUX_s_1_2_2(mux_tmp_1948, or_2042_nl, fsm_output(4));
  mux_1961_nl <= MUX_s_1_2_2(nand_252_nl, mux_1960_nl, fsm_output(6));
  and_570_nl <= (fsm_output(8)) AND (NOT mux_1961_nl);
  nand_397_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1101"))
      AND (fsm_output(2)) AND (fsm_output(7)) AND (fsm_output(9)) AND (NOT (fsm_output(5)))
      AND (fsm_output(10)));
  or_2037_nl <= (fsm_output(7)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(5)))
      OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR not_tmp_357;
  mux_1957_nl <= MUX_s_1_2_2(or_2037_nl, or_tmp_1969, fsm_output(2));
  mux_1958_nl <= MUX_s_1_2_2(nand_397_nl, mux_1957_nl, fsm_output(4));
  nor_883_nl <= NOT((fsm_output(6)) OR mux_1958_nl);
  nor_884_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(6)) OR (NOT (fsm_output(4))) OR (fsm_output(2)) OR (NOT (fsm_output(7)))
      OR (fsm_output(9)) OR (NOT (fsm_output(5))) OR (fsm_output(10)));
  mux_1959_nl <= MUX_s_1_2_2(nor_883_nl, nor_884_nl, fsm_output(8));
  mux_1962_nl <= MUX_s_1_2_2(and_570_nl, mux_1959_nl, fsm_output(0));
  mux_1970_nl <= MUX_s_1_2_2(mux_1969_nl, mux_1962_nl, fsm_output(3));
  or_2033_nl <= CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (NOT (fsm_output(2))) OR (fsm_output(7)) OR nand_334_cse;
  or_2031_nl <= (NOT (fsm_output(2))) OR (fsm_output(7)) OR (fsm_output(9)) OR (NOT
      (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR not_tmp_357;
  mux_1953_nl <= MUX_s_1_2_2(or_2033_nl, or_2031_nl, fsm_output(4));
  nor_885_nl <= NOT((fsm_output(6)) OR mux_1953_nl);
  or_2027_nl <= (fsm_output(9)) OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR not_tmp_357;
  mux_1951_nl <= MUX_s_1_2_2(or_702_cse, or_2027_nl, fsm_output(7));
  mux_1952_nl <= MUX_s_1_2_2(mux_1951_nl, or_tmp_1969, or_1912_cse);
  nor_886_nl <= NOT((NOT (fsm_output(6))) OR (NOT (fsm_output(4))) OR (fsm_output(2))
      OR mux_1952_nl);
  mux_1954_nl <= MUX_s_1_2_2(nor_885_nl, nor_886_nl, fsm_output(8));
  or_2020_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(7)) OR (fsm_output(9)) OR not_tmp_248;
  or_2018_nl <= (NOT (fsm_output(7))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1101")) OR (NOT (fsm_output(9))) OR (fsm_output(5))
      OR (fsm_output(10));
  mux_1949_nl <= MUX_s_1_2_2(or_2020_nl, or_2018_nl, fsm_output(2));
  mux_1950_nl <= MUX_s_1_2_2(mux_1949_nl, mux_tmp_1948, fsm_output(4));
  nor_887_nl <= NOT((fsm_output(8)) OR (fsm_output(6)) OR mux_1950_nl);
  mux_1955_nl <= MUX_s_1_2_2(mux_1954_nl, nor_887_nl, fsm_output(0));
  or_2013_nl <= CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (fsm_output(2)) OR (NOT (fsm_output(7))) OR (NOT (VEC_LOOP_j_sva_11_0(0)))
      OR (fsm_output(9)) OR (fsm_output(5)) OR (NOT (fsm_output(10)));
  or_2011_nl <= (fsm_output(2)) OR (NOT (fsm_output(7))) OR (NOT (fsm_output(9)))
      OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("1101")) OR (fsm_output(10));
  mux_1945_nl <= MUX_s_1_2_2(or_2013_nl, or_2011_nl, fsm_output(4));
  nand_255_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("110"))
      AND (fsm_output(2)) AND (fsm_output(7)) AND (VEC_LOOP_j_sva_11_0(0)) AND (fsm_output(9))
      AND (fsm_output(5)) AND (NOT (fsm_output(10))));
  or_2009_nl <= (NOT (fsm_output(2))) OR (NOT (fsm_output(7))) OR (fsm_output(9))
      OR (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("1101")) OR (fsm_output(10));
  mux_1944_nl <= MUX_s_1_2_2(nand_255_nl, or_2009_nl, fsm_output(4));
  mux_1946_nl <= MUX_s_1_2_2(mux_1945_nl, mux_1944_nl, fsm_output(6));
  nor_888_nl <= NOT((fsm_output(8)) OR mux_1946_nl);
  nor_889_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (NOT (fsm_output(6))) OR (fsm_output(4)) OR (fsm_output(2)) OR (NOT (fsm_output(7)))
      OR (fsm_output(9)) OR (NOT (fsm_output(5))) OR (fsm_output(10)));
  nor_890_nl <= NOT((NOT((fsm_output(4)) AND (fsm_output(2)) AND (fsm_output(7))
      AND CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1101"))
      AND (NOT (fsm_output(9))))) OR not_tmp_248);
  or_2004_nl <= (fsm_output(7)) OR (fsm_output(9)) OR (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR not_tmp_357;
  or_2002_nl <= (NOT (fsm_output(7))) OR (NOT (fsm_output(9))) OR (fsm_output(5))
      OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(10));
  mux_1941_nl <= MUX_s_1_2_2(or_2004_nl, or_2002_nl, fsm_output(2));
  nor_891_nl <= NOT((fsm_output(4)) OR mux_1941_nl);
  mux_1942_nl <= MUX_s_1_2_2(nor_890_nl, nor_891_nl, fsm_output(6));
  mux_1943_nl <= MUX_s_1_2_2(nor_889_nl, mux_1942_nl, fsm_output(8));
  mux_1947_nl <= MUX_s_1_2_2(nor_888_nl, mux_1943_nl, fsm_output(0));
  mux_1956_nl <= MUX_s_1_2_2(mux_1955_nl, mux_1947_nl, fsm_output(3));
  vec_rsc_0_13_i_wea_d_pff <= MUX_s_1_2_2(mux_1970_nl, mux_1956_nl, fsm_output(1));
  or_2111_nl <= (NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(2))) OR (fsm_output(10));
  or_2110_nl <= (fsm_output(7)) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(2)) OR (NOT (fsm_output(10)));
  mux_2001_nl <= MUX_s_1_2_2(or_2111_nl, or_2110_nl, fsm_output(5));
  nor_848_nl <= NOT((fsm_output(1)) OR mux_2001_nl);
  nor_849_nl <= NOT((fsm_output(5)) OR (NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1101")) OR (fsm_output(3)) OR (fsm_output(9))
      OR (fsm_output(2)) OR (fsm_output(10)));
  nor_850_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (NOT (fsm_output(7))) OR (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_253);
  nor_851_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(7)) OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (fsm_output(2))
      OR (NOT (fsm_output(10))));
  mux_1999_nl <= MUX_s_1_2_2(nor_850_nl, nor_851_nl, fsm_output(5));
  mux_2000_nl <= MUX_s_1_2_2(nor_849_nl, mux_1999_nl, fsm_output(1));
  mux_2002_nl <= MUX_s_1_2_2(nor_848_nl, mux_2000_nl, fsm_output(0));
  and_565_nl <= (fsm_output(6)) AND mux_2002_nl;
  nor_852_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR (fsm_output(2)) OR (fsm_output(10)));
  nor_854_nl <= NOT((fsm_output(7)) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR not_tmp_253);
  mux_1994_nl <= MUX_s_1_2_2(nor_1445_cse, nor_854_nl, fsm_output(5));
  nor_855_nl <= NOT((NOT (fsm_output(5))) OR (fsm_output(7)) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1101")) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR not_tmp_253);
  nand_243_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1101"))
      AND COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm);
  mux_1995_nl <= MUX_s_1_2_2(mux_1994_nl, nor_855_nl, nand_243_nl);
  mux_1996_nl <= MUX_s_1_2_2(nor_852_nl, mux_1995_nl, fsm_output(1));
  nor_856_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR
      (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_253);
  nor_857_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (NOT
      (fsm_output(2))) OR (fsm_output(10)));
  nor_858_nl <= NOT((fsm_output(7)) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9))) OR (fsm_output(2)) OR (fsm_output(10)));
  mux_1992_nl <= MUX_s_1_2_2(nor_857_nl, nor_858_nl, fsm_output(5));
  mux_1993_nl <= MUX_s_1_2_2(nor_856_nl, mux_1992_nl, fsm_output(1));
  mux_1997_nl <= MUX_s_1_2_2(mux_1996_nl, mux_1993_nl, fsm_output(0));
  nor_859_nl <= NOT((NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (NOT (fsm_output(5)))
      OR (fsm_output(7)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR not_tmp_253);
  nor_860_nl <= NOT((NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (NOT (fsm_output(5)))
      OR (fsm_output(7)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(3)) OR (fsm_output(9)) OR (NOT (fsm_output(2))) OR (fsm_output(10)));
  mux_1990_nl <= MUX_s_1_2_2(nor_859_nl, nor_860_nl, fsm_output(1));
  nor_861_nl <= NOT((fsm_output(1)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR mux_1925_cse);
  mux_1991_nl <= MUX_s_1_2_2(mux_1990_nl, nor_861_nl, fsm_output(0));
  mux_1998_nl <= MUX_s_1_2_2(mux_1997_nl, mux_1991_nl, fsm_output(6));
  mux_2003_nl <= MUX_s_1_2_2(and_565_nl, mux_1998_nl, fsm_output(8));
  nor_862_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (fsm_output(2))
      OR (fsm_output(10)));
  nor_863_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(7)) OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(2)))
      OR (fsm_output(10)));
  mux_1984_nl <= MUX_s_1_2_2(nor_862_nl, nor_863_nl, fsm_output(5));
  and_566_nl <= COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm AND mux_1984_nl;
  nor_864_nl <= NOT((NOT((fsm_output(7)) AND CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3
      DOWNTO 0)=STD_LOGIC_VECTOR'("1101")) AND (fsm_output(3)) AND (NOT (fsm_output(9)))))
      OR not_tmp_253);
  nor_865_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(7)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9))) OR (fsm_output(2))
      OR (NOT (fsm_output(10))));
  mux_1983_nl <= MUX_s_1_2_2(nor_864_nl, nor_865_nl, fsm_output(5));
  and_567_nl <= COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm AND mux_1983_nl;
  mux_1985_nl <= MUX_s_1_2_2(and_566_nl, and_567_nl, fsm_output(1));
  nor_866_nl <= NOT((NOT (VEC_LOOP_j_sva_11_0(3))) OR (VEC_LOOP_j_sva_11_0(1)) OR
      (NOT (VEC_LOOP_j_sva_11_0(0))) OR (NOT (fsm_output(5))) OR (NOT (VEC_LOOP_j_sva_11_0(2)))
      OR (fsm_output(7)) OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(2))
      OR (fsm_output(10)));
  nor_867_nl <= NOT(nand_332_cse OR mux_1917_cse);
  mux_1982_nl <= MUX_s_1_2_2(nor_866_nl, nor_867_nl, fsm_output(1));
  mux_1986_nl <= MUX_s_1_2_2(mux_1985_nl, mux_1982_nl, fsm_output(0));
  nor_868_nl <= NOT((NOT (fsm_output(1))) OR (fsm_output(5)) OR (fsm_output(7)) OR
      CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101")) OR (NOT (fsm_output(3)))
      OR (fsm_output(9)) OR (fsm_output(2)) OR (fsm_output(10)));
  nor_869_nl <= NOT((fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(3))) OR
      CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101")) OR (NOT (fsm_output(9)))
      OR (NOT (fsm_output(2))) OR (fsm_output(10)));
  and_568_nl <= (VEC_LOOP_j_sva_11_0(0)) AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm
      AND (fsm_output(5)) AND CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("110"))
      AND (fsm_output(7)) AND (fsm_output(3)) AND (NOT (fsm_output(9))) AND (fsm_output(2))
      AND (NOT (fsm_output(10)));
  mux_1979_nl <= MUX_s_1_2_2(nor_869_nl, and_568_nl, fsm_output(1));
  mux_1980_nl <= MUX_s_1_2_2(nor_868_nl, mux_1979_nl, fsm_output(0));
  mux_1987_nl <= MUX_s_1_2_2(mux_1986_nl, mux_1980_nl, fsm_output(6));
  nor_870_nl <= NOT((NOT (fsm_output(1))) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(3)) OR (NOT (fsm_output(9)))
      OR (fsm_output(2)) OR (fsm_output(10)));
  nor_871_nl <= NOT((fsm_output(1)) OR (fsm_output(5)) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1101")) OR (NOT (fsm_output(7))) OR (fsm_output(3))
      OR (fsm_output(9)) OR not_tmp_253);
  mux_1977_nl <= MUX_s_1_2_2(nor_870_nl, nor_871_nl, fsm_output(0));
  nor_872_nl <= NOT((NOT((fsm_output(5)) AND (fsm_output(7)) AND CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)=STD_LOGIC_VECTOR'("1101")) AND (fsm_output(3)) AND (NOT (fsm_output(9)))))
      OR not_tmp_253);
  nor_873_nl <= NOT((NOT (fsm_output(7))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1101")) OR (fsm_output(3)) OR (NOT (fsm_output(9)))
      OR (fsm_output(2)) OR (fsm_output(10)));
  nor_874_nl <= NOT((NOT((fsm_output(7)) AND CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1101"))
      AND (fsm_output(3)) AND (NOT (fsm_output(9))))) OR not_tmp_253);
  mux_1973_nl <= MUX_s_1_2_2(nor_873_nl, nor_874_nl, fsm_output(5));
  mux_1974_nl <= MUX_s_1_2_2(nor_872_nl, mux_1973_nl, COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm);
  nor_875_nl <= NOT((NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1101")) OR (fsm_output(3)) OR (fsm_output(9))
      OR (NOT (fsm_output(2))) OR (fsm_output(10)));
  mux_1975_nl <= MUX_s_1_2_2(mux_1974_nl, nor_875_nl, fsm_output(1));
  and_569_nl <= CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1101")) AND
      (fsm_output(5)) AND (fsm_output(7)) AND (fsm_output(3)) AND (fsm_output(9))
      AND (NOT (fsm_output(2))) AND (NOT (fsm_output(10)));
  nor_876_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(3)) OR (fsm_output(9))
      OR (fsm_output(2)) OR (NOT (fsm_output(10))));
  mux_1972_nl <= MUX_s_1_2_2(and_569_nl, nor_876_nl, fsm_output(1));
  mux_1976_nl <= MUX_s_1_2_2(mux_1975_nl, mux_1972_nl, fsm_output(0));
  mux_1978_nl <= MUX_s_1_2_2(mux_1977_nl, mux_1976_nl, fsm_output(6));
  mux_1988_nl <= MUX_s_1_2_2(mux_1987_nl, mux_1978_nl, fsm_output(8));
  vec_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_2003_nl, mux_1988_nl,
      fsm_output(4));
  nand_235_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)=STD_LOGIC_VECTOR'("10")) AND
      (fsm_output(9)) AND (fsm_output(5)) AND (NOT (fsm_output(10))));
  or_2164_nl <= (NOT (fsm_output(9))) OR (NOT (fsm_output(5))) OR (COMP_LOOP_acc_10_cse_12_1_1_sva(0))
      OR not_tmp_377;
  mux_2030_nl <= MUX_s_1_2_2(nand_235_nl, or_2164_nl, fsm_output(7));
  or_2162_nl <= CONV_SL_1_1(VEC_LOOP_j_sva_11_0(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("11"))
      OR (NOT (fsm_output(7))) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (fsm_output(9)) OR (fsm_output(5)) OR (fsm_output(10));
  mux_2031_nl <= MUX_s_1_2_2(mux_2030_nl, or_2162_nl, fsm_output(2));
  nor_833_nl <= NOT((fsm_output(6)) OR (fsm_output(4)) OR mux_2031_nl);
  nor_834_nl <= NOT((fsm_output(6)) OR (fsm_output(4)) OR (NOT (fsm_output(2))) OR
      (fsm_output(7)) OR (fsm_output(9)) OR (fsm_output(5)) OR (COMP_LOOP_acc_10_cse_12_1_1_sva(0))
      OR not_tmp_377);
  mux_2032_nl <= MUX_s_1_2_2(nor_833_nl, nor_834_nl, fsm_output(8));
  nor_835_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (NOT (fsm_output(6))) OR (NOT (fsm_output(4))) OR (fsm_output(2)) OR (NOT
      (fsm_output(7))) OR (fsm_output(9)) OR not_tmp_248);
  nor_836_nl <= NOT((fsm_output(4)) OR (fsm_output(2)) OR (fsm_output(7)) OR (NOT
      (fsm_output(9))) OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1110")) OR (fsm_output(10)));
  nor_837_nl <= NOT((NOT (fsm_output(2))) OR (fsm_output(7)) OR (fsm_output(9)) OR
      (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("1110")) OR (fsm_output(10)));
  nor_838_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (NOT (fsm_output(2))) OR (fsm_output(7)) OR (NOT (fsm_output(9))) OR (fsm_output(5))
      OR (fsm_output(10)));
  mux_2027_nl <= MUX_s_1_2_2(nor_837_nl, nor_838_nl, fsm_output(4));
  mux_2028_nl <= MUX_s_1_2_2(nor_836_nl, mux_2027_nl, fsm_output(6));
  mux_2029_nl <= MUX_s_1_2_2(nor_835_nl, mux_2028_nl, fsm_output(8));
  mux_2033_nl <= MUX_s_1_2_2(mux_2032_nl, mux_2029_nl, fsm_output(0));
  nand_236_nl <= NOT((COMP_LOOP_acc_16_psp_sva(0)) AND (fsm_output(4)) AND (fsm_output(2))
      AND (VEC_LOOP_j_sva_11_0(2)) AND (fsm_output(7)) AND CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1
      DOWNTO 0)=STD_LOGIC_VECTOR'("10")) AND (fsm_output(9)) AND (fsm_output(5))
      AND (NOT (fsm_output(10))));
  or_2152_nl <= CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR (fsm_output(2)) OR (fsm_output(7)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR (fsm_output(9)) OR (fsm_output(5)) OR
      (NOT (fsm_output(10)));
  mux_2024_nl <= MUX_s_1_2_2(mux_tmp_2012, or_2152_nl, fsm_output(4));
  mux_2025_nl <= MUX_s_1_2_2(nand_236_nl, mux_2024_nl, fsm_output(6));
  and_563_nl <= (fsm_output(8)) AND (NOT mux_2025_nl);
  nand_396_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1110"))
      AND (fsm_output(2)) AND (fsm_output(7)) AND (fsm_output(9)) AND (NOT (fsm_output(5)))
      AND (fsm_output(10)));
  or_2147_nl <= (fsm_output(7)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(5)))
      OR (COMP_LOOP_acc_10_cse_12_1_1_sva(0)) OR not_tmp_377;
  mux_2021_nl <= MUX_s_1_2_2(or_2147_nl, or_tmp_2082, fsm_output(2));
  mux_2022_nl <= MUX_s_1_2_2(nand_396_nl, mux_2021_nl, fsm_output(4));
  nor_839_nl <= NOT((fsm_output(6)) OR mux_2022_nl);
  nor_840_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(6)) OR (NOT (fsm_output(4))) OR (fsm_output(2)) OR (NOT (fsm_output(7)))
      OR (fsm_output(9)) OR (NOT (fsm_output(5))) OR (fsm_output(10)));
  mux_2023_nl <= MUX_s_1_2_2(nor_839_nl, nor_840_nl, fsm_output(8));
  mux_2026_nl <= MUX_s_1_2_2(and_563_nl, mux_2023_nl, fsm_output(0));
  mux_2034_nl <= MUX_s_1_2_2(mux_2033_nl, mux_2026_nl, fsm_output(3));
  or_2143_nl <= CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("111"))
      OR (NOT (fsm_output(2))) OR (fsm_output(7)) OR (VEC_LOOP_j_sva_11_0(0)) OR
      nand_337_cse;
  or_2141_nl <= (NOT (fsm_output(2))) OR (fsm_output(7)) OR (fsm_output(9)) OR (NOT
      (fsm_output(5))) OR (COMP_LOOP_acc_10_cse_12_1_1_sva(0)) OR not_tmp_377;
  mux_2017_nl <= MUX_s_1_2_2(or_2143_nl, or_2141_nl, fsm_output(4));
  nor_841_nl <= NOT((fsm_output(6)) OR mux_2017_nl);
  or_2135_nl <= (fsm_output(9)) OR (fsm_output(5)) OR (COMP_LOOP_acc_10_cse_12_1_1_sva(0))
      OR not_tmp_377;
  mux_2015_nl <= MUX_s_1_2_2(or_591_cse, or_2135_nl, fsm_output(7));
  mux_2016_nl <= MUX_s_1_2_2(or_tmp_2082, mux_2015_nl, and_564_cse);
  nor_842_nl <= NOT((NOT (fsm_output(6))) OR (NOT (fsm_output(4))) OR (fsm_output(2))
      OR mux_2016_nl);
  mux_2018_nl <= MUX_s_1_2_2(nor_841_nl, nor_842_nl, fsm_output(8));
  or_2131_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(7)) OR (fsm_output(9)) OR not_tmp_248;
  or_2129_nl <= (NOT (fsm_output(7))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1110")) OR (NOT (fsm_output(9))) OR (fsm_output(5))
      OR (fsm_output(10));
  mux_2013_nl <= MUX_s_1_2_2(or_2131_nl, or_2129_nl, fsm_output(2));
  mux_2014_nl <= MUX_s_1_2_2(mux_2013_nl, mux_tmp_2012, fsm_output(4));
  nor_843_nl <= NOT((fsm_output(8)) OR (fsm_output(6)) OR mux_2014_nl);
  mux_2019_nl <= MUX_s_1_2_2(mux_2018_nl, nor_843_nl, fsm_output(0));
  or_2124_nl <= CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("111"))
      OR (fsm_output(2)) OR (NOT (fsm_output(7))) OR (VEC_LOOP_j_sva_11_0(0)) OR
      (fsm_output(9)) OR (fsm_output(5)) OR (NOT (fsm_output(10)));
  or_2122_nl <= (fsm_output(2)) OR (NOT (fsm_output(7))) OR (NOT (fsm_output(9)))
      OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("1110")) OR (fsm_output(10));
  mux_2009_nl <= MUX_s_1_2_2(or_2124_nl, or_2122_nl, fsm_output(4));
  nand_239_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"))
      AND (fsm_output(2)) AND (fsm_output(7)) AND (NOT (VEC_LOOP_j_sva_11_0(0)))
      AND (fsm_output(9)) AND (fsm_output(5)) AND (NOT (fsm_output(10))));
  or_2120_nl <= (NOT (fsm_output(2))) OR (NOT (fsm_output(7))) OR (fsm_output(9))
      OR (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("1110")) OR (fsm_output(10));
  mux_2008_nl <= MUX_s_1_2_2(nand_239_nl, or_2120_nl, fsm_output(4));
  mux_2010_nl <= MUX_s_1_2_2(mux_2009_nl, mux_2008_nl, fsm_output(6));
  nor_844_nl <= NOT((fsm_output(8)) OR mux_2010_nl);
  nor_845_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (NOT (fsm_output(6))) OR (fsm_output(4)) OR (fsm_output(2)) OR (NOT (fsm_output(7)))
      OR (fsm_output(9)) OR (NOT (fsm_output(5))) OR (fsm_output(10)));
  nor_846_nl <= NOT((NOT((fsm_output(4)) AND (fsm_output(2)) AND (fsm_output(7))
      AND CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1110"))
      AND (NOT (fsm_output(9))))) OR not_tmp_248);
  or_2115_nl <= (fsm_output(7)) OR (fsm_output(9)) OR (NOT (fsm_output(5))) OR (COMP_LOOP_acc_10_cse_12_1_1_sva(0))
      OR not_tmp_377;
  or_2113_nl <= (NOT (fsm_output(7))) OR (NOT (fsm_output(9))) OR (fsm_output(5))
      OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(10));
  mux_2005_nl <= MUX_s_1_2_2(or_2115_nl, or_2113_nl, fsm_output(2));
  nor_847_nl <= NOT((fsm_output(4)) OR mux_2005_nl);
  mux_2006_nl <= MUX_s_1_2_2(nor_846_nl, nor_847_nl, fsm_output(6));
  mux_2007_nl <= MUX_s_1_2_2(nor_845_nl, mux_2006_nl, fsm_output(8));
  mux_2011_nl <= MUX_s_1_2_2(nor_844_nl, mux_2007_nl, fsm_output(0));
  mux_2020_nl <= MUX_s_1_2_2(mux_2019_nl, mux_2011_nl, fsm_output(3));
  vec_rsc_0_14_i_wea_d_pff <= MUX_s_1_2_2(mux_2034_nl, mux_2020_nl, fsm_output(1));
  or_2221_nl <= (NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(2))) OR (fsm_output(10));
  or_2220_nl <= (fsm_output(7)) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(2)) OR (NOT (fsm_output(10)));
  mux_2065_nl <= MUX_s_1_2_2(or_2221_nl, or_2220_nl, fsm_output(5));
  nor_804_nl <= NOT((fsm_output(1)) OR mux_2065_nl);
  nor_805_nl <= NOT((fsm_output(5)) OR (NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1110")) OR (fsm_output(3)) OR (fsm_output(9))
      OR (fsm_output(2)) OR (fsm_output(10)));
  nor_806_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (NOT (fsm_output(7))) OR (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_253);
  nor_807_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(7)) OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (fsm_output(2))
      OR (NOT (fsm_output(10))));
  mux_2063_nl <= MUX_s_1_2_2(nor_806_nl, nor_807_nl, fsm_output(5));
  mux_2064_nl <= MUX_s_1_2_2(nor_805_nl, mux_2063_nl, fsm_output(1));
  mux_2066_nl <= MUX_s_1_2_2(nor_804_nl, mux_2064_nl, fsm_output(0));
  and_558_nl <= (fsm_output(6)) AND mux_2066_nl;
  nor_808_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR (fsm_output(2)) OR (fsm_output(10)));
  nor_810_nl <= NOT((fsm_output(7)) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR not_tmp_253);
  mux_2058_nl <= MUX_s_1_2_2(nor_1445_cse, nor_810_nl, fsm_output(5));
  nor_811_nl <= NOT((NOT (fsm_output(5))) OR (fsm_output(7)) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1110")) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR not_tmp_253);
  nand_228_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1110"))
      AND COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm);
  mux_2059_nl <= MUX_s_1_2_2(mux_2058_nl, nor_811_nl, nand_228_nl);
  mux_2060_nl <= MUX_s_1_2_2(nor_808_nl, mux_2059_nl, fsm_output(1));
  nor_812_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR
      (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_253);
  nor_813_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (NOT
      (fsm_output(2))) OR (fsm_output(10)));
  nor_814_nl <= NOT((fsm_output(7)) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9))) OR (fsm_output(2)) OR (fsm_output(10)));
  mux_2056_nl <= MUX_s_1_2_2(nor_813_nl, nor_814_nl, fsm_output(5));
  mux_2057_nl <= MUX_s_1_2_2(nor_812_nl, mux_2056_nl, fsm_output(1));
  mux_2061_nl <= MUX_s_1_2_2(mux_2060_nl, mux_2057_nl, fsm_output(0));
  nor_815_nl <= NOT((NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (NOT (fsm_output(5)))
      OR (fsm_output(7)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR not_tmp_253);
  nor_816_nl <= NOT((NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (NOT (fsm_output(5)))
      OR (fsm_output(7)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(3)) OR (fsm_output(9)) OR (NOT (fsm_output(2))) OR (fsm_output(10)));
  mux_2054_nl <= MUX_s_1_2_2(nor_815_nl, nor_816_nl, fsm_output(1));
  nor_817_nl <= NOT((fsm_output(1)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR mux_1925_cse);
  mux_2055_nl <= MUX_s_1_2_2(mux_2054_nl, nor_817_nl, fsm_output(0));
  mux_2062_nl <= MUX_s_1_2_2(mux_2061_nl, mux_2055_nl, fsm_output(6));
  mux_2067_nl <= MUX_s_1_2_2(and_558_nl, mux_2062_nl, fsm_output(8));
  nor_818_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (fsm_output(2))
      OR (fsm_output(10)));
  nor_819_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(7)) OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(2)))
      OR (fsm_output(10)));
  mux_2048_nl <= MUX_s_1_2_2(nor_818_nl, nor_819_nl, fsm_output(5));
  and_559_nl <= COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm AND mux_2048_nl;
  nor_820_nl <= NOT((NOT((fsm_output(7)) AND CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3
      DOWNTO 0)=STD_LOGIC_VECTOR'("1110")) AND (fsm_output(3)) AND (NOT (fsm_output(9)))))
      OR not_tmp_253);
  nor_821_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(7)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9))) OR (fsm_output(2))
      OR (NOT (fsm_output(10))));
  mux_2047_nl <= MUX_s_1_2_2(nor_820_nl, nor_821_nl, fsm_output(5));
  and_560_nl <= COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm AND mux_2047_nl;
  mux_2049_nl <= MUX_s_1_2_2(and_559_nl, and_560_nl, fsm_output(1));
  nor_822_nl <= NOT((NOT (VEC_LOOP_j_sva_11_0(3))) OR (NOT (VEC_LOOP_j_sva_11_0(1)))
      OR (VEC_LOOP_j_sva_11_0(0)) OR (NOT (fsm_output(5))) OR (NOT (VEC_LOOP_j_sva_11_0(2)))
      OR (fsm_output(7)) OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(2))
      OR (fsm_output(10)));
  nor_823_nl <= NOT((VEC_LOOP_j_sva_11_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR mux_2045_cse);
  mux_2046_nl <= MUX_s_1_2_2(nor_822_nl, nor_823_nl, fsm_output(1));
  mux_2050_nl <= MUX_s_1_2_2(mux_2049_nl, mux_2046_nl, fsm_output(0));
  nor_824_nl <= NOT((NOT (fsm_output(1))) OR (fsm_output(5)) OR (fsm_output(7)) OR
      CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110")) OR (NOT (fsm_output(3)))
      OR (fsm_output(9)) OR (fsm_output(2)) OR (fsm_output(10)));
  nor_825_nl <= NOT((fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(3))) OR
      CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110")) OR (NOT (fsm_output(9)))
      OR (NOT (fsm_output(2))) OR (fsm_output(10)));
  and_561_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"))
      AND (NOT (VEC_LOOP_j_sva_11_0(0))) AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm
      AND (fsm_output(5)) AND (fsm_output(7)) AND (fsm_output(3)) AND (NOT (fsm_output(9)))
      AND (fsm_output(2)) AND (NOT (fsm_output(10)));
  mux_2043_nl <= MUX_s_1_2_2(nor_825_nl, and_561_nl, fsm_output(1));
  mux_2044_nl <= MUX_s_1_2_2(nor_824_nl, mux_2043_nl, fsm_output(0));
  mux_2051_nl <= MUX_s_1_2_2(mux_2050_nl, mux_2044_nl, fsm_output(6));
  nor_826_nl <= NOT((NOT (fsm_output(1))) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(3)) OR (NOT (fsm_output(9)))
      OR (fsm_output(2)) OR (fsm_output(10)));
  nor_827_nl <= NOT((fsm_output(1)) OR (fsm_output(5)) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1110")) OR (NOT (fsm_output(7))) OR (fsm_output(3))
      OR (fsm_output(9)) OR not_tmp_253);
  mux_2041_nl <= MUX_s_1_2_2(nor_826_nl, nor_827_nl, fsm_output(0));
  nor_828_nl <= NOT((NOT((fsm_output(5)) AND (fsm_output(7)) AND CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)=STD_LOGIC_VECTOR'("1110")) AND (fsm_output(3)) AND (NOT (fsm_output(9)))))
      OR not_tmp_253);
  nor_829_nl <= NOT((NOT (fsm_output(7))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1110")) OR (fsm_output(3)) OR (NOT (fsm_output(9)))
      OR (fsm_output(2)) OR (fsm_output(10)));
  nor_830_nl <= NOT((NOT((fsm_output(7)) AND CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1110"))
      AND (fsm_output(3)) AND (NOT (fsm_output(9))))) OR not_tmp_253);
  mux_2037_nl <= MUX_s_1_2_2(nor_829_nl, nor_830_nl, fsm_output(5));
  mux_2038_nl <= MUX_s_1_2_2(nor_828_nl, mux_2037_nl, COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm);
  nor_831_nl <= NOT((NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1110")) OR (fsm_output(3)) OR (fsm_output(9))
      OR (NOT (fsm_output(2))) OR (fsm_output(10)));
  mux_2039_nl <= MUX_s_1_2_2(mux_2038_nl, nor_831_nl, fsm_output(1));
  and_562_nl <= CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1110")) AND
      (fsm_output(5)) AND (fsm_output(7)) AND (fsm_output(3)) AND (fsm_output(9))
      AND (NOT (fsm_output(2))) AND (NOT (fsm_output(10)));
  nor_832_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("111"))
      OR (VEC_LOOP_j_sva_11_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR
      (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(3)) OR (fsm_output(9))
      OR (fsm_output(2)) OR (NOT (fsm_output(10))));
  mux_2036_nl <= MUX_s_1_2_2(and_562_nl, nor_832_nl, fsm_output(1));
  mux_2040_nl <= MUX_s_1_2_2(mux_2039_nl, mux_2036_nl, fsm_output(0));
  mux_2042_nl <= MUX_s_1_2_2(mux_2041_nl, mux_2040_nl, fsm_output(6));
  mux_2052_nl <= MUX_s_1_2_2(mux_2051_nl, mux_2042_nl, fsm_output(8));
  vec_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_2067_nl, mux_2052_nl,
      fsm_output(4));
  and_554_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND
      (fsm_output(9)) AND (fsm_output(5)) AND (NOT (fsm_output(10)));
  mux_2094_nl <= MUX_s_1_2_2(and_554_nl, nor_tmp_265, fsm_output(7));
  or_2271_nl <= CONV_SL_1_1(VEC_LOOP_j_sva_11_0(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("11"))
      OR (NOT (fsm_output(7))) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR (fsm_output(9)) OR (fsm_output(5)) OR (fsm_output(10));
  mux_2095_nl <= MUX_s_1_2_2((NOT mux_2094_nl), or_2271_nl, fsm_output(2));
  nor_789_nl <= NOT((fsm_output(6)) OR (fsm_output(4)) OR mux_2095_nl);
  nor_790_nl <= NOT((fsm_output(6)) OR (fsm_output(4)) OR (NOT (fsm_output(2))) OR
      (fsm_output(7)) OR (fsm_output(9)) OR (fsm_output(5)) OR not_tmp_390);
  mux_2096_nl <= MUX_s_1_2_2(nor_789_nl, nor_790_nl, fsm_output(8));
  nor_791_nl <= NOT((NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (fsm_output(6)) AND (fsm_output(4)) AND (NOT (fsm_output(2))) AND (fsm_output(7))
      AND (NOT (fsm_output(9))))) OR not_tmp_248);
  nor_792_nl <= NOT((fsm_output(4)) OR (fsm_output(2)) OR (fsm_output(7)) OR (NOT
      (fsm_output(9))) OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1111")) OR (fsm_output(10)));
  nor_793_nl <= NOT((NOT (fsm_output(2))) OR (fsm_output(7)) OR (fsm_output(9)) OR
      (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("1111")) OR (fsm_output(10)));
  nor_794_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1111"))
      OR (NOT (fsm_output(2))) OR (fsm_output(7)) OR (NOT (fsm_output(9))) OR (fsm_output(5))
      OR (fsm_output(10)));
  mux_2091_nl <= MUX_s_1_2_2(nor_793_nl, nor_794_nl, fsm_output(4));
  mux_2092_nl <= MUX_s_1_2_2(nor_792_nl, mux_2091_nl, fsm_output(6));
  mux_2093_nl <= MUX_s_1_2_2(nor_791_nl, mux_2092_nl, fsm_output(8));
  mux_2097_nl <= MUX_s_1_2_2(mux_2096_nl, mux_2093_nl, fsm_output(0));
  nand_215_nl <= NOT((COMP_LOOP_acc_16_psp_sva(0)) AND (fsm_output(4)) AND (fsm_output(2))
      AND (VEC_LOOP_j_sva_11_0(2)) AND (fsm_output(7)) AND CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1
      DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND (fsm_output(9)) AND (fsm_output(5))
      AND (NOT (fsm_output(10))));
  or_2261_nl <= CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR (fsm_output(2)) OR (fsm_output(7)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("11")) OR (fsm_output(9)) OR (fsm_output(5)) OR
      (NOT (fsm_output(10)));
  mux_2088_nl <= MUX_s_1_2_2(mux_tmp_2076, or_2261_nl, fsm_output(4));
  mux_2089_nl <= MUX_s_1_2_2(nand_215_nl, mux_2088_nl, fsm_output(6));
  and_555_nl <= (fsm_output(8)) AND (NOT mux_2089_nl);
  nand_395_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (fsm_output(2)) AND (fsm_output(7)) AND (fsm_output(9)) AND (NOT (fsm_output(5)))
      AND (fsm_output(10)));
  or_2256_nl <= (fsm_output(7)) OR (NOT nor_tmp_265);
  mux_2085_nl <= MUX_s_1_2_2(or_2256_nl, or_tmp_2192, fsm_output(2));
  mux_2086_nl <= MUX_s_1_2_2(nand_395_nl, mux_2085_nl, fsm_output(4));
  nor_795_nl <= NOT((fsm_output(6)) OR mux_2086_nl);
  nor_796_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1111"))
      OR (fsm_output(6)) OR (NOT (fsm_output(4))) OR (fsm_output(2)) OR (NOT (fsm_output(7)))
      OR (fsm_output(9)) OR (NOT (fsm_output(5))) OR (fsm_output(10)));
  mux_2087_nl <= MUX_s_1_2_2(nor_795_nl, nor_796_nl, fsm_output(8));
  mux_2090_nl <= MUX_s_1_2_2(and_555_nl, mux_2087_nl, fsm_output(0));
  mux_2098_nl <= MUX_s_1_2_2(mux_2097_nl, mux_2090_nl, fsm_output(3));
  or_2253_nl <= (NOT(CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"))
      AND (fsm_output(2)) AND (NOT (fsm_output(7))))) OR nand_334_cse;
  or_2251_nl <= (NOT (fsm_output(2))) OR (fsm_output(7)) OR (fsm_output(9)) OR not_tmp_387;
  mux_2081_nl <= MUX_s_1_2_2(or_2253_nl, or_2251_nl, fsm_output(4));
  nor_797_nl <= NOT((fsm_output(6)) OR mux_2081_nl);
  or_2245_nl <= (fsm_output(9)) OR (fsm_output(5)) OR not_tmp_390;
  mux_2079_nl <= MUX_s_1_2_2(or_702_cse, or_2245_nl, fsm_output(7));
  mux_2080_nl <= MUX_s_1_2_2(or_tmp_2192, mux_2079_nl, and_564_cse);
  nor_798_nl <= NOT((NOT (fsm_output(6))) OR (NOT (fsm_output(4))) OR (fsm_output(2))
      OR mux_2080_nl);
  mux_2082_nl <= MUX_s_1_2_2(nor_797_nl, nor_798_nl, fsm_output(8));
  or_2241_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1111"))
      OR (fsm_output(7)) OR (fsm_output(9)) OR not_tmp_248;
  nand_219_nl <= NOT((fsm_output(7)) AND CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3
      DOWNTO 0)=STD_LOGIC_VECTOR'("1111")) AND (fsm_output(9)) AND (NOT (fsm_output(5)))
      AND (NOT (fsm_output(10))));
  mux_2077_nl <= MUX_s_1_2_2(or_2241_nl, nand_219_nl, fsm_output(2));
  mux_2078_nl <= MUX_s_1_2_2(mux_2077_nl, mux_tmp_2076, fsm_output(4));
  nor_799_nl <= NOT((fsm_output(8)) OR (fsm_output(6)) OR mux_2078_nl);
  mux_2083_nl <= MUX_s_1_2_2(mux_2082_nl, nor_799_nl, fsm_output(0));
  or_2234_nl <= CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("111"))
      OR (fsm_output(2)) OR (NOT (fsm_output(7))) OR (NOT (VEC_LOOP_j_sva_11_0(0)))
      OR (fsm_output(9)) OR (fsm_output(5)) OR (NOT (fsm_output(10)));
  or_2232_nl <= (fsm_output(2)) OR (NOT (fsm_output(7))) OR (NOT (fsm_output(9)))
      OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("1111")) OR (fsm_output(10));
  mux_2073_nl <= MUX_s_1_2_2(or_2234_nl, or_2232_nl, fsm_output(4));
  nand_220_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"))
      AND (fsm_output(2)) AND (fsm_output(7)) AND (VEC_LOOP_j_sva_11_0(0)) AND (fsm_output(9))
      AND (fsm_output(5)) AND (NOT (fsm_output(10))));
  nand_221_nl <= NOT((fsm_output(2)) AND (fsm_output(7)) AND (NOT (fsm_output(9)))
      AND (fsm_output(5)) AND CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO
      0)=STD_LOGIC_VECTOR'("1111")) AND (NOT (fsm_output(10))));
  mux_2072_nl <= MUX_s_1_2_2(nand_220_nl, nand_221_nl, fsm_output(4));
  mux_2074_nl <= MUX_s_1_2_2(mux_2073_nl, mux_2072_nl, fsm_output(6));
  nor_800_nl <= NOT((fsm_output(8)) OR mux_2074_nl);
  nor_801_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1111"))
      OR (NOT (fsm_output(6))) OR (fsm_output(4)) OR (fsm_output(2)) OR (NOT (fsm_output(7)))
      OR (fsm_output(9)) OR (NOT (fsm_output(5))) OR (fsm_output(10)));
  nor_802_nl <= NOT((NOT((fsm_output(4)) AND (fsm_output(2)) AND (fsm_output(7))
      AND CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (NOT (fsm_output(9))))) OR not_tmp_248);
  or_2225_nl <= (fsm_output(7)) OR (fsm_output(9)) OR not_tmp_387;
  nand_223_nl <= NOT((fsm_output(7)) AND (fsm_output(9)) AND (NOT (fsm_output(5)))
      AND CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (NOT (fsm_output(10))));
  mux_2069_nl <= MUX_s_1_2_2(or_2225_nl, nand_223_nl, fsm_output(2));
  nor_803_nl <= NOT((fsm_output(4)) OR mux_2069_nl);
  mux_2070_nl <= MUX_s_1_2_2(nor_802_nl, nor_803_nl, fsm_output(6));
  mux_2071_nl <= MUX_s_1_2_2(nor_801_nl, mux_2070_nl, fsm_output(8));
  mux_2075_nl <= MUX_s_1_2_2(nor_800_nl, mux_2071_nl, fsm_output(0));
  mux_2084_nl <= MUX_s_1_2_2(mux_2083_nl, mux_2075_nl, fsm_output(3));
  vec_rsc_0_15_i_wea_d_pff <= MUX_s_1_2_2(mux_2098_nl, mux_2084_nl, fsm_output(1));
  nand_199_nl <= NOT((fsm_output(7)) AND CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (NOT (fsm_output(3))) AND (fsm_output(9)) AND (fsm_output(2)) AND (NOT
      (fsm_output(10))));
  or_2327_nl <= (fsm_output(7)) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1111"))
      OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(2)) OR (NOT (fsm_output(10)));
  mux_2129_nl <= MUX_s_1_2_2(nand_199_nl, or_2327_nl, fsm_output(5));
  nor_763_nl <= NOT((fsm_output(1)) OR mux_2129_nl);
  nor_764_nl <= NOT((fsm_output(5)) OR (NOT (fsm_output(7))) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1111")) OR (fsm_output(3)) OR (fsm_output(9))
      OR (fsm_output(2)) OR (fsm_output(10)));
  nor_765_nl <= NOT((NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (fsm_output(7)) AND (NOT (fsm_output(3))) AND (NOT (fsm_output(9))))) OR
      not_tmp_253);
  nor_766_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1111"))
      OR (fsm_output(7)) OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (fsm_output(2))
      OR (NOT (fsm_output(10))));
  mux_2127_nl <= MUX_s_1_2_2(nor_765_nl, nor_766_nl, fsm_output(5));
  mux_2128_nl <= MUX_s_1_2_2(nor_764_nl, mux_2127_nl, fsm_output(1));
  mux_2130_nl <= MUX_s_1_2_2(nor_763_nl, mux_2128_nl, fsm_output(0));
  and_546_nl <= (fsm_output(6)) AND mux_2130_nl;
  nor_767_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1111"))
      OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR (fsm_output(2)) OR (fsm_output(10)));
  nor_769_nl <= NOT((NOT((NOT (fsm_output(7))) AND CONV_SL_1_1(z_out_2_12_1(3 DOWNTO
      0)=STD_LOGIC_VECTOR'("1111")) AND (fsm_output(3)) AND (NOT (fsm_output(9)))))
      OR not_tmp_253);
  mux_2122_nl <= MUX_s_1_2_2(nor_1445_cse, nor_769_nl, fsm_output(5));
  nor_770_nl <= NOT((NOT((fsm_output(5)) AND (NOT (fsm_output(7))) AND CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)=STD_LOGIC_VECTOR'("1111")) AND (fsm_output(3)) AND (NOT (fsm_output(9)))))
      OR not_tmp_253);
  nand_203_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm);
  mux_2123_nl <= MUX_s_1_2_2(mux_2122_nl, nor_770_nl, nand_203_nl);
  mux_2124_nl <= MUX_s_1_2_2(nor_767_nl, mux_2123_nl, fsm_output(1));
  nor_771_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11")) OR
      (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_253);
  and_547_nl <= CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111")) AND
      (fsm_output(7)) AND (fsm_output(3)) AND (NOT (fsm_output(9))) AND (fsm_output(2))
      AND (NOT (fsm_output(10)));
  nor_772_nl <= NOT((fsm_output(7)) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1111"))
      OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9))) OR (fsm_output(2)) OR (fsm_output(10)));
  mux_2120_nl <= MUX_s_1_2_2(and_547_nl, nor_772_nl, fsm_output(5));
  mux_2121_nl <= MUX_s_1_2_2(nor_771_nl, mux_2120_nl, fsm_output(1));
  mux_2125_nl <= MUX_s_1_2_2(mux_2124_nl, mux_2121_nl, fsm_output(0));
  nor_773_nl <= NOT((NOT(COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm AND (fsm_output(5))
      AND (NOT (fsm_output(7))) AND CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO
      0)=STD_LOGIC_VECTOR'("1111")) AND (fsm_output(3)) AND (NOT (fsm_output(9)))))
      OR not_tmp_253);
  nor_774_nl <= NOT((NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (NOT (fsm_output(5)))
      OR (fsm_output(7)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1111"))
      OR (fsm_output(3)) OR (fsm_output(9)) OR (NOT (fsm_output(2))) OR (fsm_output(10)));
  mux_2118_nl <= MUX_s_1_2_2(nor_773_nl, nor_774_nl, fsm_output(1));
  nor_775_nl <= NOT(nand_324_cse OR mux_1925_cse);
  mux_2119_nl <= MUX_s_1_2_2(mux_2118_nl, nor_775_nl, fsm_output(0));
  mux_2126_nl <= MUX_s_1_2_2(mux_2125_nl, mux_2119_nl, fsm_output(6));
  mux_2131_nl <= MUX_s_1_2_2(and_546_nl, mux_2126_nl, fsm_output(8));
  nor_776_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1111"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (fsm_output(2))
      OR (fsm_output(10)));
  nor_777_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1111"))
      OR (fsm_output(7)) OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(2)))
      OR (fsm_output(10)));
  mux_2112_nl <= MUX_s_1_2_2(nor_776_nl, nor_777_nl, fsm_output(5));
  and_548_nl <= COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm AND mux_2112_nl;
  nor_778_nl <= NOT((NOT((fsm_output(7)) AND CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3
      DOWNTO 0)=STD_LOGIC_VECTOR'("1111")) AND (fsm_output(3)) AND (NOT (fsm_output(9)))))
      OR not_tmp_253);
  and_759_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (NOT (fsm_output(7))) AND (fsm_output(3)) AND (fsm_output(9)) AND (NOT
      (fsm_output(2))) AND (fsm_output(10));
  mux_2111_nl <= MUX_s_1_2_2(nor_778_nl, and_759_nl, fsm_output(5));
  and_549_nl <= COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm AND mux_2111_nl;
  mux_2113_nl <= MUX_s_1_2_2(and_548_nl, and_549_nl, fsm_output(1));
  nor_780_nl <= NOT((NOT (VEC_LOOP_j_sva_11_0(3))) OR (NOT (VEC_LOOP_j_sva_11_0(1)))
      OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR (NOT (fsm_output(5))) OR (fsm_output(7))
      OR (NOT (VEC_LOOP_j_sva_11_0(2))) OR (fsm_output(3)) OR (fsm_output(9)) OR
      (fsm_output(2)) OR (fsm_output(10)));
  nor_781_nl <= NOT(nand_332_cse OR mux_2045_cse);
  mux_2110_nl <= MUX_s_1_2_2(nor_780_nl, nor_781_nl, fsm_output(1));
  mux_2114_nl <= MUX_s_1_2_2(mux_2113_nl, mux_2110_nl, fsm_output(0));
  nor_782_nl <= NOT((NOT (fsm_output(1))) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1111"))
      OR (fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR (fsm_output(2)) OR (fsm_output(10)));
  and_550_nl <= (NOT (fsm_output(5))) AND (NOT (fsm_output(7))) AND (fsm_output(3))
      AND CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111")) AND (fsm_output(9))
      AND (fsm_output(2)) AND (NOT (fsm_output(10)));
  and_551_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"))
      AND (VEC_LOOP_j_sva_11_0(0)) AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm AND (fsm_output(5))
      AND (fsm_output(7)) AND (fsm_output(3)) AND (NOT (fsm_output(9))) AND (fsm_output(2))
      AND (NOT (fsm_output(10)));
  mux_2107_nl <= MUX_s_1_2_2(and_550_nl, and_551_nl, fsm_output(1));
  mux_2108_nl <= MUX_s_1_2_2(nor_782_nl, mux_2107_nl, fsm_output(0));
  mux_2115_nl <= MUX_s_1_2_2(mux_2114_nl, mux_2108_nl, fsm_output(6));
  nor_783_nl <= NOT((NOT (fsm_output(1))) OR CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1111"))
      OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(3)) OR (NOT (fsm_output(9)))
      OR (fsm_output(2)) OR (fsm_output(10)));
  nor_784_nl <= NOT((fsm_output(1)) OR (fsm_output(5)) OR CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1111")) OR (NOT (fsm_output(7))) OR (fsm_output(3))
      OR (fsm_output(9)) OR not_tmp_253);
  mux_2105_nl <= MUX_s_1_2_2(nor_783_nl, nor_784_nl, fsm_output(0));
  nor_785_nl <= NOT((NOT((fsm_output(5)) AND (fsm_output(7)) AND CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)=STD_LOGIC_VECTOR'("1111")) AND (fsm_output(3)) AND (NOT (fsm_output(9)))))
      OR not_tmp_253);
  nor_786_nl <= NOT((NOT (fsm_output(7))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1111")) OR (fsm_output(3)) OR (NOT (fsm_output(9)))
      OR (fsm_output(2)) OR (fsm_output(10)));
  nor_787_nl <= NOT((NOT((fsm_output(7)) AND CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (fsm_output(3)) AND (NOT (fsm_output(9))))) OR not_tmp_253);
  mux_2101_nl <= MUX_s_1_2_2(nor_786_nl, nor_787_nl, fsm_output(5));
  mux_2102_nl <= MUX_s_1_2_2(nor_785_nl, mux_2101_nl, COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm);
  and_552_nl <= (fsm_output(5)) AND (fsm_output(7)) AND CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)=STD_LOGIC_VECTOR'("1111")) AND (NOT (fsm_output(3))) AND (NOT (fsm_output(9)))
      AND (fsm_output(2)) AND (NOT (fsm_output(10)));
  mux_2103_nl <= MUX_s_1_2_2(mux_2102_nl, and_552_nl, fsm_output(1));
  and_553_nl <= (fsm_output(5)) AND (fsm_output(7)) AND CONV_SL_1_1(z_out_2_12_1(3
      DOWNTO 0)=STD_LOGIC_VECTOR'("1111")) AND (fsm_output(3)) AND (fsm_output(9))
      AND (NOT (fsm_output(2))) AND (NOT (fsm_output(10)));
  nor_788_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("111"))
      OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(3)) OR (fsm_output(9))
      OR (fsm_output(2)) OR (NOT (fsm_output(10))));
  mux_2100_nl <= MUX_s_1_2_2(and_553_nl, nor_788_nl, fsm_output(1));
  mux_2104_nl <= MUX_s_1_2_2(mux_2103_nl, mux_2100_nl, fsm_output(0));
  mux_2106_nl <= MUX_s_1_2_2(mux_2105_nl, mux_2104_nl, fsm_output(6));
  mux_2116_nl <= MUX_s_1_2_2(mux_2115_nl, mux_2106_nl, fsm_output(8));
  vec_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_2131_nl, mux_2116_nl,
      fsm_output(4));
  and_dcpl_332 <= CONV_SL_1_1(fsm_output=STD_LOGIC_VECTOR'("11010100010"));
  and_dcpl_333 <= (NOT (fsm_output(6))) AND (fsm_output(0));
  and_dcpl_338 <= (NOT (fsm_output(3))) AND (fsm_output(5)) AND (NOT (fsm_output(8)));
  and_dcpl_340 <= NOT((fsm_output(2)) OR (fsm_output(9)) OR (fsm_output(10)));
  and_dcpl_342 <= and_dcpl_340 AND and_dcpl_338 AND (fsm_output(4)) AND (NOT (fsm_output(7)))
      AND (NOT (fsm_output(1))) AND and_dcpl_333;
  and_dcpl_344 <= NOT((fsm_output(4)) OR (fsm_output(7)));
  and_dcpl_345 <= and_dcpl_344 AND (fsm_output(1));
  and_dcpl_349 <= and_dcpl_340 AND (fsm_output(3)) AND (NOT (fsm_output(5))) AND
      (NOT (fsm_output(8)));
  and_dcpl_350 <= and_dcpl_349 AND and_dcpl_345 AND (NOT (fsm_output(6))) AND (NOT
      (fsm_output(0)));
  and_dcpl_356 <= (NOT (fsm_output(2))) AND (fsm_output(9)) AND (fsm_output(10))
      AND and_dcpl_338 AND and_dcpl_345 AND (fsm_output(6)) AND (fsm_output(0));
  and_dcpl_359 <= and_dcpl_349 AND and_dcpl_344 AND (NOT (fsm_output(1))) AND and_dcpl_333;
  and_815_cse <= (fsm_output(6)) AND (NOT (fsm_output(0)));
  and_816_cse <= (fsm_output(4)) AND (NOT (fsm_output(7)));
  and_820_cse <= and_dcpl_114 AND (NOT (fsm_output(8)));
  and_dcpl_367 <= nor_609_cse AND (NOT (fsm_output(2)));
  and_825_cse <= (fsm_output(6)) AND (fsm_output(0));
  and_dcpl_371 <= (NOT (fsm_output(4))) AND (fsm_output(7));
  and_827_cse <= and_dcpl_371 AND (NOT (fsm_output(1)));
  and_830_cse <= and_dcpl_91 AND (NOT (fsm_output(8)));
  nor_1670_cse <= NOT((fsm_output(6)) OR (fsm_output(0)));
  and_835_cse <= and_dcpl_344 AND (NOT (fsm_output(1)));
  and_dcpl_383 <= (fsm_output(3)) AND (fsm_output(5)) AND (fsm_output(8));
  and_842_cse <= and_dcpl_371 AND (fsm_output(1));
  and_dcpl_390 <= nor_609_cse AND (fsm_output(2));
  and_dcpl_393 <= (fsm_output(4)) AND (fsm_output(7));
  and_849_cse <= and_dcpl_393 AND (fsm_output(1));
  and_dcpl_403 <= and_dcpl_33 AND (fsm_output(2));
  and_dcpl_411 <= and_dcpl_33 AND (NOT (fsm_output(2)));
  and_dcpl_412 <= and_dcpl_411 AND and_dcpl_383;
  and_870_cse <= and_dcpl_91 AND (fsm_output(8));
  and_873_cse <= and_dcpl_393 AND (NOT (fsm_output(1)));
  and_dcpl_422 <= and_dcpl_39 AND (NOT (fsm_output(8)));
  and_dcpl_428 <= and_dcpl_59 AND (fsm_output(2));
  and_dcpl_432 <= and_dcpl_428 AND and_dcpl_383;
  and_dcpl_446 <= and_816_cse AND (NOT (fsm_output(1)));
  and_dcpl_453 <= and_dcpl_340 AND and_dcpl_39 AND (NOT (fsm_output(8))) AND and_dcpl_446
      AND and_dcpl_333;
  and_dcpl_460 <= and_dcpl_340 AND and_820_cse AND and_816_cse AND (fsm_output(1))
      AND and_815_cse;
  and_dcpl_468 <= and_dcpl_340 AND and_830_cse AND and_dcpl_371 AND (NOT (fsm_output(1)))
      AND and_825_cse;
  and_dcpl_472 <= (fsm_output(2)) AND (NOT (fsm_output(9)));
  and_dcpl_473 <= and_dcpl_472 AND (NOT (fsm_output(10)));
  and_dcpl_475 <= and_dcpl_473 AND and_dcpl_114 AND (fsm_output(8)) AND and_842_cse
      AND and_dcpl_333;
  and_dcpl_481 <= and_dcpl_473 AND and_dcpl_39 AND (fsm_output(8)) AND and_849_cse
      AND and_815_cse;
  and_dcpl_486 <= (fsm_output(2)) AND (fsm_output(9)) AND (NOT (fsm_output(10)))
      AND and_820_cse AND and_dcpl_446 AND and_825_cse;
  and_dcpl_488 <= (NOT (fsm_output(4))) AND (NOT (fsm_output(7))) AND (fsm_output(1));
  and_dcpl_493 <= (NOT (fsm_output(2))) AND (fsm_output(9)) AND (NOT (fsm_output(10)));
  and_dcpl_494 <= and_dcpl_493 AND and_dcpl_383;
  and_dcpl_495 <= and_dcpl_494 AND and_dcpl_488 AND and_dcpl_333;
  and_dcpl_500 <= and_dcpl_493 AND and_870_cse AND and_849_cse AND nor_1670_cse;
  and_dcpl_503 <= and_dcpl_494 AND and_873_cse AND and_825_cse;
  and_dcpl_505 <= and_dcpl_472 AND (fsm_output(10));
  and_dcpl_507 <= and_dcpl_505 AND and_830_cse AND and_842_cse AND and_825_cse;
  and_dcpl_510 <= and_dcpl_505 AND and_dcpl_383 AND and_dcpl_488 AND nor_1670_cse;
  and_dcpl_513 <= and_dcpl_505 AND and_870_cse AND and_873_cse AND and_dcpl_333;
  and_dcpl_531 <= nor_609_cse AND (fsm_output(2)) AND and_dcpl_39 AND (fsm_output(8))
      AND and_dcpl_393 AND (fsm_output(1)) AND (fsm_output(6)) AND (NOT (fsm_output(0)));
  and_dcpl_539 <= (NOT (fsm_output(10))) AND (fsm_output(9)) AND (NOT (fsm_output(2)))
      AND and_dcpl_383;
  and_dcpl_540 <= and_dcpl_539 AND and_dcpl_488 AND and_dcpl_333;
  and_dcpl_544 <= and_dcpl_539 AND and_873_cse AND and_825_cse;
  and_dcpl_551 <= (fsm_output(10)) AND (NOT (fsm_output(9))) AND (fsm_output(2));
  and_dcpl_553 <= and_dcpl_551 AND and_dcpl_91 AND (NOT (fsm_output(8))) AND (NOT
      (fsm_output(4))) AND (fsm_output(7)) AND (fsm_output(1)) AND and_825_cse;
  and_dcpl_557 <= and_dcpl_551 AND and_dcpl_383 AND and_dcpl_488 AND (NOT (fsm_output(6)))
      AND (NOT (fsm_output(0)));
  and_dcpl_561 <= and_dcpl_551 AND and_dcpl_91 AND (fsm_output(8)) AND and_873_cse
      AND and_dcpl_333;
  and_dcpl_567 <= NOT((fsm_output(3)) OR (fsm_output(5)) OR (fsm_output(8)));
  and_dcpl_568 <= NOT((fsm_output(2)) OR (fsm_output(9)));
  and_dcpl_569 <= and_dcpl_568 AND (NOT (fsm_output(10)));
  and_dcpl_594 <= (fsm_output(2)) AND (fsm_output(9)) AND (NOT (fsm_output(10)));
  and_dcpl_627 <= and_dcpl_340 AND and_dcpl_338;
  and_dcpl_628 <= and_dcpl_627 AND and_816_cse AND (NOT (fsm_output(1))) AND and_dcpl_333;
  and_dcpl_631 <= NOT((fsm_output(4)) OR (fsm_output(7)) OR (fsm_output(1)));
  and_dcpl_636 <= and_dcpl_340 AND (fsm_output(3)) AND (fsm_output(5)) AND (fsm_output(8))
      AND and_dcpl_631 AND (NOT (fsm_output(6))) AND (NOT (fsm_output(0)));
  and_dcpl_642 <= (fsm_output(10)) AND (NOT (fsm_output(9))) AND (NOT (fsm_output(2)))
      AND and_dcpl_338 AND and_dcpl_631 AND (fsm_output(6)) AND (NOT (fsm_output(0)));
  or_tmp_3282 <= (fsm_output(1)) OR (NOT (fsm_output(2))) OR (NOT (fsm_output(9)))
      OR (fsm_output(8)) OR (fsm_output(6));
  not_tmp_834 <= NOT((fsm_output(8)) AND (fsm_output(6)));
  not_tmp_835 <= NOT((fsm_output(9)) AND (fsm_output(8)) AND (fsm_output(6)));
  nor_1657_cse <= NOT((fsm_output(3)) OR (fsm_output(4)) OR (NOT (fsm_output(10)))
      OR (fsm_output(0)) OR (fsm_output(1)) OR (fsm_output(2)) OR (fsm_output(9))
      OR (fsm_output(8)) OR (fsm_output(6)));
  or_3467_nl <= (fsm_output(1)) OR (NOT (fsm_output(2))) OR (NOT (fsm_output(9)))
      OR (NOT (fsm_output(8))) OR (fsm_output(6));
  or_3466_nl <= (fsm_output(1)) OR (fsm_output(2)) OR (fsm_output(9)) OR (NOT (fsm_output(8)))
      OR (fsm_output(6));
  mux_3809_nl <= MUX_s_1_2_2(or_3467_nl, or_3466_nl, fsm_output(0));
  or_3465_nl <= (NOT (fsm_output(0))) OR (NOT (fsm_output(1))) OR (NOT (fsm_output(2)))
      OR (fsm_output(9)) OR (NOT (fsm_output(8))) OR (fsm_output(6));
  mux_3810_nl <= MUX_s_1_2_2(mux_3809_nl, or_3465_nl, fsm_output(10));
  nor_1648_nl <= NOT(CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("00"))
      OR mux_3810_nl);
  nor_1649_nl <= NOT((NOT (fsm_output(4))) OR (fsm_output(10)) OR (fsm_output(0))
      OR (NOT (fsm_output(1))) OR (NOT (fsm_output(2))) OR (NOT (fsm_output(9)))
      OR (fsm_output(8)) OR (fsm_output(6)));
  nor_1650_nl <= NOT((fsm_output(1)) OR (fsm_output(2)) OR (fsm_output(9)) OR not_tmp_834);
  nor_1651_nl <= NOT(CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("01"))
      OR not_tmp_835);
  mux_3805_nl <= MUX_s_1_2_2(nor_1650_nl, nor_1651_nl, fsm_output(0));
  nor_1652_nl <= NOT((fsm_output(0)) OR (NOT (fsm_output(1))) OR (NOT (fsm_output(2)))
      OR (fsm_output(9)) OR not_tmp_834);
  mux_3806_nl <= MUX_s_1_2_2(mux_3805_nl, nor_1652_nl, fsm_output(10));
  or_3456_nl <= (fsm_output(1)) OR (fsm_output(2)) OR (fsm_output(9)) OR (fsm_output(8))
      OR (fsm_output(6));
  mux_3804_nl <= MUX_s_1_2_2(or_tmp_3282, or_3456_nl, fsm_output(0));
  and_nl <= (fsm_output(10)) AND (NOT mux_3804_nl);
  mux_3807_nl <= MUX_s_1_2_2(mux_3806_nl, and_nl, fsm_output(4));
  mux_3808_nl <= MUX_s_1_2_2(nor_1649_nl, mux_3807_nl, fsm_output(3));
  mux_3811_nl <= MUX_s_1_2_2(nor_1648_nl, mux_3808_nl, fsm_output(5));
  nor_1653_nl <= NOT(CONV_SL_1_1(fsm_output(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR not_tmp_835);
  nor_1654_nl <= NOT((NOT (fsm_output(0))) OR (fsm_output(1)) OR (NOT (fsm_output(2)))
      OR (fsm_output(9)) OR not_tmp_834);
  mux_3801_nl <= MUX_s_1_2_2(nor_1653_nl, nor_1654_nl, fsm_output(10));
  and_1158_nl <= (fsm_output(4)) AND mux_3801_nl;
  nor_1655_nl <= NOT((fsm_output(10)) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(1)))
      OR (NOT (fsm_output(2))) OR (fsm_output(9)) OR not_tmp_834);
  or_3448_nl <= (NOT (fsm_output(1))) OR (fsm_output(2)) OR (fsm_output(9)) OR (fsm_output(8))
      OR (fsm_output(6));
  mux_3828_nl <= MUX_s_1_2_2(or_3448_nl, or_tmp_3282, fsm_output(0));
  nor_1656_nl <= NOT((fsm_output(10)) OR mux_3828_nl);
  mux_3800_nl <= MUX_s_1_2_2(nor_1655_nl, nor_1656_nl, fsm_output(4));
  mux_3802_nl <= MUX_s_1_2_2(and_1158_nl, mux_3800_nl, fsm_output(3));
  mux_3803_nl <= MUX_s_1_2_2(mux_3802_nl, nor_1657_cse, fsm_output(5));
  not_tmp_838 <= MUX_s_1_2_2(mux_3811_nl, mux_3803_nl, fsm_output(7));
  and_dcpl_647 <= and_dcpl_340 AND (NOT (fsm_output(3))) AND (NOT (fsm_output(5)))
      AND (NOT (fsm_output(8))) AND and_dcpl_631 AND and_dcpl_333;
  and_dcpl_650 <= and_dcpl_627 AND and_816_cse AND (fsm_output(1)) AND and_dcpl_333;
  and_dcpl_660 <= (fsm_output(2)) AND (fsm_output(9)) AND (NOT (fsm_output(10)))
      AND and_dcpl_91 AND (NOT (fsm_output(8))) AND (NOT (fsm_output(4))) AND (fsm_output(7))
      AND (NOT (fsm_output(1))) AND and_815_cse;
  and_dcpl_669 <= (fsm_output(2)) AND (NOT (fsm_output(9))) AND (fsm_output(10))
      AND (fsm_output(3)) AND (fsm_output(5)) AND (fsm_output(8)) AND and_dcpl_393
      AND (NOT (fsm_output(1))) AND and_815_cse;
  and_dcpl_678 <= (NOT (fsm_output(2))) AND (NOT (fsm_output(9))) AND (NOT (fsm_output(10)))
      AND (fsm_output(3)) AND (NOT (fsm_output(5))) AND (NOT (fsm_output(8))) AND
      (fsm_output(4)) AND (NOT (fsm_output(7))) AND (fsm_output(1)) AND and_815_cse;
  and_dcpl_686 <= (NOT (fsm_output(2))) AND (fsm_output(9)) AND (NOT (fsm_output(10)))
      AND and_dcpl_91 AND (fsm_output(8)) AND and_dcpl_393 AND (fsm_output(1)) AND
      (NOT (fsm_output(6))) AND (NOT (fsm_output(0)));
  or_tmp_3307 <= (NOT (fsm_output(9))) OR (fsm_output(10)) OR (fsm_output(1)) OR
      (NOT (fsm_output(2)));
  or_tmp_3312 <= (NOT (fsm_output(9))) OR (fsm_output(10)) OR (NOT (fsm_output(1)))
      OR (fsm_output(2));
  mux_3821_nl <= MUX_s_1_2_2(nor_758_cse, and_529_cse, fsm_output(10));
  or_tmp_3326 <= (fsm_output(9)) OR (NOT mux_3821_nl);
  and_978_ssc <= nor_609_cse AND (NOT (fsm_output(2))) AND and_dcpl_39 AND (NOT (fsm_output(8)))
      AND (fsm_output(4)) AND (NOT (fsm_output(7))) AND (NOT (fsm_output(1))) AND
      and_dcpl_333;
  and_824_ssc <= and_dcpl_367 AND and_820_cse AND and_816_cse AND (fsm_output(1))
      AND and_815_cse;
  COMP_LOOP_or_54_ssc <= (and_dcpl_367 AND and_830_cse AND and_827_cse AND and_825_cse)
      OR (and_dcpl_367 AND and_dcpl_383 AND and_835_cse AND nor_1670_cse) OR (and_dcpl_390
      AND and_dcpl_114 AND (fsm_output(8)) AND and_842_cse AND and_dcpl_333) OR (and_dcpl_403
      AND and_820_cse AND and_816_cse AND (NOT (fsm_output(1))) AND and_825_cse)
      OR (and_dcpl_403 AND and_830_cse AND and_827_cse AND and_815_cse) OR (and_dcpl_59
      AND (NOT (fsm_output(2))) AND and_dcpl_422 AND and_835_cse AND and_815_cse)
      OR (and_dcpl_432 AND and_873_cse AND and_815_cse) OR ((fsm_output(10)) AND
      (fsm_output(9)) AND (NOT (fsm_output(2))) AND and_dcpl_422 AND and_dcpl_345
      AND and_825_cse);
  COMP_LOOP_or_55_ssc <= (and_dcpl_390 AND and_dcpl_39 AND (fsm_output(8)) AND and_849_cse
      AND and_815_cse) OR (and_dcpl_412 AND and_dcpl_345 AND and_dcpl_333) OR (and_dcpl_412
      AND and_873_cse AND and_825_cse) OR (and_dcpl_428 AND and_830_cse AND and_842_cse
      AND and_825_cse) OR (and_dcpl_432 AND and_dcpl_345 AND nor_1670_cse) OR (and_dcpl_428
      AND and_870_cse AND and_873_cse AND and_dcpl_333);
  and_872_ssc <= and_dcpl_411 AND and_870_cse AND and_849_cse AND nor_1670_cse;
  mux_3829_nl <= MUX_s_1_2_2(mux_tmp_227, or_tmp_104, and_526_cse);
  or_3510_nl <= (fsm_output(1)) OR (fsm_output(9)) OR (NOT (fsm_output(10)));
  mux_tmp_3828 <= MUX_s_1_2_2(mux_3829_nl, or_3510_nl, fsm_output(2));
  mux_tmp_3830 <= MUX_s_1_2_2(mux_tmp_227, or_tmp_104, fsm_output(1));
  nor_tmp_549 <= or_2400_cse AND (fsm_output(10));
  or_tmp_3337 <= nor_753_cse OR CONV_SL_1_1(fsm_output(10 DOWNTO 9)/=STD_LOGIC_VECTOR'("00"));
  or_tmp_3339 <= nor_297_cse OR (fsm_output(10));
  mux_tmp_3839 <= MUX_s_1_2_2(or_tmp_3339, and_757_cse, or_2644_cse);
  mux_3842_nl <= MUX_s_1_2_2(and_757_cse, mux_tmp_227, or_3388_cse);
  or_3520_nl <= and_526_cse OR CONV_SL_1_1(fsm_output(10 DOWNTO 9)/=STD_LOGIC_VECTOR'("10"));
  mux_tmp_3841 <= MUX_s_1_2_2(mux_3842_nl, or_3520_nl, fsm_output(2));
  or_tmp_3344 <= (NOT (fsm_output(3))) OR (NOT (fsm_output(2))) OR (NOT (fsm_output(1)))
      OR (fsm_output(9)) OR (fsm_output(10));
  nor_tmp_552 <= or_2421_cse AND (fsm_output(10));
  or_tmp_3347 <= nor_303_cse OR (fsm_output(10));
  or_3527_nl <= (NOT (fsm_output(2))) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(1)))
      OR (fsm_output(9)) OR (fsm_output(10));
  mux_3849_nl <= MUX_s_1_2_2(or_tmp_3347, nor_tmp_552, fsm_output(2));
  mux_tmp_3848 <= MUX_s_1_2_2(or_3527_nl, mux_3849_nl, fsm_output(3));
  nor_tmp_554 <= or_2419_cse AND (fsm_output(10));
  or_tmp_3352 <= and_521_cse OR (fsm_output(10));
  mux_tmp_3856 <= MUX_s_1_2_2(or_tmp_3352, nor_tmp_554, fsm_output(2));
  mux_tmp_3864 <= MUX_s_1_2_2(or_tmp_3337, nor_tmp_549, fsm_output(2));
  or_tmp_3357 <= (fsm_output(2)) OR and_526_cse OR (NOT and_757_cse);
  nor_1704_cse <= NOT(COMP_LOOP_nor_11_itm OR (fsm_output(6)));
  or_tmp_3381 <= (fsm_output(10)) OR nor_1704_cse OR (fsm_output(2)) OR (NOT (fsm_output(9)));
  or_tmp_3382 <= NOT((fsm_output(10)) AND COMP_LOOP_nor_11_itm AND (fsm_output(6))
      AND (fsm_output(2)) AND (NOT (fsm_output(9))));
  or_tmp_3384 <= nor_1704_cse OR (NOT (fsm_output(2))) OR (fsm_output(9));
  or_3564_nl <= (NOT COMP_LOOP_nor_11_itm) OR (NOT (fsm_output(6))) OR (fsm_output(2))
      OR (fsm_output(9));
  mux_3893_nl <= MUX_s_1_2_2(or_3564_nl, or_tmp_3384, fsm_output(10));
  mux_tmp_3892 <= MUX_s_1_2_2(mux_3893_nl, or_tmp_3382, fsm_output(1));
  not_tmp_882 <= NOT(COMP_LOOP_nor_11_itm AND (fsm_output(6)) AND (fsm_output(2))
      AND (fsm_output(9)));
  not_tmp_883 <= NOT((fsm_output(2)) AND (fsm_output(9)));
  or_tmp_3402 <= (NOT (fsm_output(6))) OR (fsm_output(2)) OR (NOT (fsm_output(9)));
  mux_3904_nl <= MUX_s_1_2_2(not_tmp_883, or_2855_cse, fsm_output(6));
  mux_tmp_3903 <= MUX_s_1_2_2(or_tmp_3402, mux_3904_nl, COMP_LOOP_nor_11_itm);
  or_tmp_3403 <= (fsm_output(10)) OR mux_tmp_3903;
  or_3586_nl <= (fsm_output(6)) OR (fsm_output(2)) OR (fsm_output(9));
  or_3585_nl <= (NOT (fsm_output(6))) OR (NOT (fsm_output(2))) OR (fsm_output(9));
  mux_tmp_3906 <= MUX_s_1_2_2(or_3586_nl, or_3585_nl, fsm_output(10));
  or_3584_nl <= (NOT COMP_LOOP_nor_11_itm) OR (fsm_output(6)) OR (fsm_output(2))
      OR (fsm_output(9));
  or_3583_nl <= (fsm_output(6)) OR (NOT (fsm_output(2))) OR (fsm_output(9));
  mux_3907_nl <= MUX_s_1_2_2(or_3584_nl, or_3583_nl, fsm_output(10));
  mux_tmp_3907 <= MUX_s_1_2_2(mux_tmp_3906, mux_3907_nl, fsm_output(1));
  or_tmp_3409 <= (fsm_output(10)) OR (fsm_output(6)) OR not_tmp_883;
  COMP_LOOP_or_61_itm <= and_dcpl_460 OR and_dcpl_468 OR and_dcpl_475 OR and_dcpl_481
      OR and_dcpl_486 OR and_dcpl_495 OR and_dcpl_500 OR and_dcpl_503 OR and_dcpl_507
      OR and_dcpl_510 OR and_dcpl_513;
  COMP_LOOP_or_24_itm <= and_dcpl_531 OR and_dcpl_540 OR and_dcpl_544 OR and_dcpl_553
      OR and_dcpl_557 OR and_dcpl_561;
  COMP_LOOP_nor_633_itm <= NOT(and_dcpl_628 OR and_dcpl_636 OR and_dcpl_642);
  COMP_LOOP_nor_685_itm <= NOT(and_dcpl_636 OR and_dcpl_642);
  COMP_LOOP_or_65_itm <= and_dcpl_636 OR and_dcpl_642;
  COMP_LOOP_nor_687_itm <= NOT(and_dcpl_636 OR and_dcpl_642 OR not_tmp_838 OR and_dcpl_650);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( not_tmp_208 = '0' ) THEN
        p_sva <= p_rsci_idat;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( ((and_dcpl_93 AND and_dcpl_88) OR STAGE_LOOP_i_3_0_sva_mx0c1) = '1' )
          THEN
        STAGE_LOOP_i_3_0_sva <= MUX_v_4_2_2(STD_LOGIC_VECTOR'( "0001"), STAGE_LOOP_i_3_0_sva_2,
            STAGE_LOOP_i_3_0_sva_mx0c1);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( not_tmp_208 = '0' ) THEN
        r_sva <= r_rsci_idat;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_vec_rsc_triosy_0_15_obj_ld_cse <= '0';
        COMP_LOOP_nor_11_itm <= '0';
        modExp_exp_1_7_1_sva <= '0';
        COMP_LOOP_nor_12_itm <= '0';
        COMP_LOOP_nor_134_itm <= '0';
        COMP_LOOP_nor_137_itm <= '0';
        COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm <= '0';
        COMP_LOOP_COMP_LOOP_nor_1_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_139_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_140_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_141_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_143_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_144_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_145_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_146_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_147_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_148_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_149_itm <= '0';
      ELSE
        reg_vec_rsc_triosy_0_15_obj_ld_cse <= and_dcpl_103 AND and_dcpl_2 AND and_757_cse
            AND (NOT STAGE_LOOP_acc_itm_2_1);
        COMP_LOOP_nor_11_itm <= (COMP_LOOP_mux1h_428_nl AND (mux_2989_nl OR (fsm_output(0))))
            OR (mux_3077_nl AND (fsm_output(0)));
        modExp_exp_1_7_1_sva <= COMP_LOOP_mux1h_464_nl AND mux_3521_nl;
        COMP_LOOP_nor_12_itm <= (COMP_LOOP_mux1h_474_nl AND mux_3542_nl) OR mux_3636_nl;
        COMP_LOOP_nor_134_itm <= (COMP_LOOP_mux1h_477_nl AND mux_3649_nl) OR mux_3656_nl;
        COMP_LOOP_nor_137_itm <= (COMP_LOOP_mux1h_479_nl AND (mux_3663_nl OR (fsm_output(10))))
            OR mux_3670_nl;
        COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm <= COMP_LOOP_mux1h_480_nl AND (NOT and_dcpl_257);
        COMP_LOOP_COMP_LOOP_nor_1_itm <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")));
        COMP_LOOP_COMP_LOOP_and_139_itm <= CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0101"));
        COMP_LOOP_COMP_LOOP_and_140_itm <= CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0110"));
        COMP_LOOP_COMP_LOOP_and_141_itm <= CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0111"));
        COMP_LOOP_COMP_LOOP_and_143_itm <= CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1001"));
        COMP_LOOP_COMP_LOOP_and_144_itm <= CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1010"));
        COMP_LOOP_COMP_LOOP_and_145_itm <= CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1011"));
        COMP_LOOP_COMP_LOOP_and_146_itm <= CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1100"));
        COMP_LOOP_COMP_LOOP_and_147_itm <= CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1101"));
        COMP_LOOP_COMP_LOOP_and_148_itm <= CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1110"));
        COMP_LOOP_COMP_LOOP_and_149_itm <= CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      modulo_result_rem_cmp_a <= MUX1HOT_v_64_6_2(z_out_8, operator_64_false_acc_mut_63_0,
          COMP_LOOP_10_acc_8_itm, COMP_LOOP_1_modExp_1_while_if_mul_mut_1, COMP_LOOP_10_mul_mut,
          COMP_LOOP_1_acc_5_mut_mx0w5, STD_LOGIC_VECTOR'( modulo_result_or_nl & (NOT
          mux_2231_nl) & (NOT mux_2331_nl) & (NOT mux_2346_nl) & (NOT mux_2418_nl)
          & not_tmp_441));
      modulo_result_rem_cmp_b <= p_sva;
      operator_66_true_div_cmp_a <= MUX_v_65_2_2(z_out_6, (operator_64_false_acc_mut_64
          & operator_64_false_acc_mut_63_0), and_dcpl_241);
      operator_66_true_div_cmp_b_9_0 <= MUX_v_10_2_2(STAGE_LOOP_lshift_psp_sva_mx0w0,
          STAGE_LOOP_lshift_psp_sva, and_dcpl_241);
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( mux_2452_nl = '0' ) THEN
        STAGE_LOOP_lshift_psp_sva <= STAGE_LOOP_lshift_psp_sva_mx0w0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( mux_3889_nl = '0' ) THEN
        operator_64_false_acc_mut_64 <= operator_64_false_mux1h_2_rgt(64);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( mux_3943_nl = '0' ) THEN
        operator_64_false_acc_mut_63_0 <= operator_64_false_mux1h_2_rgt(63 DOWNTO
            0);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        VEC_LOOP_j_sva_11_0 <= STD_LOGIC_VECTOR'( "000000000000");
      ELSIF ( (and_dcpl_247 OR VEC_LOOP_j_sva_11_0_mx0c1) = '1' ) THEN
        VEC_LOOP_j_sva_11_0 <= MUX_v_12_2_2(STD_LOGIC_VECTOR'("000000000000"), (z_out(11
            DOWNTO 0)), VEC_LOOP_j_sva_11_0_mx0c1);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_k_9_4_sva_4_0 <= STD_LOGIC_VECTOR'( "00000");
      ELSIF ( (mux_3946_nl AND (NOT((fsm_output(8)) OR (fsm_output(2))))) = '1' )
          THEN
        COMP_LOOP_k_9_4_sva_4_0 <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), (z_out_1(4
            DOWNTO 0)), or_3508_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( ((modExp_while_and_3 OR modExp_while_and_5 OR modExp_result_sva_mx0c0
          OR (NOT mux_2668_nl)) AND (modExp_result_sva_mx0c0 OR modExp_result_and_rgt
          OR modExp_result_and_1_rgt)) = '1' ) THEN
        modExp_result_sva <= MUX1HOT_v_64_3_2(STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000001"),
            modulo_result_rem_cmp_z, modulo_qr_sva_1_mx0w6, STD_LOGIC_VECTOR'( modExp_result_sva_mx0c0
            & modExp_result_and_rgt & modExp_result_and_1_rgt));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        tmp_10_lpi_4_dfm <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
      ELSIF ( (MUX_s_1_2_2(mux_2741_nl, mux_2714_nl, fsm_output(4))) = '1' ) THEN
        tmp_10_lpi_4_dfm <= MUX1HOT_v_64_17_2(('0' & operator_64_false_slc_modExp_exp_63_1_3),
            vec_rsc_0_0_i_qa_d, vec_rsc_0_1_i_qa_d, vec_rsc_0_2_i_qa_d, vec_rsc_0_3_i_qa_d,
            vec_rsc_0_4_i_qa_d, vec_rsc_0_5_i_qa_d, vec_rsc_0_6_i_qa_d, vec_rsc_0_7_i_qa_d,
            vec_rsc_0_8_i_qa_d, vec_rsc_0_9_i_qa_d, vec_rsc_0_10_i_qa_d, vec_rsc_0_11_i_qa_d,
            vec_rsc_0_12_i_qa_d, vec_rsc_0_13_i_qa_d, vec_rsc_0_14_i_qa_d, vec_rsc_0_15_i_qa_d,
            STD_LOGIC_VECTOR'( and_dcpl_247 & COMP_LOOP_or_8_nl & COMP_LOOP_or_9_nl
            & COMP_LOOP_or_10_nl & COMP_LOOP_or_11_nl & COMP_LOOP_or_12_nl & COMP_LOOP_or_13_nl
            & COMP_LOOP_or_14_nl & COMP_LOOP_or_15_nl & COMP_LOOP_or_16_nl & COMP_LOOP_or_17_nl
            & COMP_LOOP_or_18_nl & COMP_LOOP_or_19_nl & COMP_LOOP_or_20_nl & COMP_LOOP_or_21_nl
            & COMP_LOOP_or_22_nl & COMP_LOOP_or_23_nl));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (MUX_s_1_2_2(mux_2981_nl, mux_2925_nl, fsm_output(1))) = '1' ) THEN
        COMP_LOOP_10_mul_mut <= MUX1HOT_v_64_21_2(r_sva, modulo_result_rem_cmp_z,
            modulo_qr_sva_1_mx0w6, modExp_result_sva, vec_rsc_0_0_i_qa_d, vec_rsc_0_1_i_qa_d,
            vec_rsc_0_2_i_qa_d, vec_rsc_0_3_i_qa_d, vec_rsc_0_4_i_qa_d, vec_rsc_0_5_i_qa_d,
            vec_rsc_0_6_i_qa_d, vec_rsc_0_7_i_qa_d, vec_rsc_0_8_i_qa_d, vec_rsc_0_9_i_qa_d,
            vec_rsc_0_10_i_qa_d, vec_rsc_0_11_i_qa_d, vec_rsc_0_12_i_qa_d, vec_rsc_0_13_i_qa_d,
            vec_rsc_0_14_i_qa_d, vec_rsc_0_15_i_qa_d, COMP_LOOP_1_modExp_1_while_if_mul_mut_1,
            STD_LOGIC_VECTOR'( and_312_nl & COMP_LOOP_or_29_nl & COMP_LOOP_or_30_nl
            & (NOT mux_2757_itm) & COMP_LOOP_and_277_nl & COMP_LOOP_COMP_LOOP_and_932_nl
            & COMP_LOOP_COMP_LOOP_and_934_nl & COMP_LOOP_and_1_nl & COMP_LOOP_COMP_LOOP_and_936_nl
            & COMP_LOOP_and_2_nl & COMP_LOOP_and_3_nl & COMP_LOOP_and_4_nl & COMP_LOOP_COMP_LOOP_and_930_nl
            & COMP_LOOP_and_5_nl & COMP_LOOP_and_6_nl & COMP_LOOP_and_7_nl & COMP_LOOP_and_8_nl
            & COMP_LOOP_and_9_nl & COMP_LOOP_and_10_nl & COMP_LOOP_and_11_nl & (NOT
            mux_129_nl)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_137_itm <= '0';
      ELSIF ( (and_dcpl_237 OR and_dcpl_304 OR and_dcpl_117 OR and_dcpl_130 OR and_dcpl_140
          OR and_dcpl_149 OR and_dcpl_155 OR and_dcpl_164 OR and_dcpl_171 OR and_dcpl_178
          OR and_dcpl_185 OR and_dcpl_189 OR and_dcpl_197 OR and_dcpl_202 OR and_dcpl_211
          OR and_dcpl_219 OR and_dcpl_226 OR and_dcpl_231) = '1' ) THEN
        COMP_LOOP_COMP_LOOP_and_137_itm <= MUX1HOT_s_1_3_2((NOT (z_out_1(63))), (NOT
            (z_out_6(8))), COMP_LOOP_COMP_LOOP_and_17_nl, STD_LOGIC_VECTOR'( and_dcpl_237
            & and_dcpl_304 & COMP_LOOP_or_32_cse));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (mux_3288_nl OR not_tmp_441) = '1' ) THEN
        COMP_LOOP_10_acc_8_itm <= MUX_v_64_2_2(z_out_8, STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(COMP_LOOP_1_acc_8_nl),
            64)), not_tmp_441);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (NOT((fsm_output(3)) OR (NOT (fsm_output(5))) OR (fsm_output(2)) OR or_3079_cse
          OR (NOT (fsm_output(4))) OR (fsm_output(1)) OR (NOT (fsm_output(0))) OR
          (fsm_output(9)) OR (fsm_output(10)))) = '1' ) THEN
        COMP_LOOP_acc_psp_sva <= COMP_LOOP_acc_psp_sva_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_nor_itm <= '0';
      ELSIF ( not_tmp_619 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_nor_itm <= NOT(CONV_SL_1_1(VEC_LOOP_j_sva_11_0(3 DOWNTO
            0)/=STD_LOGIC_VECTOR'("0000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_305_itm <= '0';
      ELSIF ( not_tmp_619 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_305_itm <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_62_itm <= '0';
      ELSIF ( not_tmp_619 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_62_itm <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_2_itm <= '0';
      ELSIF ( not_tmp_619 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_2_itm <= CONV_SL_1_1(VEC_LOOP_j_sva_11_0(3 DOWNTO
            0)=STD_LOGIC_VECTOR'("0011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_64_itm <= '0';
      ELSIF ( not_tmp_619 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_64_itm <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_4_itm <= '0';
      ELSIF ( not_tmp_619 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_4_itm <= CONV_SL_1_1(VEC_LOOP_j_sva_11_0(3 DOWNTO
            0)=STD_LOGIC_VECTOR'("0101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_5_itm <= '0';
      ELSIF ( not_tmp_619 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_5_itm <= CONV_SL_1_1(VEC_LOOP_j_sva_11_0(3 DOWNTO
            0)=STD_LOGIC_VECTOR'("0110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_6_itm <= '0';
      ELSIF ( not_tmp_619 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_6_itm <= CONV_SL_1_1(VEC_LOOP_j_sva_11_0(3 DOWNTO
            0)=STD_LOGIC_VECTOR'("0111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_68_itm <= '0';
      ELSIF ( not_tmp_619 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_68_itm <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1001"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_8_itm <= '0';
      ELSIF ( not_tmp_619 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_8_itm <= CONV_SL_1_1(VEC_LOOP_j_sva_11_0(3 DOWNTO
            0)=STD_LOGIC_VECTOR'("1001"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_9_itm <= '0';
      ELSIF ( not_tmp_619 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_9_itm <= CONV_SL_1_1(VEC_LOOP_j_sva_11_0(3 DOWNTO
            0)=STD_LOGIC_VECTOR'("1010"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_10_itm <= '0';
      ELSIF ( (MUX_s_1_2_2(mux_3334_nl, and_757_cse, fsm_output(8))) = '1' ) THEN
        COMP_LOOP_COMP_LOOP_and_10_itm <= MUX_s_1_2_2(COMP_LOOP_COMP_LOOP_and_10_nl,
            (NOT (COMP_LOOP_1_acc_nl(9))), and_dcpl_231);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_11_itm <= '0';
      ELSIF ( not_tmp_619 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_11_itm <= CONV_SL_1_1(VEC_LOOP_j_sva_11_0(3 DOWNTO
            0)=STD_LOGIC_VECTOR'("1100"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_12_itm <= '0';
      ELSIF ( not_tmp_619 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_12_itm <= CONV_SL_1_1(VEC_LOOP_j_sva_11_0(3 DOWNTO
            0)=STD_LOGIC_VECTOR'("1101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_13_itm <= '0';
      ELSIF ( not_tmp_619 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_13_itm <= CONV_SL_1_1(VEC_LOOP_j_sva_11_0(3 DOWNTO
            0)=STD_LOGIC_VECTOR'("1110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_14_itm <= '0';
      ELSIF ( not_tmp_619 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_14_itm <= CONV_SL_1_1(VEC_LOOP_j_sva_11_0(3 DOWNTO
            0)=STD_LOGIC_VECTOR'("1111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_1_cse_6_sva <= STD_LOGIC_VECTOR'( "000000000000");
      ELSIF ( (mux_3340_nl OR (fsm_output(10))) = '1' ) THEN
        COMP_LOOP_acc_1_cse_6_sva <= COMP_LOOP_acc_1_cse_6_sva_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_1_cse_2_sva <= STD_LOGIC_VECTOR'( "000000000000");
      ELSIF ( (mux_3350_nl OR CONV_SL_1_1(fsm_output(10 DOWNTO 8)/=STD_LOGIC_VECTOR'("000")))
          = '1' ) THEN
        COMP_LOOP_acc_1_cse_2_sva <= COMP_LOOP_acc_1_cse_2_sva_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_11_psp_sva <= STD_LOGIC_VECTOR'( "00000000000");
      ELSIF ( (NOT((NOT mux_3355_nl) AND nor_609_cse)) = '1' ) THEN
        COMP_LOOP_acc_11_psp_sva <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_sva_11_0(11
            DOWNTO 1)) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0
            & STD_LOGIC_VECTOR'( "001")), 8), 11), 11));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_1_cse_4_sva <= STD_LOGIC_VECTOR'( "000000000000");
      ELSIF ( (NOT((NOT mux_3359_nl) AND nor_609_cse)) = '1' ) THEN
        COMP_LOOP_acc_1_cse_4_sva <= z_out_6(11 DOWNTO 0);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_13_psp_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (NOT(mux_3364_nl AND (NOT (fsm_output(10))))) = '1' ) THEN
        COMP_LOOP_acc_13_psp_sva <= z_out_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_14_psp_sva <= STD_LOGIC_VECTOR'( "00000000000");
      ELSIF ( (mux_3367_nl OR (fsm_output(10))) = '1' ) THEN
        COMP_LOOP_acc_14_psp_sva <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_sva_11_0(11
            DOWNTO 1)) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0
            & STD_LOGIC_VECTOR'( "011")), 8), 11), 11));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_1_cse_8_sva <= STD_LOGIC_VECTOR'( "000000000000");
      ELSIF ( (mux_3372_nl OR (fsm_output(10))) = '1' ) THEN
        COMP_LOOP_acc_1_cse_8_sva <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_sva_11_0)
            + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0 & STD_LOGIC_VECTOR'(
            "0111")), 9), 12), 12));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_16_psp_sva <= STD_LOGIC_VECTOR'( "000000000");
      ELSIF ( (mux_3375_nl OR (fsm_output(10))) = '1' ) THEN
        COMP_LOOP_acc_16_psp_sva <= z_out_1(8 DOWNTO 0);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_1_cse_10_sva <= STD_LOGIC_VECTOR'( "000000000000");
      ELSIF ( (MUX_s_1_2_2(mux_tmp_3378, mux_3381_nl, fsm_output(5))) = '1' ) THEN
        COMP_LOOP_acc_1_cse_10_sva <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_sva_11_0)
            + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0 & STD_LOGIC_VECTOR'(
            "1001")), 9), 12), 12));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_17_psp_sva <= STD_LOGIC_VECTOR'( "00000000000");
      ELSIF ( (MUX_s_1_2_2(mux_3386_nl, (fsm_output(10)), or_470_cse)) = '1' ) THEN
        COMP_LOOP_acc_17_psp_sva <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_sva_11_0(11
            DOWNTO 1)) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0
            & STD_LOGIC_VECTOR'( "101")), 8), 11), 11));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_1_cse_12_sva <= STD_LOGIC_VECTOR'( "000000000000");
      ELSIF ( (MUX_s_1_2_2(mux_3391_nl, (fsm_output(10)), or_470_cse)) = '1' ) THEN
        COMP_LOOP_acc_1_cse_12_sva <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_sva_11_0)
            + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0 & STD_LOGIC_VECTOR'(
            "1011")), 9), 12), 12));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_19_psp_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (MUX_s_1_2_2(mux_3396_nl, (fsm_output(10)), fsm_output(9))) = '1' )
          THEN
        COMP_LOOP_acc_19_psp_sva <= z_out_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_1_cse_14_sva <= STD_LOGIC_VECTOR'( "000000000000");
      ELSIF ( (MUX_s_1_2_2(mux_3400_nl, (fsm_output(10)), fsm_output(9))) = '1' )
          THEN
        COMP_LOOP_acc_1_cse_14_sva <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_sva_11_0)
            + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0 & STD_LOGIC_VECTOR'(
            "1101")), 9), 12), 12));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_20_psp_sva <= STD_LOGIC_VECTOR'( "00000000000");
      ELSIF ( (MUX_s_1_2_2(nor_1680_nl, and_1162_nl, fsm_output(9))) = '1' ) THEN
        COMP_LOOP_acc_20_psp_sva <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_sva_11_0(11
            DOWNTO 1)) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0
            & STD_LOGIC_VECTOR'( "111")), 8), 11), 11));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_1_cse_sva <= STD_LOGIC_VECTOR'( "000000000000");
      ELSIF ( (MUX_s_1_2_2(mux_3408_nl, and_757_cse, fsm_output(8))) = '1' ) THEN
        COMP_LOOP_acc_1_cse_sva <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_sva_11_0)
            + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0 & STD_LOGIC_VECTOR'(
            "1111")), 9), 12), 12));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        modExp_exp_1_6_1_sva <= '0';
        modExp_exp_1_5_1_sva <= '0';
        modExp_exp_1_4_1_sva <= '0';
      ELSIF ( mux_3494_itm = '1' ) THEN
        modExp_exp_1_6_1_sva <= MUX1HOT_s_1_3_2((COMP_LOOP_k_9_4_sva_4_0(2)), modExp_exp_1_7_1_sva,
            (COMP_LOOP_k_9_4_sva_4_0(3)), STD_LOGIC_VECTOR'( and_dcpl_257 & not_tmp_701
            & not_tmp_688));
        modExp_exp_1_5_1_sva <= MUX1HOT_s_1_3_2((COMP_LOOP_k_9_4_sva_4_0(1)), modExp_exp_1_6_1_sva,
            (COMP_LOOP_k_9_4_sva_4_0(2)), STD_LOGIC_VECTOR'( and_dcpl_257 & not_tmp_701
            & not_tmp_688));
        modExp_exp_1_4_1_sva <= MUX1HOT_s_1_3_2((COMP_LOOP_k_9_4_sva_4_0(0)), modExp_exp_1_5_1_sva,
            (COMP_LOOP_k_9_4_sva_4_0(1)), STD_LOGIC_VECTOR'( and_dcpl_257 & not_tmp_701
            & not_tmp_688));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_10_cse_12_1_1_sva <= STD_LOGIC_VECTOR'( "000000000000");
      ELSIF ( COMP_LOOP_or_32_cse = '1' ) THEN
        COMP_LOOP_acc_10_cse_12_1_1_sva <= z_out_2_12_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (and_dcpl_117 OR not_tmp_446 OR and_dcpl_130 OR and_dcpl_149 OR and_dcpl_155
          OR and_dcpl_164 OR and_dcpl_178 OR and_dcpl_185 OR and_dcpl_189 OR and_dcpl_202
          OR and_dcpl_211 OR and_dcpl_219) = '1' ) THEN
        COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm <= MUX_s_1_2_2((z_out_3(9)), (z_out_6(8)),
            not_tmp_446);
      END IF;
    END IF;
  END PROCESS;
  modulo_result_or_nl <= and_dcpl_237 OR not_tmp_446;
  mux_2225_nl <= MUX_s_1_2_2((fsm_output(7)), and_395_cse, or_2377_cse);
  mux_2226_nl <= MUX_s_1_2_2(mux_2225_nl, mux_tmp_2172, fsm_output(9));
  nand_195_nl <= NOT(nand_196_cse AND mux_2926_cse);
  mux_2224_nl <= MUX_s_1_2_2(nand_195_nl, or_tmp_2277, fsm_output(9));
  mux_2227_nl <= MUX_s_1_2_2((NOT mux_2226_nl), mux_2224_nl, fsm_output(6));
  or_2375_nl <= CONV_SL_1_1(fsm_output(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"));
  mux_2221_nl <= MUX_s_1_2_2(or_tmp_2280, (NOT (fsm_output(7))), or_2375_nl);
  mux_2222_nl <= MUX_s_1_2_2(mux_2221_nl, or_tmp_2280, fsm_output(9));
  mux_2219_nl <= MUX_s_1_2_2(or_tmp_2276, (fsm_output(7)), and_527_cse);
  mux_2220_nl <= MUX_s_1_2_2(mux_2219_nl, or_tmp_2297, fsm_output(9));
  mux_2223_nl <= MUX_s_1_2_2(mux_2222_nl, mux_2220_nl, fsm_output(6));
  mux_2228_nl <= MUX_s_1_2_2(mux_2227_nl, mux_2223_nl, fsm_output(8));
  or_2373_nl <= (fsm_output(1)) OR (fsm_output(2)) OR (fsm_output(7)) OR (NOT (fsm_output(10)));
  or_2371_nl <= and_527_cse OR (fsm_output(7)) OR (NOT (fsm_output(10)));
  mux_2216_nl <= MUX_s_1_2_2(or_2373_nl, or_2371_nl, fsm_output(9));
  mux_2214_nl <= MUX_s_1_2_2(mux_2926_cse, or_tmp_2280, or_2368_cse);
  mux_2215_nl <= MUX_s_1_2_2((NOT (fsm_output(7))), mux_2214_nl, fsm_output(9));
  mux_2217_nl <= MUX_s_1_2_2(mux_2216_nl, mux_2215_nl, fsm_output(6));
  mux_2210_nl <= MUX_s_1_2_2((fsm_output(7)), mux_2926_cse, and_529_cse);
  mux_2211_nl <= MUX_s_1_2_2(mux_tmp_2172, mux_2210_nl, fsm_output(0));
  mux_2212_nl <= MUX_s_1_2_2(mux_2211_nl, or_tmp_2276, fsm_output(9));
  or_2367_nl <= nor_758_cse OR (NOT (fsm_output(7))) OR (fsm_output(10));
  mux_2209_nl <= MUX_s_1_2_2(or_2367_nl, or_tmp_2294, fsm_output(9));
  mux_2213_nl <= MUX_s_1_2_2(mux_2212_nl, mux_2209_nl, fsm_output(6));
  mux_2218_nl <= MUX_s_1_2_2(mux_2217_nl, mux_2213_nl, fsm_output(8));
  mux_2229_nl <= MUX_s_1_2_2(mux_2228_nl, mux_2218_nl, fsm_output(5));
  mux_2204_nl <= MUX_s_1_2_2(or_tmp_2276, (fsm_output(7)), or_2377_cse);
  mux_2205_nl <= MUX_s_1_2_2((fsm_output(7)), mux_2204_nl, fsm_output(9));
  mux_2206_nl <= MUX_s_1_2_2(mux_2205_nl, mux_2203_cse, fsm_output(6));
  or_2364_nl <= (fsm_output(1)) OR (fsm_output(2)) OR (NOT (fsm_output(7))) OR (fsm_output(10));
  mux_2200_nl <= MUX_s_1_2_2(or_2364_nl, or_tmp_2274, fsm_output(0));
  mux_2201_nl <= MUX_s_1_2_2(mux_tmp_2178, mux_2200_nl, fsm_output(9));
  mux_2197_nl <= MUX_s_1_2_2((fsm_output(7)), or_tmp_2281, or_2368_cse);
  or_2362_nl <= and_529_cse OR (fsm_output(7)) OR (NOT (fsm_output(10)));
  mux_2198_nl <= MUX_s_1_2_2(mux_2197_nl, or_2362_nl, fsm_output(0));
  or_2360_nl <= (fsm_output(2)) OR (fsm_output(7)) OR (fsm_output(10));
  mux_2199_nl <= MUX_s_1_2_2(mux_2198_nl, or_2360_nl, fsm_output(9));
  mux_2202_nl <= MUX_s_1_2_2(mux_2201_nl, mux_2199_nl, fsm_output(6));
  mux_2207_nl <= MUX_s_1_2_2(mux_2206_nl, mux_2202_nl, fsm_output(8));
  mux_2192_nl <= MUX_s_1_2_2((NOT or_tmp_2280), or_tmp_2281, fsm_output(2));
  mux_2191_nl <= MUX_s_1_2_2((fsm_output(7)), or_tmp_2281, fsm_output(2));
  mux_2193_nl <= MUX_s_1_2_2(mux_2192_nl, mux_2191_nl, and_526_cse);
  mux_2194_nl <= MUX_s_1_2_2((NOT mux_2193_nl), or_tmp_2280, fsm_output(9));
  mux_2190_nl <= MUX_s_1_2_2(mux_tmp_2176, or_tmp_2302, fsm_output(9));
  mux_2195_nl <= MUX_s_1_2_2(mux_2194_nl, mux_2190_nl, fsm_output(6));
  mux_2187_nl <= MUX_s_1_2_2((fsm_output(7)), and_395_cse, and_527_cse);
  mux_2188_nl <= MUX_s_1_2_2((NOT mux_2187_nl), or_tmp_2280, fsm_output(9));
  mux_2189_nl <= MUX_s_1_2_2(mux_tmp_2159, mux_2188_nl, fsm_output(6));
  mux_2196_nl <= MUX_s_1_2_2(mux_2195_nl, mux_2189_nl, fsm_output(8));
  mux_2208_nl <= MUX_s_1_2_2(mux_2207_nl, mux_2196_nl, fsm_output(5));
  mux_2230_nl <= MUX_s_1_2_2(mux_2229_nl, mux_2208_nl, fsm_output(4));
  mux_2180_nl <= MUX_s_1_2_2(mux_tmp_2178, or_tmp_2302, fsm_output(1));
  mux_2181_nl <= MUX_s_1_2_2(mux_2180_nl, or_tmp_2297, fsm_output(0));
  or_2357_nl <= (fsm_output(2)) OR (NOT and_395_cse);
  mux_2179_nl <= MUX_s_1_2_2(or_2357_nl, mux_tmp_2178, or_3388_cse);
  mux_2182_nl <= MUX_s_1_2_2(mux_2181_nl, mux_2179_nl, fsm_output(9));
  or_2355_nl <= (NOT (fsm_output(2))) OR (fsm_output(7)) OR (NOT (fsm_output(10)));
  mux_2177_nl <= MUX_s_1_2_2(or_2355_nl, mux_tmp_2176, fsm_output(9));
  mux_2183_nl <= MUX_s_1_2_2(mux_2182_nl, mux_2177_nl, fsm_output(6));
  mux_2173_nl <= MUX_s_1_2_2((NOT mux_tmp_2172), or_tmp_2280, fsm_output(9));
  mux_2174_nl <= MUX_s_1_2_2(mux_2173_nl, mux_2171_cse, fsm_output(6));
  mux_2184_nl <= MUX_s_1_2_2(mux_2183_nl, mux_2174_nl, fsm_output(8));
  or_2351_nl <= (fsm_output(9)) OR or_tmp_2294;
  mux_2167_nl <= MUX_s_1_2_2((fsm_output(7)), and_395_cse, or_2368_cse);
  or_2347_nl <= and_527_cse OR (NOT (fsm_output(7))) OR (fsm_output(10));
  mux_2168_nl <= MUX_s_1_2_2((NOT mux_2167_nl), or_2347_nl, fsm_output(9));
  mux_2169_nl <= MUX_s_1_2_2(or_2351_nl, mux_2168_nl, fsm_output(6));
  mux_2163_nl <= MUX_s_1_2_2((NOT mux_2926_cse), or_tmp_2276, fsm_output(2));
  mux_2162_nl <= MUX_s_1_2_2((NOT mux_2926_cse), (fsm_output(7)), fsm_output(2));
  mux_2164_nl <= MUX_s_1_2_2(mux_2163_nl, mux_2162_nl, or_3388_cse);
  mux_2160_nl <= MUX_s_1_2_2(or_tmp_2276, or_tmp_2280, or_2368_cse);
  or_2343_nl <= (NOT(nor_758_cse OR (fsm_output(7)))) OR (fsm_output(10));
  mux_2161_nl <= MUX_s_1_2_2(mux_2160_nl, or_2343_nl, fsm_output(0));
  mux_2165_nl <= MUX_s_1_2_2((NOT mux_2164_nl), mux_2161_nl, fsm_output(9));
  mux_2166_nl <= MUX_s_1_2_2(mux_2165_nl, mux_tmp_2159, fsm_output(6));
  mux_2170_nl <= MUX_s_1_2_2(mux_2169_nl, mux_2166_nl, fsm_output(8));
  mux_2185_nl <= MUX_s_1_2_2(mux_2184_nl, mux_2170_nl, fsm_output(5));
  mux_2154_nl <= MUX_s_1_2_2((fsm_output(7)), or_tmp_2281, and_527_cse);
  mux_2153_nl <= MUX_s_1_2_2((fsm_output(7)), or_tmp_2281, and_536_cse);
  mux_2155_nl <= MUX_s_1_2_2(mux_2154_nl, mux_2153_nl, fsm_output(9));
  mux_2150_nl <= MUX_s_1_2_2((NOT mux_2926_cse), or_tmp_2276, and_529_cse);
  mux_2149_nl <= MUX_s_1_2_2((NOT mux_2926_cse), (fsm_output(7)), and_529_cse);
  mux_2151_nl <= MUX_s_1_2_2(mux_2150_nl, mux_2149_nl, fsm_output(0));
  mux_2147_nl <= MUX_s_1_2_2((fsm_output(7)), mux_2926_cse, fsm_output(2));
  mux_2146_nl <= MUX_s_1_2_2(and_395_cse, mux_2926_cse, fsm_output(2));
  mux_2148_nl <= MUX_s_1_2_2(mux_2147_nl, mux_2146_nl, and_526_cse);
  mux_2152_nl <= MUX_s_1_2_2((NOT mux_2151_nl), mux_2148_nl, fsm_output(9));
  mux_2156_nl <= MUX_s_1_2_2(mux_2155_nl, mux_2152_nl, fsm_output(6));
  mux_2143_nl <= MUX_s_1_2_2(or_tmp_2276, (fsm_output(7)), or_2368_cse);
  mux_2144_nl <= MUX_s_1_2_2(mux_2143_nl, or_tmp_2276, fsm_output(9));
  or_2339_nl <= (fsm_output(6)) OR mux_2144_nl;
  mux_2157_nl <= MUX_s_1_2_2(mux_2156_nl, or_2339_nl, fsm_output(8));
  mux_2140_nl <= MUX_s_1_2_2((NOT or_tmp_2281), or_tmp_2280, fsm_output(9));
  or_2335_nl <= (NOT (fsm_output(9))) OR (fsm_output(1)) OR (fsm_output(2));
  mux_2139_nl <= MUX_s_1_2_2(or_tmp_2276, (fsm_output(7)), or_2335_nl);
  mux_2141_nl <= MUX_s_1_2_2(mux_2140_nl, mux_2139_nl, fsm_output(6));
  nand_197_nl <= NOT(nand_196_cse AND and_395_cse);
  mux_2135_nl <= MUX_s_1_2_2((NOT and_395_cse), or_tmp_2276, and_529_cse);
  mux_2136_nl <= MUX_s_1_2_2(nand_197_nl, mux_2135_nl, fsm_output(0));
  mux_2137_nl <= MUX_s_1_2_2(mux_2136_nl, or_tmp_2277, fsm_output(9));
  mux_2133_nl <= MUX_s_1_2_2((NOT and_395_cse), or_tmp_2276, or_2377_cse);
  mux_2134_nl <= MUX_s_1_2_2(mux_2133_nl, or_tmp_2274, fsm_output(9));
  mux_2138_nl <= MUX_s_1_2_2(mux_2137_nl, mux_2134_nl, fsm_output(6));
  mux_2142_nl <= MUX_s_1_2_2(mux_2141_nl, mux_2138_nl, fsm_output(8));
  mux_2158_nl <= MUX_s_1_2_2(mux_2157_nl, mux_2142_nl, fsm_output(5));
  mux_2186_nl <= MUX_s_1_2_2(mux_2185_nl, mux_2158_nl, fsm_output(4));
  mux_2231_nl <= MUX_s_1_2_2(mux_2230_nl, mux_2186_nl, fsm_output(3));
  mux_2324_nl <= MUX_s_1_2_2(or_3008_cse, or_259_cse, fsm_output(1));
  mux_2325_nl <= MUX_s_1_2_2(mux_2324_nl, mux_tmp_2311, fsm_output(0));
  mux_2326_nl <= MUX_s_1_2_2(mux_2325_nl, mux_tmp_130, fsm_output(3));
  and_519_nl <= or_3388_cse AND (fsm_output(9));
  mux_2322_nl <= MUX_s_1_2_2((fsm_output(8)), or_tmp_93, and_519_nl);
  mux_2323_nl <= MUX_s_1_2_2(mux_3555_cse, mux_2322_nl, fsm_output(3));
  mux_2327_nl <= MUX_s_1_2_2(mux_2326_nl, mux_2323_nl, fsm_output(6));
  mux_2319_nl <= MUX_s_1_2_2(or_tmp_2360, or_tmp_2341, fsm_output(0));
  mux_2318_nl <= MUX_s_1_2_2((fsm_output(8)), or_tmp_94, or_2421_cse);
  mux_2320_nl <= MUX_s_1_2_2(mux_2319_nl, mux_2318_nl, fsm_output(3));
  mux_2321_nl <= MUX_s_1_2_2(mux_2320_nl, mux_tmp_2287, fsm_output(6));
  mux_2328_nl <= MUX_s_1_2_2(mux_2327_nl, mux_2321_nl, fsm_output(7));
  mux_2314_nl <= MUX_s_1_2_2((fsm_output(8)), or_tmp_94, or_2419_cse);
  mux_2315_nl <= MUX_s_1_2_2(mux_2314_nl, (fsm_output(8)), fsm_output(3));
  mux_2312_nl <= MUX_s_1_2_2(mux_tmp_2311, mux_tmp_2293, fsm_output(0));
  mux_2313_nl <= MUX_s_1_2_2(mux_tmp_130, mux_2312_nl, fsm_output(3));
  mux_2316_nl <= MUX_s_1_2_2(mux_2315_nl, mux_2313_nl, fsm_output(6));
  or_2418_nl <= (NOT((fsm_output(3)) OR (fsm_output(0)) OR (fsm_output(1)))) OR (fsm_output(9));
  mux_2309_nl <= MUX_s_1_2_2((fsm_output(8)), or_tmp_94, or_2418_nl);
  mux_2307_nl <= MUX_s_1_2_2(mux_tmp_130, mux_tmp_141, fsm_output(1));
  mux_2308_nl <= MUX_s_1_2_2(mux_2307_nl, or_tmp_2341, fsm_output(3));
  mux_2310_nl <= MUX_s_1_2_2(mux_2309_nl, mux_2308_nl, fsm_output(6));
  mux_2317_nl <= MUX_s_1_2_2(mux_2316_nl, mux_2310_nl, fsm_output(7));
  mux_2329_nl <= MUX_s_1_2_2(mux_2328_nl, mux_2317_nl, fsm_output(5));
  mux_2303_nl <= MUX_s_1_2_2(mux_tmp_130, or_tmp_2360, fsm_output(3));
  mux_2301_nl <= MUX_s_1_2_2(or_2998_cse, or_2414_cse, or_3388_cse);
  mux_2300_nl <= MUX_s_1_2_2(mux_1036_cse, mux_tmp_130, or_3388_cse);
  mux_2302_nl <= MUX_s_1_2_2(mux_2301_nl, mux_2300_nl, fsm_output(3));
  mux_2304_nl <= MUX_s_1_2_2(mux_2303_nl, mux_2302_nl, fsm_output(6));
  mux_2296_nl <= MUX_s_1_2_2((fsm_output(8)), or_tmp_93, or_2419_cse);
  mux_2297_nl <= MUX_s_1_2_2(mux_tmp_2289, mux_2296_nl, fsm_output(0));
  mux_2298_nl <= MUX_s_1_2_2((fsm_output(8)), mux_2297_nl, fsm_output(3));
  or_2408_nl <= nor_303_cse OR (NOT (fsm_output(8))) OR (fsm_output(10));
  mux_2294_nl <= MUX_s_1_2_2(mux_tmp_2293, or_2408_nl, fsm_output(0));
  mux_2295_nl <= MUX_s_1_2_2(mux_2294_nl, mux_tmp_130, fsm_output(3));
  mux_2299_nl <= MUX_s_1_2_2(mux_2298_nl, mux_2295_nl, fsm_output(6));
  mux_2305_nl <= MUX_s_1_2_2(mux_2304_nl, mux_2299_nl, fsm_output(7));
  mux_2288_nl <= MUX_s_1_2_2(or_2407_cse, mux_tmp_165, fsm_output(1));
  mux_2290_nl <= MUX_s_1_2_2(mux_tmp_2289, mux_2288_nl, fsm_output(3));
  mux_2291_nl <= MUX_s_1_2_2(mux_2290_nl, mux_tmp_2287, fsm_output(6));
  or_2406_nl <= and_526_cse OR CONV_SL_1_1(fsm_output(10 DOWNTO 8)/=STD_LOGIC_VECTOR'("100"));
  or_2404_nl <= and_521_cse OR (NOT (fsm_output(8))) OR (fsm_output(10));
  mux_2285_nl <= MUX_s_1_2_2(or_2406_nl, or_2404_nl, fsm_output(3));
  mux_2286_nl <= MUX_s_1_2_2(mux_2285_nl, mux_tmp_139, fsm_output(6));
  mux_2292_nl <= MUX_s_1_2_2(mux_2291_nl, mux_2286_nl, fsm_output(7));
  mux_2306_nl <= MUX_s_1_2_2(mux_2305_nl, mux_2292_nl, fsm_output(5));
  mux_2330_nl <= MUX_s_1_2_2(mux_2329_nl, mux_2306_nl, fsm_output(4));
  or_2403_nl <= nor_297_cse OR (NOT (fsm_output(8))) OR (fsm_output(10));
  mux_2280_nl <= MUX_s_1_2_2(or_2403_nl, mux_tmp_130, fsm_output(3));
  or_2402_nl <= (fsm_output(1)) OR (fsm_output(9));
  mux_2278_nl <= MUX_s_1_2_2(or_tmp_93, (fsm_output(8)), or_2402_nl);
  mux_2277_nl <= MUX_s_1_2_2(mux_981_cse, or_2998_cse, and_526_cse);
  mux_2279_nl <= MUX_s_1_2_2(mux_2278_nl, mux_2277_nl, fsm_output(3));
  mux_2281_nl <= MUX_s_1_2_2(mux_2280_nl, mux_2279_nl, fsm_output(6));
  mux_2275_nl <= MUX_s_1_2_2(or_tmp_2340, (fsm_output(8)), fsm_output(3));
  mux_2276_nl <= MUX_s_1_2_2(mux_2275_nl, mux_tmp_2241, fsm_output(6));
  mux_2282_nl <= MUX_s_1_2_2(mux_2281_nl, mux_2276_nl, fsm_output(7));
  nor_295_nl <= NOT((fsm_output(3)) OR (fsm_output(0)) OR (fsm_output(1)) OR (NOT
      (fsm_output(9))));
  mux_2272_nl <= MUX_s_1_2_2((fsm_output(8)), or_tmp_94, nor_295_nl);
  mux_2270_nl <= MUX_s_1_2_2((NOT (fsm_output(8))), or_tmp_88, or_2400_cse);
  mux_2271_nl <= MUX_s_1_2_2(mux_tmp_2262, mux_2270_nl, fsm_output(3));
  mux_2273_nl <= MUX_s_1_2_2(mux_2272_nl, mux_2271_nl, fsm_output(6));
  mux_2267_nl <= MUX_s_1_2_2(mux_tmp_141, or_3008_cse, or_3388_cse);
  or_2398_nl <= nor_297_cse OR (fsm_output(8)) OR (fsm_output(10));
  mux_2268_nl <= MUX_s_1_2_2(mux_2267_nl, or_2398_nl, fsm_output(3));
  mux_2269_nl <= MUX_s_1_2_2(mux_tmp_2235, mux_2268_nl, fsm_output(6));
  mux_2274_nl <= MUX_s_1_2_2(mux_2273_nl, mux_2269_nl, fsm_output(7));
  mux_2283_nl <= MUX_s_1_2_2(mux_2282_nl, mux_2274_nl, fsm_output(5));
  mux_2261_nl <= MUX_s_1_2_2(or_tmp_2341, or_tmp_2340, fsm_output(0));
  mux_2263_nl <= MUX_s_1_2_2(mux_tmp_2262, mux_2261_nl, fsm_output(3));
  or_2395_nl <= (NOT(CONV_SL_1_1(fsm_output(9 DOWNTO 8)/=STD_LOGIC_VECTOR'("10"))))
      OR (fsm_output(10));
  mux_2259_nl <= MUX_s_1_2_2(or_2395_nl, mux_1036_cse, and_526_cse);
  mux_2260_nl <= MUX_s_1_2_2(mux_2259_nl, mux_tmp_130, fsm_output(3));
  mux_2264_nl <= MUX_s_1_2_2(mux_2263_nl, mux_2260_nl, fsm_output(6));
  mux_2255_nl <= MUX_s_1_2_2(or_tmp_93, (fsm_output(8)), or_2419_cse);
  mux_2251_nl <= MUX_s_1_2_2(or_tmp_94, (fsm_output(8)), fsm_output(9));
  mux_2253_nl <= MUX_s_1_2_2(mux_981_cse, mux_2251_nl, fsm_output(1));
  mux_2250_nl <= MUX_s_1_2_2(or_tmp_94, or_tmp_93, nor_303_cse);
  mux_2254_nl <= MUX_s_1_2_2(mux_2253_nl, mux_2250_nl, fsm_output(0));
  mux_2256_nl <= MUX_s_1_2_2(mux_2255_nl, mux_2254_nl, fsm_output(3));
  or_2392_nl <= (NOT((fsm_output(3)) OR (fsm_output(1)))) OR (fsm_output(9));
  mux_2249_nl <= MUX_s_1_2_2((NOT (fsm_output(8))), or_tmp_88, or_2392_nl);
  mux_2257_nl <= MUX_s_1_2_2(mux_2256_nl, mux_2249_nl, fsm_output(6));
  mux_2265_nl <= MUX_s_1_2_2(mux_2264_nl, mux_2257_nl, fsm_output(7));
  or_2390_nl <= (NOT((NOT (fsm_output(1))) OR (fsm_output(9)))) OR (fsm_output(8))
      OR (NOT (fsm_output(10)));
  or_2385_nl <= CONV_SL_1_1(fsm_output(9 DOWNTO 8)/=STD_LOGIC_VECTOR'("10"));
  mux_2244_nl <= MUX_s_1_2_2(or_2387_cse, or_2385_nl, fsm_output(1));
  mux_2245_nl <= MUX_s_1_2_2(or_2390_nl, mux_2244_nl, fsm_output(0));
  mux_2243_nl <= MUX_s_1_2_2(mux_tmp_165, mux_3555_cse, or_3388_cse);
  mux_2246_nl <= MUX_s_1_2_2(mux_2245_nl, mux_2243_nl, fsm_output(3));
  mux_2247_nl <= MUX_s_1_2_2(mux_2246_nl, mux_tmp_2241, fsm_output(6));
  mux_2236_nl <= MUX_s_1_2_2((fsm_output(8)), (NOT or_tmp_88), or_2419_cse);
  nand_51_nl <= NOT((fsm_output(3)) AND mux_2236_nl);
  mux_2237_nl <= MUX_s_1_2_2(nand_51_nl, mux_tmp_2235, fsm_output(6));
  mux_2248_nl <= MUX_s_1_2_2(mux_2247_nl, mux_2237_nl, fsm_output(7));
  mux_2266_nl <= MUX_s_1_2_2(mux_2265_nl, mux_2248_nl, fsm_output(5));
  mux_2284_nl <= MUX_s_1_2_2(mux_2283_nl, mux_2266_nl, fsm_output(4));
  mux_2331_nl <= MUX_s_1_2_2(mux_2330_nl, mux_2284_nl, fsm_output(2));
  and_517_nl <= (fsm_output(4)) AND mux_125_cse;
  nor_752_nl <= NOT((fsm_output(4)) OR (fsm_output(7)) OR mux_tmp_119);
  mux_2343_nl <= MUX_s_1_2_2(and_517_nl, nor_752_nl, fsm_output(1));
  nand_189_nl <= NOT((fsm_output(5)) AND mux_2343_nl);
  or_3386_nl <= (fsm_output(1)) OR (NOT (fsm_output(4))) OR (fsm_output(7)) OR (NOT
      (fsm_output(3))) OR (fsm_output(8)) OR (NOT (fsm_output(6))) OR (fsm_output(10));
  nand_190_nl <= NOT((fsm_output(1)) AND (fsm_output(4)) AND (fsm_output(7)) AND
      (fsm_output(3)) AND (fsm_output(8)) AND (fsm_output(6)) AND (fsm_output(10)));
  mux_2341_nl <= MUX_s_1_2_2(or_3386_nl, nand_190_nl, fsm_output(5));
  mux_2344_nl <= MUX_s_1_2_2(nand_189_nl, mux_2341_nl, fsm_output(2));
  or_2437_nl <= (NOT (fsm_output(4))) OR (NOT (fsm_output(7))) OR (fsm_output(3))
      OR (NOT (fsm_output(8))) OR (fsm_output(6)) OR (fsm_output(10));
  mux_2340_nl <= MUX_s_1_2_2(or_2437_nl, or_tmp_2376, fsm_output(1));
  or_2438_nl <= (NOT (fsm_output(2))) OR (fsm_output(5)) OR mux_2340_nl;
  mux_2345_nl <= MUX_s_1_2_2(mux_2344_nl, or_2438_nl, fsm_output(9));
  or_2435_nl <= (NOT (fsm_output(7))) OR (NOT (fsm_output(3))) OR (fsm_output(8))
      OR not_tmp_49;
  or_2433_nl <= (NOT (fsm_output(7))) OR (fsm_output(3)) OR (NOT (fsm_output(8)))
      OR (fsm_output(6)) OR (fsm_output(10));
  mux_2335_nl <= MUX_s_1_2_2(or_2435_nl, or_2433_nl, fsm_output(4));
  mux_2336_nl <= MUX_s_1_2_2(mux_2335_nl, or_tmp_2376, fsm_output(1));
  or_2431_nl <= (NOT (fsm_output(1))) OR (NOT (fsm_output(4))) OR (fsm_output(7))
      OR (fsm_output(3)) OR (fsm_output(8)) OR (fsm_output(6)) OR (fsm_output(10));
  mux_2337_nl <= MUX_s_1_2_2(mux_2336_nl, or_2431_nl, fsm_output(5));
  or_2430_nl <= (fsm_output(5)) OR (NOT (fsm_output(1))) OR (NOT (fsm_output(4)))
      OR (NOT (fsm_output(7))) OR (fsm_output(3)) OR (NOT (fsm_output(8))) OR (fsm_output(6))
      OR (NOT (fsm_output(10)));
  mux_2338_nl <= MUX_s_1_2_2(mux_2337_nl, or_2430_nl, fsm_output(2));
  nand_191_nl <= NOT((fsm_output(5)) AND (fsm_output(1)) AND (fsm_output(4)) AND
      (fsm_output(7)) AND (fsm_output(3)) AND (fsm_output(8)) AND (fsm_output(6))
      AND (NOT (fsm_output(10))));
  or_2427_nl <= (NOT (fsm_output(1))) OR (NOT (fsm_output(4))) OR (fsm_output(7))
      OR (NOT (fsm_output(3))) OR (fsm_output(8)) OR (NOT (fsm_output(6))) OR (fsm_output(10));
  or_2426_nl <= (fsm_output(1)) OR (fsm_output(4)) OR (fsm_output(7)) OR mux_tmp_119;
  mux_2333_nl <= MUX_s_1_2_2(or_2427_nl, or_2426_nl, fsm_output(5));
  mux_2334_nl <= MUX_s_1_2_2(nand_191_nl, mux_2333_nl, fsm_output(2));
  mux_2339_nl <= MUX_s_1_2_2(mux_2338_nl, mux_2334_nl, fsm_output(9));
  mux_2346_nl <= MUX_s_1_2_2(mux_2345_nl, mux_2339_nl, fsm_output(0));
  mux_2414_nl <= MUX_s_1_2_2(mux_tmp_2389, or_tmp_2396, fsm_output(7));
  mux_2413_nl <= MUX_s_1_2_2(mux_tmp_2386, mux_tmp_2353, fsm_output(7));
  mux_2415_nl <= MUX_s_1_2_2(mux_2414_nl, mux_2413_nl, fsm_output(2));
  mux_2411_nl <= MUX_s_1_2_2(mux_tmp_2378, mux_tmp_2382, fsm_output(7));
  mux_2410_nl <= MUX_s_1_2_2(mux_tmp_2376, nand_tmp_54, fsm_output(7));
  mux_2412_nl <= MUX_s_1_2_2(mux_2411_nl, mux_2410_nl, fsm_output(2));
  mux_2416_nl <= MUX_s_1_2_2(mux_2415_nl, mux_2412_nl, fsm_output(3));
  mux_2405_nl <= MUX_s_1_2_2(mux_tmp_2347, mux_tmp_2369, fsm_output(6));
  mux_2406_nl <= MUX_s_1_2_2(mux_tmp_2371, mux_2405_nl, fsm_output(0));
  mux_2407_nl <= MUX_s_1_2_2(mux_2406_nl, nand_tmp_54, fsm_output(7));
  mux_2403_nl <= MUX_s_1_2_2(mux_tmp_2365, mux_tmp_2361, fsm_output(0));
  mux_2401_nl <= MUX_s_1_2_2(or_tmp_2390, mux_tmp_2363, fsm_output(6));
  mux_2402_nl <= MUX_s_1_2_2(mux_tmp_2364, mux_2401_nl, fsm_output(0));
  mux_2404_nl <= MUX_s_1_2_2(mux_2403_nl, mux_2402_nl, fsm_output(7));
  mux_2408_nl <= MUX_s_1_2_2(mux_2407_nl, mux_2404_nl, fsm_output(2));
  mux_2397_nl <= MUX_s_1_2_2(mux_tmp_2348, mux_tmp_2359, fsm_output(6));
  mux_2398_nl <= MUX_s_1_2_2(mux_2397_nl, mux_tmp_2356, fsm_output(0));
  mux_2399_nl <= MUX_s_1_2_2(or_tmp_2396, mux_2398_nl, fsm_output(7));
  mux_2395_nl <= MUX_s_1_2_2(or_tmp_2396, mux_tmp_2353, fsm_output(0));
  mux_2396_nl <= MUX_s_1_2_2(mux_2395_nl, mux_tmp_2350, fsm_output(7));
  mux_2400_nl <= MUX_s_1_2_2(mux_2399_nl, mux_2396_nl, fsm_output(2));
  mux_2409_nl <= MUX_s_1_2_2(mux_2408_nl, mux_2400_nl, fsm_output(3));
  mux_2417_nl <= MUX_s_1_2_2(mux_2416_nl, mux_2409_nl, fsm_output(4));
  mux_2390_nl <= MUX_s_1_2_2(mux_tmp_2389, mux_tmp_2386, fsm_output(0));
  mux_2391_nl <= MUX_s_1_2_2(mux_2390_nl, or_tmp_2396, fsm_output(7));
  mux_2383_nl <= MUX_s_1_2_2(mux_tmp_2353, mux_tmp_2382, fsm_output(0));
  mux_2384_nl <= MUX_s_1_2_2(mux_tmp_2378, mux_2383_nl, fsm_output(7));
  mux_2392_nl <= MUX_s_1_2_2(mux_2391_nl, mux_2384_nl, fsm_output(2));
  mux_2379_nl <= MUX_s_1_2_2(mux_tmp_2378, mux_tmp_2376, fsm_output(0));
  mux_2380_nl <= MUX_s_1_2_2(mux_2379_nl, nand_tmp_54, fsm_output(7));
  mux_2372_nl <= MUX_s_1_2_2(mux_tmp_2370, or_tmp_2405, fsm_output(6));
  mux_2373_nl <= MUX_s_1_2_2(mux_2372_nl, mux_tmp_2371, fsm_output(0));
  mux_2374_nl <= MUX_s_1_2_2(mux_2373_nl, nand_tmp_54, fsm_output(7));
  mux_2381_nl <= MUX_s_1_2_2(mux_2380_nl, mux_2374_nl, fsm_output(2));
  mux_2393_nl <= MUX_s_1_2_2(mux_2392_nl, mux_2381_nl, fsm_output(3));
  mux_2366_nl <= MUX_s_1_2_2(mux_tmp_2365, mux_tmp_2364, fsm_output(7));
  mux_2360_nl <= MUX_s_1_2_2(or_tmp_2390, mux_tmp_2359, fsm_output(6));
  mux_2362_nl <= MUX_s_1_2_2(mux_tmp_2361, mux_2360_nl, fsm_output(7));
  mux_2367_nl <= MUX_s_1_2_2(mux_2366_nl, mux_2362_nl, fsm_output(2));
  mux_2357_nl <= MUX_s_1_2_2(or_tmp_2396, mux_tmp_2356, fsm_output(7));
  mux_2349_nl <= MUX_s_1_2_2(mux_tmp_2348, mux_tmp_2347, fsm_output(6));
  mux_2351_nl <= MUX_s_1_2_2(mux_tmp_2350, mux_2349_nl, fsm_output(0));
  mux_2354_nl <= MUX_s_1_2_2(mux_tmp_2353, mux_2351_nl, fsm_output(7));
  mux_2358_nl <= MUX_s_1_2_2(mux_2357_nl, mux_2354_nl, fsm_output(2));
  mux_2368_nl <= MUX_s_1_2_2(mux_2367_nl, mux_2358_nl, fsm_output(3));
  mux_2394_nl <= MUX_s_1_2_2(mux_2393_nl, mux_2368_nl, fsm_output(4));
  mux_2418_nl <= MUX_s_1_2_2(mux_2417_nl, mux_2394_nl, fsm_output(1));
  COMP_LOOP_nor_11_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("000")));
  COMP_LOOP_and_274_nl <= (NOT and_dcpl_256) AND and_dcpl_247;
  or_2881_nl <= nor_653_cse OR (NOT (fsm_output(8))) OR (fsm_output(10));
  mux_3065_nl <= MUX_s_1_2_2(or_2881_nl, mux_tmp_3049, fsm_output(1));
  mux_3066_nl <= MUX_s_1_2_2(mux_3065_nl, mux_1036_cse, fsm_output(4));
  mux_3063_nl <= MUX_s_1_2_2(mux_tmp_3024, or_tmp_2802, or_3388_cse);
  mux_3064_nl <= MUX_s_1_2_2(mux_tmp_130, mux_3063_nl, fsm_output(4));
  mux_3067_nl <= MUX_s_1_2_2(mux_3066_nl, mux_3064_nl, fsm_output(7));
  mux_3060_nl <= MUX_s_1_2_2(mux_tmp_130, mux_tmp_3032, and_526_cse);
  or_449_nl <= (NOT (fsm_output(2))) OR (fsm_output(9)) OR (fsm_output(8)) OR (fsm_output(10));
  or_2876_nl <= nor_653_cse OR (fsm_output(8)) OR (fsm_output(10));
  mux_3059_nl <= MUX_s_1_2_2(or_449_nl, or_2876_nl, fsm_output(1));
  mux_3061_nl <= MUX_s_1_2_2(mux_3060_nl, mux_3059_nl, fsm_output(4));
  mux_3062_nl <= MUX_s_1_2_2(mux_3061_nl, mux_tmp_139, fsm_output(7));
  mux_3068_nl <= MUX_s_1_2_2(mux_3067_nl, mux_3062_nl, fsm_output(5));
  nor_407_nl <= NOT((fsm_output(4)) OR (NOT (fsm_output(1))) OR (fsm_output(0)) OR
      (fsm_output(9)) OR (NOT (fsm_output(2))));
  mux_3056_nl <= MUX_s_1_2_2((fsm_output(8)), or_tmp_93, nor_407_nl);
  mux_3053_nl <= MUX_s_1_2_2(or_tmp_93, or_tmp_2814, fsm_output(9));
  mux_3051_nl <= MUX_s_1_2_2(or_tmp_2795, or_tmp_2814, fsm_output(9));
  or_439_nl <= (fsm_output(2)) OR (fsm_output(9)) OR (fsm_output(8)) OR (NOT (fsm_output(10)));
  mux_3052_nl <= MUX_s_1_2_2(mux_3051_nl, or_439_nl, fsm_output(0));
  mux_3054_nl <= MUX_s_1_2_2(mux_3053_nl, mux_3052_nl, fsm_output(1));
  mux_3050_nl <= MUX_s_1_2_2(mux_tmp_3049, mux_tmp_3007, fsm_output(1));
  mux_3055_nl <= MUX_s_1_2_2(mux_3054_nl, mux_3050_nl, fsm_output(4));
  mux_3057_nl <= MUX_s_1_2_2(mux_3056_nl, mux_3055_nl, fsm_output(7));
  or_2870_nl <= (fsm_output(1)) OR (NOT (fsm_output(9))) OR (fsm_output(2)) OR (fsm_output(8))
      OR (NOT (fsm_output(10)));
  mux_3047_nl <= MUX_s_1_2_2(or_2870_nl, mux_tmp_130, fsm_output(4));
  mux_3045_nl <= MUX_s_1_2_2(mux_tmp_130, mux_tmp_3032, or_3388_cse);
  mux_3046_nl <= MUX_s_1_2_2(mux_tmp_130, mux_3045_nl, fsm_output(4));
  mux_3048_nl <= MUX_s_1_2_2(mux_3047_nl, mux_3046_nl, fsm_output(7));
  mux_3058_nl <= MUX_s_1_2_2(mux_3057_nl, mux_3048_nl, fsm_output(5));
  mux_3069_nl <= MUX_s_1_2_2(mux_3068_nl, mux_3058_nl, fsm_output(6));
  mux_3039_nl <= MUX_s_1_2_2((NOT mux_tmp_3014), or_tmp_88, fsm_output(9));
  mux_3040_nl <= MUX_s_1_2_2(mux_3039_nl, mux_1036_cse, fsm_output(1));
  mux_3035_nl <= MUX_s_1_2_2(or_tmp_93, (fsm_output(8)), fsm_output(2));
  mux_3036_nl <= MUX_s_1_2_2((NOT mux_3035_nl), or_tmp_88, fsm_output(9));
  mux_3038_nl <= MUX_s_1_2_2(mux_1036_cse, mux_3036_nl, or_3388_cse);
  mux_3041_nl <= MUX_s_1_2_2(mux_3040_nl, mux_3038_nl, fsm_output(4));
  mux_3033_nl <= MUX_s_1_2_2(mux_tmp_130, mux_tmp_3032, fsm_output(1));
  or_2866_nl <= (NOT((fsm_output(0)) OR (NOT (fsm_output(9))))) OR (NOT (fsm_output(2)))
      OR (fsm_output(8)) OR (fsm_output(10));
  or_2865_nl <= nor_657_cse OR (fsm_output(8)) OR (fsm_output(10));
  mux_3030_nl <= MUX_s_1_2_2(or_2866_nl, or_2865_nl, fsm_output(1));
  mux_3034_nl <= MUX_s_1_2_2(mux_3033_nl, mux_3030_nl, fsm_output(4));
  mux_3042_nl <= MUX_s_1_2_2(mux_3041_nl, mux_3034_nl, fsm_output(7));
  mux_3025_nl <= MUX_s_1_2_2((NOT nor_tmp_405), or_tmp_2803, fsm_output(9));
  mux_3026_nl <= MUX_s_1_2_2(mux_3025_nl, mux_tmp_3024, fsm_output(0));
  mux_3027_nl <= MUX_s_1_2_2(mux_3026_nl, or_tmp_2802, fsm_output(1));
  or_2859_nl <= (NOT(nor_753_cse OR (fsm_output(9)))) OR (fsm_output(2));
  mux_3023_nl <= MUX_s_1_2_2(or_tmp_94, (fsm_output(8)), or_2859_nl);
  mux_3028_nl <= MUX_s_1_2_2(mux_3027_nl, mux_3023_nl, fsm_output(4));
  mux_3029_nl <= MUX_s_1_2_2(mux_3028_nl, mux_tmp_139, fsm_output(7));
  mux_3043_nl <= MUX_s_1_2_2(mux_3042_nl, mux_3029_nl, fsm_output(5));
  mux_3016_nl <= MUX_s_1_2_2((fsm_output(8)), or_tmp_93, or_2855_cse);
  mux_3015_nl <= MUX_s_1_2_2(or_tmp_2795, mux_tmp_3014, fsm_output(9));
  mux_3017_nl <= MUX_s_1_2_2(mux_3016_nl, mux_3015_nl, fsm_output(0));
  mux_3018_nl <= MUX_s_1_2_2(mux_tmp_3014, mux_3017_nl, fsm_output(1));
  mux_3019_nl <= MUX_s_1_2_2((fsm_output(8)), mux_3018_nl, fsm_output(4));
  or_2851_nl <= (NOT (fsm_output(1))) OR (NOT (fsm_output(0))) OR (fsm_output(9))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(8))) OR (fsm_output(10));
  mux_3013_nl <= MUX_s_1_2_2(or_2851_nl, mux_tmp_130, fsm_output(4));
  mux_3020_nl <= MUX_s_1_2_2(mux_3019_nl, mux_3013_nl, fsm_output(7));
  mux_3009_nl <= MUX_s_1_2_2(mux_tmp_3008, mux_tmp_3007, fsm_output(0));
  mux_3010_nl <= MUX_s_1_2_2(or_tmp_2791, mux_3009_nl, fsm_output(1));
  mux_3011_nl <= MUX_s_1_2_2(mux_3010_nl, mux_tmp_130, fsm_output(4));
  or_2846_nl <= and_526_cse OR (fsm_output(9)) OR (fsm_output(2)) OR (NOT nor_tmp_405);
  mux_3005_nl <= MUX_s_1_2_2(mux_tmp_130, or_2846_nl, fsm_output(4));
  mux_3012_nl <= MUX_s_1_2_2(mux_3011_nl, mux_3005_nl, fsm_output(7));
  mux_3021_nl <= MUX_s_1_2_2(mux_3020_nl, mux_3012_nl, fsm_output(5));
  mux_3044_nl <= MUX_s_1_2_2(mux_3043_nl, mux_3021_nl, fsm_output(6));
  mux_3070_nl <= MUX_s_1_2_2(mux_3069_nl, mux_3044_nl, fsm_output(3));
  COMP_LOOP_mux1h_428_nl <= MUX1HOT_s_1_6_2((operator_66_true_div_cmp_z(0)), (tmp_10_lpi_4_dfm(0)),
      (z_out(5)), COMP_LOOP_nor_12_itm, COMP_LOOP_nor_11_itm, COMP_LOOP_nor_11_nl,
      STD_LOGIC_VECTOR'( COMP_LOOP_and_274_nl & and_dcpl_256 & and_dcpl_109 & not_tmp_557
      & (NOT mux_3070_nl) & COMP_LOOP_or_32_cse));
  or_2821_nl <= (fsm_output(9)) OR (NOT (fsm_output(8))) OR (fsm_output(4)) OR (fsm_output(1))
      OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(10));
  nor_671_nl <= NOT((fsm_output(6)) OR nand_159_cse);
  nor_672_nl <= NOT((fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(10)));
  mux_2986_nl <= MUX_s_1_2_2(nor_671_nl, nor_672_nl, fsm_output(1));
  nand_74_nl <= NOT((NOT((fsm_output(8)) OR (NOT (fsm_output(4))))) AND mux_2986_nl);
  or_2818_nl <= (NOT (fsm_output(8))) OR (fsm_output(4)) OR (NOT (fsm_output(1)))
      OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3))) OR (fsm_output(10));
  mux_2987_nl <= MUX_s_1_2_2(nand_74_nl, or_2818_nl, fsm_output(9));
  mux_2988_nl <= MUX_s_1_2_2(or_2821_nl, mux_2987_nl, fsm_output(5));
  or_3440_nl <= (fsm_output(7)) OR mux_2988_nl;
  or_3441_nl <= (fsm_output(5)) OR (fsm_output(9)) OR (NOT (fsm_output(8))) OR (fsm_output(4))
      OR (NOT (fsm_output(1))) OR (fsm_output(6)) OR (fsm_output(3)) OR (NOT (fsm_output(10)));
  and_447_nl <= (fsm_output(1)) AND (fsm_output(6)) AND (fsm_output(3)) AND (NOT
      (fsm_output(10)));
  nor_675_nl <= NOT((fsm_output(1)) OR (NOT (fsm_output(6))) OR (fsm_output(3)) OR
      (NOT (fsm_output(10))));
  mux_2983_nl <= MUX_s_1_2_2(and_447_nl, nor_675_nl, fsm_output(4));
  nand_73_nl <= NOT((fsm_output(8)) AND mux_2983_nl);
  or_2811_nl <= (fsm_output(8)) OR (NOT (fsm_output(4))) OR (fsm_output(1)) OR (fsm_output(6))
      OR (NOT (fsm_output(3))) OR (fsm_output(10));
  mux_2984_nl <= MUX_s_1_2_2(nand_73_nl, or_2811_nl, fsm_output(9));
  or_3442_nl <= (fsm_output(5)) OR mux_2984_nl;
  mux_2985_nl <= MUX_s_1_2_2(or_3441_nl, or_3442_nl, fsm_output(7));
  mux_2989_nl <= MUX_s_1_2_2(or_3440_nl, mux_2985_nl, fsm_output(2));
  nor_647_nl <= NOT((fsm_output(1)) OR (NOT (fsm_output(4))) OR (NOT (fsm_output(3)))
      OR (fsm_output(10)));
  mux_3075_nl <= MUX_s_1_2_2(nor_647_nl, nor_tmp_410, fsm_output(2));
  nor_646_nl <= NOT(CONV_SL_1_1(fsm_output(7 DOWNTO 5)/=STD_LOGIC_VECTOR'("100"))
      OR (NOT mux_3075_nl));
  nor_648_nl <= NOT((fsm_output(4)) OR nand_159_cse);
  nor_649_nl <= NOT((fsm_output(4)) OR (fsm_output(3)) OR (fsm_output(10)));
  mux_3074_nl <= MUX_s_1_2_2(nor_648_nl, nor_649_nl, fsm_output(1));
  and_439_nl <= (NOT (fsm_output(7))) AND (fsm_output(6)) AND (fsm_output(5)) AND
      (fsm_output(2)) AND mux_3074_nl;
  mux_3076_nl <= MUX_s_1_2_2(nor_646_nl, and_439_nl, fsm_output(8));
  nor_650_nl <= NOT((fsm_output(1)) OR (NOT (fsm_output(4))) OR (fsm_output(3)) OR
      (fsm_output(10)));
  mux_3072_nl <= MUX_s_1_2_2(nor_tmp_410, nor_650_nl, fsm_output(2));
  and_440_nl <= (NOT(CONV_SL_1_1(fsm_output(7 DOWNTO 5)/=STD_LOGIC_VECTOR'("001"))))
      AND mux_3072_nl;
  nor_651_nl <= NOT((fsm_output(6)) OR (fsm_output(5)) OR (fsm_output(2)) OR (NOT
      (fsm_output(1))) OR (fsm_output(4)) OR (fsm_output(3)) OR (fsm_output(10)));
  nor_652_nl <= NOT((NOT (fsm_output(6))) OR (fsm_output(5)) OR (fsm_output(2)) OR
      (fsm_output(1)) OR (NOT (fsm_output(4))) OR (fsm_output(3)) OR (fsm_output(10)));
  mux_3071_nl <= MUX_s_1_2_2(nor_651_nl, nor_652_nl, fsm_output(7));
  mux_3073_nl <= MUX_s_1_2_2(and_440_nl, mux_3071_nl, fsm_output(8));
  mux_3077_nl <= MUX_s_1_2_2(mux_3076_nl, mux_3073_nl, fsm_output(9));
  COMP_LOOP_mux1h_464_nl <= MUX1HOT_s_1_4_2((COMP_LOOP_k_9_4_sva_4_0(3)), COMP_LOOP_nor_134_itm,
      modExp_exp_1_7_1_sva, (COMP_LOOP_k_9_4_sva_4_0(4)), STD_LOGIC_VECTOR'( and_dcpl_257
      & and_dcpl_304 & (NOT mux_3494_itm) & not_tmp_688));
  or_3501_nl <= (NOT (fsm_output(7))) OR (fsm_output(5)) OR (fsm_output(9)) OR (NOT
      (fsm_output(2))) OR (NOT (fsm_output(8))) OR (fsm_output(6)) OR (NOT (fsm_output(10)));
  or_3502_nl <= (fsm_output(5)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(2)))
      OR (fsm_output(8)) OR (NOT (fsm_output(6))) OR (fsm_output(10));
  or_3503_nl <= (NOT (fsm_output(5))) OR (NOT (fsm_output(9))) OR (fsm_output(2))
      OR (NOT (fsm_output(8))) OR (NOT (fsm_output(6))) OR (fsm_output(10));
  mux_3517_nl <= MUX_s_1_2_2(or_3502_nl, or_3503_nl, fsm_output(7));
  mux_3518_nl <= MUX_s_1_2_2(or_3501_nl, mux_3517_nl, fsm_output(3));
  mux_3519_nl <= MUX_s_1_2_2(or_80_cse, mux_3518_nl, fsm_output(4));
  or_3133_nl <= (NOT (fsm_output(5))) OR (NOT (fsm_output(9))) OR (fsm_output(2))
      OR (fsm_output(8)) OR not_tmp_49;
  mux_3515_nl <= MUX_s_1_2_2(or_3133_nl, or_tmp_3053, fsm_output(7));
  or_3131_nl <= (NOT (fsm_output(5))) OR (NOT (fsm_output(9))) OR (fsm_output(2))
      OR (NOT (fsm_output(8))) OR (fsm_output(6)) OR (fsm_output(10));
  or_3130_nl <= (fsm_output(5)) OR (fsm_output(9)) OR (NOT (fsm_output(2))) OR (NOT
      (fsm_output(8))) OR (fsm_output(6)) OR (fsm_output(10));
  mux_3514_nl <= MUX_s_1_2_2(or_3131_nl, or_3130_nl, fsm_output(7));
  mux_3516_nl <= MUX_s_1_2_2(mux_3515_nl, mux_3514_nl, fsm_output(3));
  or_3504_nl <= (fsm_output(4)) OR mux_3516_nl;
  mux_3520_nl <= MUX_s_1_2_2(mux_3519_nl, or_3504_nl, fsm_output(1));
  or_3505_nl <= (NOT (fsm_output(3))) OR (fsm_output(7)) OR (NOT (fsm_output(5)))
      OR (fsm_output(9)) OR (NOT (fsm_output(2))) OR (NOT (fsm_output(8))) OR (fsm_output(6))
      OR (NOT (fsm_output(10)));
  nor_600_nl <= NOT((NOT (fsm_output(9))) OR (fsm_output(2)) OR (NOT (fsm_output(8)))
      OR (fsm_output(6)) OR (fsm_output(10)));
  nor_601_nl <= NOT((fsm_output(9)) OR (NOT (fsm_output(2))) OR (NOT (fsm_output(8)))
      OR (NOT (fsm_output(6))) OR (fsm_output(10)));
  mux_3511_nl <= MUX_s_1_2_2(nor_600_nl, nor_601_nl, fsm_output(5));
  nand_412_nl <= NOT((NOT((fsm_output(3)) OR (NOT (fsm_output(7))))) AND mux_3511_nl);
  mux_3512_nl <= MUX_s_1_2_2(or_3505_nl, nand_412_nl, fsm_output(4));
  or_3124_nl <= (NOT (fsm_output(5))) OR (fsm_output(9)) OR (NOT (fsm_output(2)))
      OR (NOT (fsm_output(8))) OR (fsm_output(6)) OR (fsm_output(10));
  or_3123_nl <= (fsm_output(5)) OR (NOT (fsm_output(9))) OR (fsm_output(2)) OR (fsm_output(8))
      OR (NOT (fsm_output(6))) OR (fsm_output(10));
  mux_3509_nl <= MUX_s_1_2_2(or_3124_nl, or_3123_nl, fsm_output(7));
  or_3506_nl <= (fsm_output(3)) OR mux_3509_nl;
  or_3120_nl <= (NOT (fsm_output(5))) OR (fsm_output(9)) OR (fsm_output(2)) OR nand_142_cse;
  mux_3508_nl <= MUX_s_1_2_2(or_tmp_3053, or_3120_nl, fsm_output(7));
  nand_413_nl <= NOT((fsm_output(3)) AND (NOT mux_3508_nl));
  mux_3510_nl <= MUX_s_1_2_2(or_3506_nl, nand_413_nl, fsm_output(4));
  mux_3513_nl <= MUX_s_1_2_2(mux_3512_nl, mux_3510_nl, fsm_output(1));
  mux_3521_nl <= MUX_s_1_2_2(mux_3520_nl, mux_3513_nl, fsm_output(0));
  COMP_LOOP_nor_12_nl <= NOT((z_out_2_12_1(3)) OR (z_out_2_12_1(2)) OR (z_out_2_12_1(0)));
  mux_3610_nl <= MUX_s_1_2_2(nand_tmp_4, mux_155_cse, fsm_output(2));
  mux_3611_nl <= MUX_s_1_2_2(mux_3610_nl, mux_tmp_3551, fsm_output(0));
  mux_3609_nl <= MUX_s_1_2_2(mux_tmp_3551, mux_tmp_3547, fsm_output(0));
  mux_3612_nl <= MUX_s_1_2_2(mux_3611_nl, mux_3609_nl, fsm_output(1));
  mux_3606_nl <= MUX_s_1_2_2(mux_tmp_130, mux_tmp_141, fsm_output(4));
  mux_3607_nl <= MUX_s_1_2_2(mux_3606_nl, or_tmp_96, fsm_output(2));
  mux_3605_nl <= MUX_s_1_2_2(mux_161_cse, or_tmp_96, fsm_output(2));
  mux_3608_nl <= MUX_s_1_2_2(mux_3607_nl, mux_3605_nl, or_3388_cse);
  mux_3613_nl <= MUX_s_1_2_2(mux_3612_nl, mux_3608_nl, fsm_output(7));
  mux_3602_nl <= MUX_s_1_2_2(mux_tmp_3576, mux_tmp_3574, fsm_output(0));
  mux_3603_nl <= MUX_s_1_2_2(mux_tmp_3577, mux_3602_nl, fsm_output(1));
  mux_3604_nl <= MUX_s_1_2_2(mux_3603_nl, mux_tmp_139, fsm_output(7));
  mux_3614_nl <= MUX_s_1_2_2(mux_3613_nl, mux_3604_nl, fsm_output(5));
  or_3192_nl <= (NOT(and_529_cse OR (fsm_output(4)))) OR (fsm_output(9));
  mux_3599_nl <= MUX_s_1_2_2(or_tmp_93, (fsm_output(8)), or_3192_nl);
  mux_3596_nl <= MUX_s_1_2_2(mux_498_cse, mux_171_cse, fsm_output(2));
  mux_493_nl <= MUX_s_1_2_2(or_469_cse, mux_tmp_130, fsm_output(4));
  mux_3595_nl <= MUX_s_1_2_2(mux_498_cse, mux_493_nl, fsm_output(2));
  mux_3597_nl <= MUX_s_1_2_2(mux_3596_nl, mux_3595_nl, fsm_output(0));
  mux_454_nl <= MUX_s_1_2_2(mux_tmp_165, or_tmp_88, fsm_output(4));
  mux_3591_nl <= MUX_s_1_2_2(mux_454_nl, nand_tmp_4, fsm_output(2));
  mux_3588_nl <= MUX_s_1_2_2(mux_171_cse, nand_tmp_4, fsm_output(2));
  mux_3592_nl <= MUX_s_1_2_2(mux_3591_nl, mux_3588_nl, fsm_output(0));
  mux_3598_nl <= MUX_s_1_2_2(mux_3597_nl, mux_3592_nl, fsm_output(1));
  mux_3600_nl <= MUX_s_1_2_2(mux_3599_nl, mux_3598_nl, fsm_output(7));
  mux_3584_nl <= MUX_s_1_2_2(or_2387_cse, mux_tmp_130, fsm_output(4));
  mux_3585_nl <= MUX_s_1_2_2(mux_3584_nl, nand_tmp_4, or_2368_cse);
  and_364_nl <= or_3388_cse AND (fsm_output(2)) AND (fsm_output(4));
  mux_3583_nl <= MUX_s_1_2_2(mux_tmp_130, mux_tmp_141, and_364_nl);
  mux_3586_nl <= MUX_s_1_2_2(mux_3585_nl, mux_3583_nl, fsm_output(7));
  mux_3601_nl <= MUX_s_1_2_2(mux_3600_nl, mux_3586_nl, fsm_output(5));
  mux_3615_nl <= MUX_s_1_2_2(mux_3614_nl, mux_3601_nl, fsm_output(6));
  mux_3578_nl <= MUX_s_1_2_2(mux_tmp_3577, mux_tmp_3576, fsm_output(0));
  mux_3579_nl <= MUX_s_1_2_2(mux_3578_nl, mux_tmp_3574, fsm_output(1));
  mux_3580_nl <= MUX_s_1_2_2(mux_tmp_130, mux_3579_nl, fsm_output(7));
  mux_481_nl <= MUX_s_1_2_2(or_3008_cse, (fsm_output(8)), fsm_output(4));
  mux_3569_nl <= MUX_s_1_2_2(mux_340_cse, mux_481_nl, fsm_output(2));
  mux_3565_nl <= MUX_s_1_2_2(mux_tmp_141, mux_tmp_139, fsm_output(4));
  mux_3566_nl <= MUX_s_1_2_2(mux_3565_nl, or_163_cse, fsm_output(2));
  mux_3570_nl <= MUX_s_1_2_2(mux_3569_nl, mux_3566_nl, fsm_output(0));
  mux_3562_nl <= MUX_s_1_2_2(or_3008_cse, mux_tmp_139, fsm_output(4));
  mux_3563_nl <= MUX_s_1_2_2(mux_3562_nl, or_163_cse, fsm_output(2));
  mux_3571_nl <= MUX_s_1_2_2(mux_3570_nl, mux_3563_nl, fsm_output(1));
  mux_3572_nl <= MUX_s_1_2_2(mux_3571_nl, mux_tmp_139, fsm_output(7));
  mux_3581_nl <= MUX_s_1_2_2(mux_3580_nl, mux_3572_nl, fsm_output(5));
  and_365_nl <= (NOT((fsm_output(2)) AND (fsm_output(4)))) AND (fsm_output(9));
  mux_3557_nl <= MUX_s_1_2_2(or_tmp_93, (fsm_output(8)), and_365_nl);
  mux_3556_nl <= MUX_s_1_2_2(mux_3555_cse, or_2387_cse, and_366_cse);
  mux_3558_nl <= MUX_s_1_2_2(mux_3557_nl, mux_3556_nl, and_526_cse);
  mux_3554_nl <= MUX_s_1_2_2(nand_tmp_4, mux_tmp_131, and_536_cse);
  mux_3559_nl <= MUX_s_1_2_2(mux_3558_nl, mux_3554_nl, fsm_output(7));
  or_3177_nl <= (NOT((fsm_output(2)) OR (fsm_output(4)))) OR (fsm_output(9));
  mux_3546_nl <= MUX_s_1_2_2((NOT (fsm_output(8))), or_tmp_88, or_3177_nl);
  mux_3548_nl <= MUX_s_1_2_2(mux_tmp_3547, mux_3546_nl, fsm_output(0));
  mux_3552_nl <= MUX_s_1_2_2(mux_tmp_3551, mux_3548_nl, fsm_output(1));
  mux_3545_nl <= MUX_s_1_2_2(mux_161_cse, or_tmp_96, or_2377_cse);
  mux_3553_nl <= MUX_s_1_2_2(mux_3552_nl, mux_3545_nl, fsm_output(7));
  mux_3560_nl <= MUX_s_1_2_2(mux_3559_nl, mux_3553_nl, fsm_output(5));
  mux_3582_nl <= MUX_s_1_2_2(mux_3581_nl, mux_3560_nl, fsm_output(6));
  mux_3616_nl <= MUX_s_1_2_2(mux_3615_nl, mux_3582_nl, fsm_output(3));
  mux_3627_nl <= MUX_s_1_2_2(mux_tmp_3618, or_tmp_3135, fsm_output(3));
  nor_565_nl <= NOT((fsm_output(5)) OR (NOT (fsm_output(7))) OR mux_3627_nl);
  or_3213_nl <= (fsm_output(2)) OR (NOT (fsm_output(1))) OR (fsm_output(8)) OR not_tmp_49;
  or_3211_nl <= (fsm_output(2)) OR (NOT (fsm_output(1))) OR (NOT (fsm_output(8)))
      OR (fsm_output(6)) OR (fsm_output(10));
  mux_3626_nl <= MUX_s_1_2_2(or_3213_nl, or_3211_nl, fsm_output(3));
  nor_566_nl <= NOT((NOT (fsm_output(5))) OR (fsm_output(7)) OR mux_3626_nl);
  mux_3628_nl <= MUX_s_1_2_2(nor_565_nl, nor_566_nl, fsm_output(9));
  nor_567_nl <= NOT((fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(3)) OR
      (NOT (fsm_output(2))) OR (fsm_output(1)) OR (NOT (fsm_output(8))) OR (fsm_output(6))
      OR (NOT (fsm_output(10))));
  nor_568_nl <= NOT((fsm_output(7)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(2)))
      OR (fsm_output(1)) OR (fsm_output(8)) OR (NOT (fsm_output(6))) OR (fsm_output(10)));
  nor_569_nl <= NOT((NOT (fsm_output(7))) OR (NOT (fsm_output(3))) OR (fsm_output(2))
      OR (fsm_output(1)) OR (NOT (fsm_output(8))) OR (NOT (fsm_output(6))) OR (fsm_output(10)));
  mux_3624_nl <= MUX_s_1_2_2(nor_568_nl, nor_569_nl, fsm_output(5));
  mux_3625_nl <= MUX_s_1_2_2(nor_567_nl, mux_3624_nl, fsm_output(9));
  mux_3629_nl <= MUX_s_1_2_2(mux_3628_nl, mux_3625_nl, fsm_output(4));
  or_3203_nl <= (NOT (fsm_output(2))) OR (fsm_output(1)) OR (NOT (fsm_output(8)))
      OR (fsm_output(6)) OR (NOT (fsm_output(10)));
  mux_3621_nl <= MUX_s_1_2_2(or_tmp_3135, or_3203_nl, fsm_output(3));
  nor_570_nl <= NOT((NOT (fsm_output(5))) OR (fsm_output(7)) OR mux_3621_nl);
  nor_571_nl <= NOT((fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(3)) OR
      (fsm_output(2)) OR (NOT (fsm_output(1))) OR (fsm_output(8)) OR (NOT (fsm_output(6)))
      OR (fsm_output(10)));
  mux_3622_nl <= MUX_s_1_2_2(nor_570_nl, nor_571_nl, fsm_output(9));
  nor_572_nl <= NOT((fsm_output(7)) OR (NOT (fsm_output(3))) OR mux_tmp_3618);
  nor_573_nl <= NOT((NOT (fsm_output(2))) OR (fsm_output(1)) OR (NOT (fsm_output(8)))
      OR (NOT (fsm_output(6))) OR (fsm_output(10)));
  nor_574_nl <= NOT((fsm_output(2)) OR (NOT((fsm_output(1)) AND (fsm_output(8)) AND
      (fsm_output(6)) AND (fsm_output(10)))));
  mux_3617_nl <= MUX_s_1_2_2(nor_573_nl, nor_574_nl, fsm_output(3));
  and_362_nl <= (fsm_output(7)) AND mux_3617_nl;
  mux_3619_nl <= MUX_s_1_2_2(nor_572_nl, and_362_nl, fsm_output(5));
  nor_575_nl <= NOT((fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(3)) OR
      (fsm_output(2)) OR (fsm_output(1)) OR (NOT (fsm_output(8))) OR (fsm_output(6))
      OR (fsm_output(10)));
  mux_3620_nl <= MUX_s_1_2_2(mux_3619_nl, nor_575_nl, fsm_output(9));
  mux_3623_nl <= MUX_s_1_2_2(mux_3622_nl, mux_3620_nl, fsm_output(4));
  mux_3630_nl <= MUX_s_1_2_2(mux_3629_nl, mux_3623_nl, fsm_output(0));
  COMP_LOOP_mux1h_474_nl <= MUX1HOT_s_1_3_2(COMP_LOOP_nor_12_itm, COMP_LOOP_nor_134_itm,
      COMP_LOOP_nor_12_nl, STD_LOGIC_VECTOR'( (NOT mux_3616_nl) & mux_3630_nl & COMP_LOOP_or_32_cse));
  or_3171_nl <= (fsm_output(4)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(6)))
      OR (NOT (fsm_output(8))) OR (fsm_output(10));
  mux_3540_nl <= MUX_s_1_2_2(or_tmp_3095, or_3171_nl, fsm_output(3));
  nor_578_nl <= NOT((fsm_output(7)) OR (NOT (fsm_output(5))) OR mux_3540_nl);
  nor_579_nl <= NOT((fsm_output(5)) OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(9))
      OR (fsm_output(6)) OR nand_138_cse);
  nor_580_nl <= NOT((fsm_output(5)) OR (NOT (fsm_output(3))) OR (fsm_output(4)) OR
      (fsm_output(9)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(8))) OR (fsm_output(10)));
  mux_3539_nl <= MUX_s_1_2_2(nor_579_nl, nor_580_nl, fsm_output(7));
  mux_3541_nl <= MUX_s_1_2_2(nor_578_nl, mux_3539_nl, fsm_output(2));
  nand_411_nl <= NOT((fsm_output(1)) AND mux_3541_nl);
  nand_139_nl <= NOT((fsm_output(4)) AND (fsm_output(9)) AND (fsm_output(6)) AND
      (fsm_output(8)) AND (NOT (fsm_output(10))));
  mux_3537_nl <= MUX_s_1_2_2(nand_139_nl, or_tmp_3095, fsm_output(3));
  or_3166_nl <= (NOT (fsm_output(7))) OR (fsm_output(5)) OR mux_3537_nl;
  nor_582_nl <= NOT((NOT (fsm_output(4))) OR (NOT (fsm_output(9))) OR (fsm_output(6))
      OR (fsm_output(8)) OR (fsm_output(10)));
  nor_583_nl <= NOT((fsm_output(4)) OR (fsm_output(9)) OR nand_142_cse);
  mux_3536_nl <= MUX_s_1_2_2(nor_582_nl, nor_583_nl, fsm_output(3));
  nand_104_nl <= NOT((NOT((fsm_output(7)) OR (NOT (fsm_output(5))))) AND mux_3536_nl);
  mux_3538_nl <= MUX_s_1_2_2(or_3166_nl, nand_104_nl, fsm_output(2));
  or_3499_nl <= (fsm_output(1)) OR mux_3538_nl;
  mux_3542_nl <= MUX_s_1_2_2(nand_411_nl, or_3499_nl, fsm_output(0));
  or_3228_nl <= (fsm_output(9)) OR (fsm_output(6)) OR mux_tmp_3632;
  or_3226_nl <= (NOT (fsm_output(6))) OR (fsm_output(5)) OR (NOT (fsm_output(7)))
      OR (fsm_output(3)) OR (NOT((fsm_output(8)) AND (fsm_output(4)) AND (fsm_output(10))));
  or_3224_nl <= (fsm_output(6)) OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR (NOT
      (fsm_output(3))) OR (fsm_output(8)) OR (NOT (fsm_output(4))) OR (fsm_output(10));
  mux_3634_nl <= MUX_s_1_2_2(or_3226_nl, or_3224_nl, fsm_output(9));
  mux_3635_nl <= MUX_s_1_2_2(or_3228_nl, mux_3634_nl, fsm_output(2));
  nor_562_nl <= NOT((fsm_output(1)) OR mux_3635_nl);
  nor_563_nl <= NOT((NOT (fsm_output(9))) OR (fsm_output(6)) OR mux_tmp_3632);
  or_3217_nl <= (fsm_output(5)) OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3)))
      OR (fsm_output(8)) OR not_tmp_39;
  or_3215_nl <= (NOT (fsm_output(5))) OR (fsm_output(7)) OR (fsm_output(3)) OR (NOT
      (fsm_output(8))) OR (fsm_output(4)) OR (fsm_output(10));
  mux_3631_nl <= MUX_s_1_2_2(or_3217_nl, or_3215_nl, fsm_output(6));
  nor_564_nl <= NOT((fsm_output(9)) OR mux_3631_nl);
  mux_3633_nl <= MUX_s_1_2_2(nor_563_nl, nor_564_nl, fsm_output(2));
  and_361_nl <= (fsm_output(1)) AND mux_3633_nl;
  mux_3636_nl <= MUX_s_1_2_2(nor_562_nl, and_361_nl, fsm_output(0));
  COMP_LOOP_nor_14_nl <= NOT((z_out_2_12_1(3)) OR (z_out_2_12_1(1)) OR (z_out_2_12_1(0)));
  mux_3637_nl <= MUX_s_1_2_2(mux_tmp_3457, mux_tmp_3474, fsm_output(6));
  mux_3638_nl <= MUX_s_1_2_2((NOT mux_3485_itm), mux_3637_nl, fsm_output(4));
  mux_3639_nl <= MUX_s_1_2_2(mux_3638_nl, mux_tmp_3481, fsm_output(1));
  mux_3640_nl <= MUX_s_1_2_2(mux_tmp_3491, mux_3639_nl, fsm_output(0));
  mux_3641_nl <= MUX_s_1_2_2(mux_3640_nl, mux_tmp_3472, fsm_output(9));
  mux_3642_nl <= MUX_s_1_2_2(mux_3641_nl, mux_tmp_3453, fsm_output(10));
  COMP_LOOP_mux1h_477_nl <= MUX1HOT_s_1_4_2((COMP_LOOP_k_9_4_sva_4_0(4)), COMP_LOOP_nor_137_itm,
      COMP_LOOP_nor_134_itm, COMP_LOOP_nor_14_nl, STD_LOGIC_VECTOR'( and_dcpl_257
      & not_tmp_701 & (NOT mux_3642_nl) & COMP_LOOP_or_32_cse));
  or_3240_nl <= (fsm_output(9)) OR (fsm_output(3)) OR (fsm_output(4)) OR (NOT (fsm_output(8)))
      OR (fsm_output(10));
  or_3239_nl <= (fsm_output(9)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(4)))
      OR (fsm_output(8)) OR (NOT (fsm_output(10)));
  mux_3647_nl <= MUX_s_1_2_2(or_3240_nl, or_3239_nl, fsm_output(5));
  or_3241_nl <= CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00")) OR mux_3647_nl;
  or_3236_nl <= (NOT (fsm_output(6))) OR (fsm_output(5)) OR (fsm_output(9)) OR (NOT
      (fsm_output(3))) OR (NOT (fsm_output(4))) OR (fsm_output(8)) OR (fsm_output(10));
  or_3235_nl <= (fsm_output(5)) OR (fsm_output(9)) OR (NOT (fsm_output(3))) OR (NOT
      (fsm_output(4))) OR (fsm_output(8)) OR (fsm_output(10));
  or_3234_nl <= (fsm_output(5)) OR (NOT (fsm_output(9))) OR (fsm_output(3)) OR (NOT
      (fsm_output(4))) OR (NOT (fsm_output(8))) OR (fsm_output(10));
  mux_3645_nl <= MUX_s_1_2_2(or_3235_nl, or_3234_nl, fsm_output(6));
  mux_3646_nl <= MUX_s_1_2_2(or_3236_nl, mux_3645_nl, fsm_output(7));
  mux_3648_nl <= MUX_s_1_2_2(or_3241_nl, mux_3646_nl, fsm_output(0));
  or_3497_nl <= (fsm_output(2)) OR mux_3648_nl;
  or_3498_nl <= (fsm_output(0)) OR (fsm_output(7)) OR (NOT (fsm_output(6))) OR (NOT
      (fsm_output(5))) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(3))) OR (fsm_output(4))
      OR (NOT (fsm_output(8))) OR (fsm_output(10));
  nor_560_nl <= NOT((NOT (fsm_output(6))) OR (NOT (fsm_output(5))) OR (fsm_output(9))
      OR (fsm_output(3)) OR (fsm_output(4)) OR (NOT (fsm_output(8))) OR (fsm_output(10)));
  nor_561_nl <= NOT((fsm_output(6)) OR (fsm_output(5)) OR (fsm_output(9)) OR (NOT
      (fsm_output(3))) OR (NOT (fsm_output(4))) OR (fsm_output(8)) OR (NOT (fsm_output(10))));
  mux_3643_nl <= MUX_s_1_2_2(nor_560_nl, nor_561_nl, fsm_output(7));
  nand_410_nl <= NOT((fsm_output(0)) AND mux_3643_nl);
  mux_3644_nl <= MUX_s_1_2_2(or_3498_nl, nand_410_nl, fsm_output(2));
  mux_3649_nl <= MUX_s_1_2_2(or_3497_nl, mux_3644_nl, fsm_output(1));
  nor_555_nl <= NOT((fsm_output(5)) OR (NOT (fsm_output(2))) OR (NOT (fsm_output(1)))
      OR (fsm_output(3)) OR (fsm_output(4)) OR (NOT (fsm_output(8))) OR (fsm_output(9))
      OR (fsm_output(6)) OR (NOT (fsm_output(10))));
  or_3253_nl <= (NOT (fsm_output(4))) OR (NOT (fsm_output(8))) OR (fsm_output(9))
      OR not_tmp_49;
  mux_3653_nl <= MUX_s_1_2_2(or_3253_nl, or_tmp_3176, fsm_output(3));
  or_3251_nl <= (NOT (fsm_output(3))) OR (fsm_output(4)) OR (NOT (fsm_output(8)))
      OR (fsm_output(9)) OR (NOT (fsm_output(6))) OR (fsm_output(10));
  mux_3654_nl <= MUX_s_1_2_2(mux_3653_nl, or_3251_nl, fsm_output(1));
  nor_556_nl <= NOT((fsm_output(5)) OR (NOT (fsm_output(2))) OR mux_3654_nl);
  mux_3655_nl <= MUX_s_1_2_2(nor_555_nl, nor_556_nl, fsm_output(7));
  or_3249_nl <= (fsm_output(2)) OR (NOT (fsm_output(1))) OR (fsm_output(3)) OR (fsm_output(4))
      OR (NOT (fsm_output(8))) OR (NOT (fsm_output(9))) OR (fsm_output(6)) OR (fsm_output(10));
  nand_383_nl <= NOT((fsm_output(1)) AND (fsm_output(3)) AND (fsm_output(4)) AND
      (NOT (fsm_output(8))) AND (fsm_output(9)) AND (NOT (fsm_output(6))) AND (fsm_output(10)));
  or_3244_nl <= (fsm_output(4)) OR (NOT (fsm_output(8))) OR (fsm_output(9)) OR not_tmp_49;
  mux_3650_nl <= MUX_s_1_2_2(or_tmp_3176, or_3244_nl, fsm_output(3));
  or_3246_nl <= (fsm_output(1)) OR mux_3650_nl;
  mux_3651_nl <= MUX_s_1_2_2(nand_383_nl, or_3246_nl, fsm_output(2));
  mux_3652_nl <= MUX_s_1_2_2(or_3249_nl, mux_3651_nl, fsm_output(5));
  nor_557_nl <= NOT((fsm_output(7)) OR mux_3652_nl);
  mux_3656_nl <= MUX_s_1_2_2(mux_3655_nl, nor_557_nl, fsm_output(0));
  COMP_LOOP_nor_17_nl <= NOT(CONV_SL_1_1(z_out_2_12_1(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000")));
  COMP_LOOP_mux1h_479_nl <= MUX1HOT_s_1_3_2(COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm,
      COMP_LOOP_nor_137_itm, COMP_LOOP_nor_17_nl, STD_LOGIC_VECTOR'( not_tmp_701
      & (NOT mux_3494_itm) & COMP_LOOP_or_32_cse));
  or_3266_nl <= (NOT (fsm_output(1))) OR (fsm_output(2)) OR (fsm_output(6)) OR (NOT
      (fsm_output(9)));
  mux_3660_nl <= MUX_s_1_2_2(or_3417_cse, or_3266_nl, fsm_output(0));
  nand_130_nl <= NOT((fsm_output(0)) AND (fsm_output(1)) AND (fsm_output(2)) AND
      (fsm_output(6)) AND (NOT (fsm_output(9))));
  mux_3661_nl <= MUX_s_1_2_2(mux_3660_nl, nand_130_nl, fsm_output(5));
  nor_552_nl <= NOT((fsm_output(7)) OR mux_3661_nl);
  nor_553_nl <= NOT((NOT (fsm_output(7))) OR (fsm_output(5)) OR (fsm_output(0)) OR
      (NOT (fsm_output(1))) OR (NOT (fsm_output(2))) OR (NOT (fsm_output(6))) OR
      (fsm_output(9)));
  mux_3662_nl <= MUX_s_1_2_2(nor_552_nl, nor_553_nl, fsm_output(3));
  nand_389_nl <= NOT((fsm_output(8)) AND mux_3662_nl);
  or_3261_nl <= (NOT (fsm_output(1))) OR (fsm_output(2)) OR (fsm_output(6)) OR (fsm_output(9));
  mux_3658_nl <= MUX_s_1_2_2(or_3261_nl, or_tmp_3190, fsm_output(0));
  or_3353_nl <= (fsm_output(7)) OR (NOT (fsm_output(5))) OR mux_3658_nl;
  mux_3657_nl <= MUX_s_1_2_2(or_tmp_3190, or_3417_cse, fsm_output(0));
  or_3260_nl <= (NOT (fsm_output(7))) OR (fsm_output(5)) OR mux_3657_nl;
  mux_3659_nl <= MUX_s_1_2_2(or_3353_nl, or_3260_nl, fsm_output(3));
  or_3443_nl <= (fsm_output(8)) OR mux_3659_nl;
  mux_3663_nl <= MUX_s_1_2_2(nand_389_nl, or_3443_nl, fsm_output(4));
  nor_547_nl <= NOT((fsm_output(3)) OR (NOT (fsm_output(8))) OR (fsm_output(6)) OR
      (NOT (fsm_output(1))) OR (fsm_output(0)) OR (fsm_output(4)) OR (fsm_output(9))
      OR not_tmp_253);
  or_3282_nl <= (fsm_output(0)) OR (NOT (fsm_output(4))) OR (fsm_output(9)) OR (fsm_output(2))
      OR (NOT (fsm_output(10)));
  nand_382_nl <= NOT((fsm_output(0)) AND (fsm_output(4)) AND (fsm_output(9)) AND
      (NOT (fsm_output(2))) AND (fsm_output(10)));
  mux_3667_nl <= MUX_s_1_2_2(or_3282_nl, nand_382_nl, fsm_output(1));
  nor_548_nl <= NOT((fsm_output(6)) OR mux_3667_nl);
  nor_549_nl <= NOT((NOT (fsm_output(0))) OR (fsm_output(4)) OR (fsm_output(9)) OR
      not_tmp_253);
  nor_550_nl <= NOT((fsm_output(0)) OR (fsm_output(4)) OR (NOT (fsm_output(9))) OR
      (fsm_output(2)) OR (fsm_output(10)));
  mux_3666_nl <= MUX_s_1_2_2(nor_549_nl, nor_550_nl, fsm_output(1));
  and_358_nl <= (fsm_output(6)) AND mux_3666_nl;
  mux_3668_nl <= MUX_s_1_2_2(nor_548_nl, and_358_nl, fsm_output(8));
  and_357_nl <= (fsm_output(3)) AND mux_3668_nl;
  mux_3669_nl <= MUX_s_1_2_2(nor_547_nl, and_357_nl, fsm_output(5));
  or_3273_nl <= (NOT (fsm_output(4))) OR (fsm_output(9)) OR not_tmp_253;
  or_3271_nl <= (NOT (fsm_output(4))) OR (NOT (fsm_output(9))) OR (fsm_output(2))
      OR (fsm_output(10));
  mux_3664_nl <= MUX_s_1_2_2(or_3273_nl, or_3271_nl, fsm_output(0));
  or_3274_nl <= (NOT (fsm_output(8))) OR (NOT (fsm_output(6))) OR (fsm_output(1))
      OR mux_3664_nl;
  or_3269_nl <= (fsm_output(8)) OR (fsm_output(6)) OR (NOT (fsm_output(1))) OR (NOT
      (fsm_output(0))) OR (NOT (fsm_output(4))) OR (fsm_output(9)) OR not_tmp_253;
  mux_3665_nl <= MUX_s_1_2_2(or_3274_nl, or_3269_nl, fsm_output(3));
  nor_551_nl <= NOT((fsm_output(5)) OR mux_3665_nl);
  mux_3670_nl <= MUX_s_1_2_2(mux_3669_nl, nor_551_nl, fsm_output(7));
  mux_3761_nl <= MUX_s_1_2_2((NOT mux_tmp_236), mux_tmp_228, fsm_output(7));
  mux_3762_nl <= MUX_s_1_2_2(mux_3761_nl, mux_tmp_3720, fsm_output(1));
  mux_3763_nl <= MUX_s_1_2_2(mux_tmp_3724, mux_3762_nl, and_366_cse);
  mux_3755_nl <= MUX_s_1_2_2(or_361_cse, and_757_cse, fsm_output(5));
  mux_3756_nl <= MUX_s_1_2_2(mux_3755_nl, or_tmp_114, fsm_output(7));
  mux_3757_nl <= MUX_s_1_2_2(mux_3756_nl, mux_tmp_3753, fsm_output(0));
  mux_3758_nl <= MUX_s_1_2_2(mux_3757_nl, mux_tmp_3674, fsm_output(1));
  mux_3754_nl <= MUX_s_1_2_2(mux_tmp_3753, mux_tmp_3705, and_526_cse);
  mux_3759_nl <= MUX_s_1_2_2(mux_3758_nl, mux_3754_nl, fsm_output(2));
  or_3302_nl <= (fsm_output(5)) OR (fsm_output(9)) OR (NOT (fsm_output(10)));
  mux_3750_nl <= MUX_s_1_2_2(mux_tmp_231, or_3302_nl, fsm_output(7));
  mux_3751_nl <= MUX_s_1_2_2(mux_tmp_3698, mux_3750_nl, or_3388_cse);
  mux_3752_nl <= MUX_s_1_2_2(mux_3751_nl, or_tmp_3224, fsm_output(2));
  mux_3760_nl <= MUX_s_1_2_2(mux_3759_nl, mux_3752_nl, fsm_output(4));
  mux_3764_nl <= MUX_s_1_2_2(mux_3763_nl, mux_3760_nl, fsm_output(8));
  mux_3744_nl <= MUX_s_1_2_2((NOT nand_tmp_7), mux_tmp_3736, fsm_output(7));
  nor_546_nl <= NOT((NOT (fsm_output(5))) OR (fsm_output(10)));
  mux_3743_nl <= MUX_s_1_2_2(nor_546_nl, mux_tmp_3736, fsm_output(7));
  mux_3745_nl <= MUX_s_1_2_2(mux_3744_nl, mux_3743_nl, fsm_output(0));
  mux_3742_nl <= MUX_s_1_2_2(mux_tmp_3737, mux_tmp_3739, fsm_output(0));
  mux_3746_nl <= MUX_s_1_2_2(mux_3745_nl, mux_3742_nl, fsm_output(1));
  mux_3740_nl <= MUX_s_1_2_2(mux_tmp_3739, mux_tmp_3737, fsm_output(0));
  mux_3741_nl <= MUX_s_1_2_2(mux_3740_nl, mux_tmp_3691, fsm_output(1));
  mux_3747_nl <= MUX_s_1_2_2(mux_3746_nl, mux_3741_nl, fsm_output(2));
  mux_3748_nl <= MUX_s_1_2_2(mux_3747_nl, mux_tmp_3691, fsm_output(4));
  or_3298_nl <= (fsm_output(5)) OR (fsm_output(9)) OR (fsm_output(10));
  mux_3733_nl <= MUX_s_1_2_2(or_3298_nl, nand_tmp_7, fsm_output(7));
  mux_3734_nl <= MUX_s_1_2_2(mux_tmp_3681, mux_3733_nl, and_529_cse);
  and_349_nl <= (fsm_output(1)) AND (fsm_output(7));
  mux_3731_nl <= MUX_s_1_2_2(mux_tmp_215, nor_tmp_23, and_349_nl);
  mux_3729_nl <= MUX_s_1_2_2(mux_tmp_215, nor_tmp_23, fsm_output(7));
  mux_3728_nl <= MUX_s_1_2_2(mux_tmp_215, mux_tmp_236, fsm_output(7));
  mux_3730_nl <= MUX_s_1_2_2(mux_3729_nl, mux_3728_nl, or_3388_cse);
  mux_3732_nl <= MUX_s_1_2_2(mux_3731_nl, mux_3730_nl, fsm_output(2));
  mux_3735_nl <= MUX_s_1_2_2(mux_3734_nl, mux_3732_nl, fsm_output(4));
  mux_3749_nl <= MUX_s_1_2_2(mux_3748_nl, mux_3735_nl, fsm_output(8));
  mux_3765_nl <= MUX_s_1_2_2(mux_3764_nl, mux_3749_nl, fsm_output(6));
  mux_3719_nl <= MUX_s_1_2_2((NOT or_tmp_114), mux_tmp_228, fsm_output(7));
  mux_3721_nl <= MUX_s_1_2_2(mux_tmp_3720, mux_3719_nl, fsm_output(0));
  mux_3716_nl <= MUX_s_1_2_2((NOT and_757_cse), and_757_cse, fsm_output(5));
  mux_3717_nl <= MUX_s_1_2_2(mux_3716_nl, mux_259_cse, fsm_output(7));
  mux_3722_nl <= MUX_s_1_2_2(mux_3721_nl, mux_3717_nl, fsm_output(1));
  mux_3713_nl <= MUX_s_1_2_2((NOT or_tmp_114), mux_259_cse, fsm_output(7));
  mux_3711_nl <= MUX_s_1_2_2((NOT or_tmp_114), and_757_cse, fsm_output(7));
  mux_3714_nl <= MUX_s_1_2_2(mux_3713_nl, mux_3711_nl, fsm_output(0));
  mux_3710_nl <= MUX_s_1_2_2((NOT or_tmp_114), nor_tmp_23, fsm_output(7));
  mux_3715_nl <= MUX_s_1_2_2(mux_3714_nl, mux_3710_nl, fsm_output(1));
  mux_3723_nl <= MUX_s_1_2_2(mux_3722_nl, mux_3715_nl, fsm_output(2));
  mux_3725_nl <= MUX_s_1_2_2(mux_tmp_3724, mux_3723_nl, fsm_output(4));
  or_3295_nl <= and_350_cse OR and_757_cse;
  mux_3706_nl <= MUX_s_1_2_2(mux_tmp_3705, or_3295_nl, fsm_output(0));
  mux_3707_nl <= MUX_s_1_2_2(mux_3706_nl, mux_tmp_3701, fsm_output(1));
  mux_3699_nl <= MUX_s_1_2_2(mux_tmp_231, or_tmp_114, fsm_output(7));
  mux_3702_nl <= MUX_s_1_2_2(mux_tmp_3701, mux_3699_nl, fsm_output(0));
  mux_3703_nl <= MUX_s_1_2_2(mux_3702_nl, mux_tmp_3698, fsm_output(1));
  mux_3708_nl <= MUX_s_1_2_2(mux_3707_nl, mux_3703_nl, fsm_output(2));
  mux_3709_nl <= MUX_s_1_2_2(mux_3708_nl, or_tmp_3224, fsm_output(4));
  mux_3726_nl <= MUX_s_1_2_2(mux_3725_nl, mux_3709_nl, fsm_output(8));
  mux_3689_nl <= MUX_s_1_2_2((NOT or_2414_cse), or_tmp_104, fsm_output(5));
  mux_3690_nl <= MUX_s_1_2_2(mux_3689_nl, or_361_cse, fsm_output(7));
  mux_3692_nl <= MUX_s_1_2_2(mux_tmp_3691, mux_3690_nl, fsm_output(1));
  nand_380_nl <= NOT((NOT((fsm_output(5)) AND (fsm_output(9)))) AND (fsm_output(10)));
  mux_3687_nl <= MUX_s_1_2_2(nand_380_nl, or_361_cse, fsm_output(7));
  mux_3685_nl <= MUX_s_1_2_2((NOT and_757_cse), or_tmp_104, fsm_output(5));
  mux_3686_nl <= MUX_s_1_2_2(mux_3685_nl, or_361_cse, fsm_output(7));
  mux_3688_nl <= MUX_s_1_2_2(mux_3687_nl, mux_3686_nl, and_526_cse);
  mux_3693_nl <= MUX_s_1_2_2(mux_3692_nl, mux_3688_nl, fsm_output(2));
  mux_3694_nl <= MUX_s_1_2_2(mux_tmp_3691, mux_3693_nl, fsm_output(4));
  mux_3682_nl <= MUX_s_1_2_2(mux_tmp_3681, mux_tmp_3679, and_526_cse);
  nor_527_nl <= NOT((fsm_output(0)) OR (NOT (fsm_output(7))));
  mux_3678_nl <= MUX_s_1_2_2(mux_tmp_215, nand_tmp_7, nor_527_nl);
  mux_3680_nl <= MUX_s_1_2_2(mux_tmp_3679, mux_3678_nl, fsm_output(1));
  mux_3683_nl <= MUX_s_1_2_2(mux_3682_nl, mux_3680_nl, fsm_output(2));
  mux_3676_nl <= MUX_s_1_2_2(mux_tmp_3673, mux_tmp_3674, and_526_cse);
  mux_3675_nl <= MUX_s_1_2_2(mux_tmp_3674, mux_tmp_3673, or_3388_cse);
  mux_3677_nl <= MUX_s_1_2_2(mux_3676_nl, mux_3675_nl, fsm_output(2));
  mux_3684_nl <= MUX_s_1_2_2(mux_3683_nl, mux_3677_nl, fsm_output(4));
  mux_3695_nl <= MUX_s_1_2_2(mux_3694_nl, mux_3684_nl, fsm_output(8));
  mux_3727_nl <= MUX_s_1_2_2(mux_3726_nl, mux_3695_nl, fsm_output(6));
  mux_3766_nl <= MUX_s_1_2_2(mux_3765_nl, mux_3727_nl, fsm_output(3));
  COMP_LOOP_or_28_nl <= and_dcpl_140 OR and_dcpl_197;
  COMP_LOOP_mux1h_480_nl <= MUX1HOT_s_1_6_2(modExp_exp_1_4_1_sva, COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm,
      (COMP_LOOP_k_9_4_sva_4_0(0)), (z_out_6(7)), (z_out_7(6)), (z_out_7(5)), STD_LOGIC_VECTOR'(
      not_tmp_701 & (NOT mux_3766_nl) & not_tmp_688 & COMP_LOOP_or_28_nl & and_dcpl_171
      & and_dcpl_226));
  or_3396_nl <= (fsm_output(5)) OR (fsm_output(7)) OR (fsm_output(9)) OR (fsm_output(10));
  nand_175_nl <= NOT((fsm_output(0)) AND (fsm_output(5)) AND (fsm_output(7)) AND
      (fsm_output(9)) AND (fsm_output(10)));
  mux_2449_nl <= MUX_s_1_2_2(or_3396_nl, nand_175_nl, fsm_output(1));
  mux_2450_nl <= MUX_s_1_2_2(mux_2449_nl, nand_356_cse, or_491_cse);
  mux_2451_nl <= MUX_s_1_2_2(mux_2450_nl, nand_357_cse, fsm_output(6));
  mux_2452_nl <= MUX_s_1_2_2(mux_2451_nl, nand_358_cse, fsm_output(8));
  or_3549_nl <= (fsm_output(2)) OR (NOT (fsm_output(0))) OR (fsm_output(1)) OR (fsm_output(9))
      OR (fsm_output(10));
  mux_3885_nl <= MUX_s_1_2_2(or_3549_nl, mux_tmp_3864, fsm_output(3));
  nor_1705_nl <= NOT((fsm_output(6)) OR (NOT mux_3885_nl));
  nor_1706_nl <= NOT(CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT and_757_cse));
  and_1165_nl <= (fsm_output(2)) AND (NOT or_tmp_3347);
  mux_3883_nl <= MUX_s_1_2_2(nor_1706_nl, and_1165_nl, fsm_output(3));
  and_1166_nl <= CONV_SL_1_1(fsm_output(3 DOWNTO 2)=STD_LOGIC_VECTOR'("11")) AND
      (NOT or_tmp_3352);
  mux_3884_nl <= MUX_s_1_2_2(mux_3883_nl, and_1166_nl, fsm_output(6));
  mux_3886_nl <= MUX_s_1_2_2(nor_1705_nl, mux_3884_nl, fsm_output(4));
  or_3619_nl <= CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00")) OR (NOT
      nor_tmp_552);
  or_3543_nl <= CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR (NOT
      and_757_cse);
  mux_3880_nl <= MUX_s_1_2_2((NOT nor_tmp_554), or_3543_nl, fsm_output(2));
  or_3620_nl <= (fsm_output(3)) OR mux_3880_nl;
  mux_3881_nl <= MUX_s_1_2_2(or_3619_nl, or_3620_nl, fsm_output(6));
  or_3541_nl <= (NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))))
      OR CONV_SL_1_1(fsm_output(10 DOWNTO 9)/=STD_LOGIC_VECTOR'("00"));
  mux_3877_nl <= MUX_s_1_2_2(or_3541_nl, or_tmp_3339, fsm_output(2));
  mux_3878_nl <= MUX_s_1_2_2(mux_3877_nl, (NOT or_tmp_3357), fsm_output(3));
  nor_1708_nl <= NOT(CONV_SL_1_1(fsm_output(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (NOT and_757_cse));
  mux_3876_nl <= MUX_s_1_2_2(mux_tmp_3856, nor_1708_nl, fsm_output(3));
  mux_3879_nl <= MUX_s_1_2_2(mux_3878_nl, mux_3876_nl, fsm_output(6));
  mux_3882_nl <= MUX_s_1_2_2(mux_3881_nl, mux_3879_nl, fsm_output(4));
  mux_3887_nl <= MUX_s_1_2_2(mux_3886_nl, mux_3882_nl, fsm_output(5));
  or_3537_nl <= (NOT (fsm_output(1))) OR (fsm_output(9)) OR (fsm_output(10));
  mux_3871_nl <= MUX_s_1_2_2(or_3537_nl, or_tmp_3339, fsm_output(2));
  mux_3872_nl <= MUX_s_1_2_2((NOT mux_3871_nl), or_tmp_3357, fsm_output(3));
  mux_3868_nl <= MUX_s_1_2_2(and_757_cse, mux_tmp_227, and_526_cse);
  mux_3869_nl <= MUX_s_1_2_2(mux_3868_nl, mux_tmp_3830, fsm_output(2));
  or_3534_nl <= (fsm_output(2)) OR (fsm_output(0)) OR (fsm_output(1)) OR (fsm_output(9))
      OR (NOT (fsm_output(10)));
  mux_3870_nl <= MUX_s_1_2_2(mux_3869_nl, or_3534_nl, fsm_output(3));
  mux_3873_nl <= MUX_s_1_2_2(mux_3872_nl, mux_3870_nl, fsm_output(6));
  nand_417_nl <= NOT((fsm_output(3)) AND (NOT mux_tmp_3864));
  mux_3867_nl <= MUX_s_1_2_2(nand_417_nl, mux_tmp_3848, fsm_output(6));
  mux_3874_nl <= MUX_s_1_2_2(mux_3873_nl, mux_3867_nl, fsm_output(4));
  and_1168_nl <= (fsm_output(6)) AND (fsm_output(3));
  mux_3864_nl <= MUX_s_1_2_2(and_757_cse, mux_tmp_3841, and_1168_nl);
  mux_3865_nl <= MUX_s_1_2_2(mux_3864_nl, or_3532_cse, fsm_output(4));
  mux_3875_nl <= MUX_s_1_2_2(mux_3874_nl, mux_3865_nl, fsm_output(5));
  mux_3888_nl <= MUX_s_1_2_2(mux_3887_nl, mux_3875_nl, fsm_output(7));
  mux_3859_nl <= MUX_s_1_2_2(mux_tmp_3856, and_757_cse, fsm_output(3));
  mux_3860_nl <= MUX_s_1_2_2(mux_3859_nl, mux_tmp_3839, fsm_output(6));
  or_3529_nl <= (fsm_output(3)) OR mux_tmp_3828;
  mux_3857_nl <= MUX_s_1_2_2(and_757_cse, or_3529_nl, fsm_output(6));
  mux_3861_nl <= MUX_s_1_2_2(mux_3860_nl, mux_3857_nl, fsm_output(4));
  mux_3852_nl <= MUX_s_1_2_2(and_757_cse, mux_tmp_227, fsm_output(1));
  mux_3851_nl <= MUX_s_1_2_2(mux_tmp_227, or_tmp_104, or_3388_cse);
  mux_3853_nl <= MUX_s_1_2_2(mux_3852_nl, mux_3851_nl, fsm_output(2));
  mux_3854_nl <= MUX_s_1_2_2(and_757_cse, mux_3853_nl, fsm_output(3));
  mux_3855_nl <= MUX_s_1_2_2(mux_3854_nl, mux_tmp_3848, fsm_output(6));
  mux_3848_nl <= MUX_s_1_2_2(or_tmp_3344, and_757_cse, fsm_output(6));
  mux_3856_nl <= MUX_s_1_2_2(mux_3855_nl, mux_3848_nl, fsm_output(4));
  mux_3862_nl <= MUX_s_1_2_2(mux_3861_nl, mux_3856_nl, fsm_output(5));
  mux_3845_nl <= MUX_s_1_2_2(and_757_cse, or_tmp_3344, fsm_output(6));
  or_3522_nl <= (fsm_output(3)) OR mux_tmp_3841;
  mux_3844_nl <= MUX_s_1_2_2(or_3522_nl, mux_tmp_3839, fsm_output(6));
  mux_3846_nl <= MUX_s_1_2_2(mux_3845_nl, mux_3844_nl, fsm_output(4));
  nand_416_nl <= NOT((fsm_output(2)) AND (NOT or_tmp_3337));
  mux_3837_nl <= MUX_s_1_2_2(nor_tmp_549, and_757_cse, fsm_output(2));
  mux_3838_nl <= MUX_s_1_2_2(nand_416_nl, mux_3837_nl, fsm_output(3));
  mux_3839_nl <= MUX_s_1_2_2(mux_3838_nl, and_757_cse, fsm_output(6));
  mux_3834_nl <= MUX_s_1_2_2(and_757_cse, mux_tmp_227, and_536_cse);
  or_3513_nl <= (fsm_output(0)) OR (fsm_output(1)) OR (fsm_output(9)) OR (NOT (fsm_output(10)));
  mux_3833_nl <= MUX_s_1_2_2(mux_tmp_3830, or_3513_nl, fsm_output(2));
  mux_3835_nl <= MUX_s_1_2_2(mux_3834_nl, mux_3833_nl, fsm_output(3));
  mux_3831_nl <= MUX_s_1_2_2(and_757_cse, mux_tmp_3828, fsm_output(3));
  mux_3836_nl <= MUX_s_1_2_2(mux_3835_nl, mux_3831_nl, fsm_output(6));
  mux_3840_nl <= MUX_s_1_2_2(mux_3839_nl, mux_3836_nl, fsm_output(4));
  mux_3847_nl <= MUX_s_1_2_2(mux_3846_nl, mux_3840_nl, fsm_output(5));
  mux_3863_nl <= MUX_s_1_2_2(mux_3862_nl, mux_3847_nl, fsm_output(7));
  mux_3889_nl <= MUX_s_1_2_2(mux_3888_nl, mux_3863_nl, fsm_output(8));
  or_3612_nl <= (NOT (fsm_output(1))) OR (fsm_output(10)) OR (NOT COMP_LOOP_nor_11_itm)
      OR (NOT (fsm_output(6))) OR (NOT (fsm_output(2))) OR (fsm_output(9));
  or_3611_nl <= (fsm_output(1)) OR (fsm_output(10)) OR (fsm_output(6)) OR (fsm_output(2))
      OR (fsm_output(9));
  mux_3938_nl <= MUX_s_1_2_2(or_3612_nl, or_3611_nl, fsm_output(0));
  mux_3936_nl <= MUX_s_1_2_2(or_tmp_3409, or_2965_cse, fsm_output(1));
  mux_3937_nl <= MUX_s_1_2_2(mux_3936_nl, mux_3935_cse, fsm_output(0));
  mux_3939_nl <= MUX_s_1_2_2(mux_3938_nl, mux_3937_nl, fsm_output(3));
  or_3608_nl <= (fsm_output(3)) OR (fsm_output(0)) OR (NOT (fsm_output(1))) OR (NOT
      (fsm_output(10))) OR (NOT COMP_LOOP_nor_11_itm) OR (NOT (fsm_output(6))) OR
      (fsm_output(2)) OR (NOT (fsm_output(9)));
  mux_3940_nl <= MUX_s_1_2_2(mux_3939_nl, or_3608_nl, fsm_output(5));
  or_3606_nl <= (fsm_output(0)) OR (NOT (fsm_output(1))) OR (NOT (fsm_output(10)))
      OR (fsm_output(6)) OR (fsm_output(2)) OR (NOT (fsm_output(9)));
  or_3604_nl <= (fsm_output(1)) OR (fsm_output(10)) OR not_tmp_882;
  nand_423_nl <= NOT((fsm_output(1)) AND (fsm_output(10)) AND COMP_LOOP_nor_11_itm
      AND (fsm_output(6)) AND (fsm_output(2)) AND (NOT (fsm_output(9))));
  mux_3932_nl <= MUX_s_1_2_2(or_3604_nl, nand_423_nl, fsm_output(0));
  mux_3933_nl <= MUX_s_1_2_2(or_3606_nl, mux_3932_nl, fsm_output(3));
  or_3601_nl <= (fsm_output(10)) OR (fsm_output(2)) OR (fsm_output(9));
  mux_3929_nl <= MUX_s_1_2_2(or_3601_nl, mux_tmp_3906, fsm_output(1));
  mux_3925_nl <= MUX_s_1_2_2((fsm_output(9)), (NOT (fsm_output(9))), fsm_output(2));
  mux_3926_nl <= MUX_s_1_2_2(mux_3925_nl, or_2855_cse, fsm_output(6));
  mux_3927_nl <= MUX_s_1_2_2(or_tmp_3402, mux_3926_nl, COMP_LOOP_nor_11_itm);
  or_3600_nl <= (fsm_output(10)) OR mux_3927_nl;
  mux_3928_nl <= MUX_s_1_2_2(or_tmp_3409, or_3600_nl, fsm_output(1));
  mux_3930_nl <= MUX_s_1_2_2(mux_3929_nl, mux_3928_nl, fsm_output(0));
  or_3599_nl <= (NOT (fsm_output(10))) OR (fsm_output(6)) OR (fsm_output(2)) OR (fsm_output(9));
  or_3598_nl <= (NOT (fsm_output(10))) OR (NOT COMP_LOOP_nor_11_itm) OR (fsm_output(6))
      OR (fsm_output(2)) OR (fsm_output(9));
  mux_3923_nl <= MUX_s_1_2_2(or_3599_nl, or_3598_nl, fsm_output(1));
  nand_420_nl <= NOT((fsm_output(10)) AND (NOT mux_tmp_3903));
  or_3597_nl <= (NOT (fsm_output(10))) OR (fsm_output(6)) OR (fsm_output(2)) OR (NOT
      (fsm_output(9)));
  mux_3922_nl <= MUX_s_1_2_2(nand_420_nl, or_3597_nl, fsm_output(1));
  mux_3924_nl <= MUX_s_1_2_2(mux_3923_nl, mux_3922_nl, fsm_output(0));
  mux_3931_nl <= MUX_s_1_2_2(mux_3930_nl, mux_3924_nl, fsm_output(3));
  mux_3934_nl <= MUX_s_1_2_2(mux_3933_nl, mux_3931_nl, fsm_output(5));
  mux_3941_nl <= MUX_s_1_2_2(mux_3940_nl, mux_3934_nl, fsm_output(4));
  or_3594_nl <= (fsm_output(10)) OR (NOT COMP_LOOP_nor_11_itm) OR (NOT (fsm_output(6)))
      OR (fsm_output(2)) OR (fsm_output(9));
  mux_3918_nl <= MUX_s_1_2_2(or_3594_nl, or_tmp_3382, fsm_output(1));
  or_3593_nl <= (NOT (fsm_output(1))) OR (fsm_output(10)) OR (NOT COMP_LOOP_nor_11_itm)
      OR (NOT (fsm_output(6))) OR (fsm_output(2)) OR (NOT (fsm_output(9)));
  mux_3919_nl <= MUX_s_1_2_2(mux_3918_nl, or_3593_nl, fsm_output(0));
  or_3595_nl <= (fsm_output(3)) OR mux_3919_nl;
  or_3591_nl <= (fsm_output(3)) OR (NOT (fsm_output(0))) OR (fsm_output(1)) OR (NOT
      (fsm_output(10))) OR (NOT COMP_LOOP_nor_11_itm) OR (fsm_output(6)) OR (fsm_output(2))
      OR (fsm_output(9));
  mux_3920_nl <= MUX_s_1_2_2(or_3595_nl, or_3591_nl, fsm_output(5));
  or_3589_nl <= (NOT (fsm_output(0))) OR (NOT (fsm_output(1))) OR (fsm_output(10))
      OR (NOT (fsm_output(6))) OR (NOT (fsm_output(2))) OR (fsm_output(9));
  mux_3915_nl <= MUX_s_1_2_2(or_tmp_3409, or_tmp_3403, fsm_output(1));
  mux_3916_nl <= MUX_s_1_2_2(mux_3915_nl, mux_tmp_3907, fsm_output(0));
  mux_3917_nl <= MUX_s_1_2_2(or_3589_nl, mux_3916_nl, fsm_output(3));
  or_3590_nl <= (fsm_output(5)) OR mux_3917_nl;
  mux_3921_nl <= MUX_s_1_2_2(mux_3920_nl, or_3590_nl, fsm_output(4));
  mux_3942_nl <= MUX_s_1_2_2(mux_3941_nl, mux_3921_nl, fsm_output(7));
  or_3578_nl <= (fsm_output(10)) OR (fsm_output(6)) OR (fsm_output(2)) OR (NOT (fsm_output(9)));
  mux_3906_nl <= MUX_s_1_2_2(or_tmp_3403, or_3578_nl, fsm_output(1));
  mux_3910_nl <= MUX_s_1_2_2(mux_tmp_3907, mux_3906_nl, fsm_output(0));
  or_3576_nl <= (fsm_output(0)) OR (fsm_output(1)) OR (NOT (fsm_output(10))) OR (NOT
      COMP_LOOP_nor_11_itm) OR (fsm_output(6)) OR (fsm_output(2)) OR (fsm_output(9));
  mux_3911_nl <= MUX_s_1_2_2(mux_3910_nl, or_3576_nl, fsm_output(3));
  or_3575_nl <= (NOT (fsm_output(0))) OR (NOT (fsm_output(1))) OR (fsm_output(10))
      OR or_tmp_3384;
  or_3573_nl <= (fsm_output(10)) OR not_tmp_882;
  mux_3901_nl <= MUX_s_1_2_2(or_3573_nl, or_tmp_3381, fsm_output(1));
  mux_3902_nl <= MUX_s_1_2_2(mux_3901_nl, mux_tmp_3892, fsm_output(0));
  mux_3903_nl <= MUX_s_1_2_2(or_3575_nl, mux_3902_nl, fsm_output(3));
  mux_3912_nl <= MUX_s_1_2_2(mux_3911_nl, mux_3903_nl, fsm_output(5));
  or_3572_nl <= (NOT (fsm_output(5))) OR (NOT (fsm_output(3))) OR (fsm_output(0))
      OR (NOT (fsm_output(1))) OR (fsm_output(10)) OR (fsm_output(6)) OR (NOT (fsm_output(2)))
      OR (fsm_output(9));
  mux_3913_nl <= MUX_s_1_2_2(mux_3912_nl, or_3572_nl, fsm_output(4));
  or_3571_nl <= (NOT (fsm_output(3))) OR (fsm_output(0)) OR (NOT (fsm_output(1)))
      OR (fsm_output(10)) OR or_tmp_3384;
  or_3569_nl <= (NOT (fsm_output(0))) OR (fsm_output(1)) OR (fsm_output(10)) OR (fsm_output(6))
      OR (NOT (fsm_output(2))) OR (fsm_output(9));
  or_3568_nl <= (fsm_output(1)) OR (fsm_output(10)) OR (fsm_output(6)) OR (fsm_output(2))
      OR (NOT (fsm_output(9)));
  mux_3897_nl <= MUX_s_1_2_2(or_3568_nl, or_2914_cse, fsm_output(0));
  mux_3898_nl <= MUX_s_1_2_2(or_3569_nl, mux_3897_nl, fsm_output(3));
  mux_3899_nl <= MUX_s_1_2_2(or_3571_nl, mux_3898_nl, fsm_output(5));
  or_3556_nl <= (fsm_output(10)) OR (NOT COMP_LOOP_nor_11_itm) OR (NOT (fsm_output(6)))
      OR (fsm_output(2)) OR (NOT (fsm_output(9)));
  mux_3892_nl <= MUX_s_1_2_2(or_tmp_3381, or_3556_nl, fsm_output(1));
  mux_3895_nl <= MUX_s_1_2_2(mux_tmp_3892, mux_3892_nl, fsm_output(0));
  or_3565_nl <= (fsm_output(3)) OR mux_3895_nl;
  or_3554_nl <= (NOT (fsm_output(0))) OR (fsm_output(1)) OR (fsm_output(10)) OR (NOT
      COMP_LOOP_nor_11_itm) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(2))) OR
      (fsm_output(9));
  or_3553_nl <= (fsm_output(1)) OR (fsm_output(10)) OR (NOT COMP_LOOP_nor_11_itm)
      OR (NOT (fsm_output(6))) OR (fsm_output(2)) OR (NOT (fsm_output(9)));
  or_3551_nl <= (NOT (fsm_output(1))) OR (NOT (fsm_output(10))) OR (NOT COMP_LOOP_nor_11_itm)
      OR (NOT (fsm_output(6))) OR (fsm_output(2)) OR (fsm_output(9));
  mux_3890_nl <= MUX_s_1_2_2(or_3553_nl, or_3551_nl, fsm_output(0));
  mux_3891_nl <= MUX_s_1_2_2(or_3554_nl, mux_3890_nl, fsm_output(3));
  mux_3896_nl <= MUX_s_1_2_2(or_3565_nl, mux_3891_nl, fsm_output(5));
  mux_3900_nl <= MUX_s_1_2_2(mux_3899_nl, mux_3896_nl, fsm_output(4));
  mux_3914_nl <= MUX_s_1_2_2(mux_3913_nl, mux_3900_nl, fsm_output(7));
  mux_3943_nl <= MUX_s_1_2_2(mux_3942_nl, mux_3914_nl, fsm_output(8));
  or_2641_nl <= (fsm_output(1)) OR (NOT (fsm_output(4))) OR (fsm_output(7)) OR (NOT
      (fsm_output(5))) OR (fsm_output(3));
  or_2640_nl <= (fsm_output(1)) OR (fsm_output(4)) OR (fsm_output(7)) OR (fsm_output(5))
      OR (NOT (fsm_output(3)));
  mux_2638_nl <= MUX_s_1_2_2(or_2641_nl, or_2640_nl, fsm_output(0));
  or_2642_nl <= (fsm_output(9)) OR mux_2638_nl;
  or_2638_nl <= (NOT (fsm_output(9))) OR (fsm_output(0)) OR (NOT (fsm_output(1)))
      OR (fsm_output(4)) OR (NOT (fsm_output(7))) OR (NOT (fsm_output(5))) OR (fsm_output(3));
  mux_2639_nl <= MUX_s_1_2_2(or_2642_nl, or_2638_nl, fsm_output(10));
  or_3508_nl <= mux_2639_nl OR (fsm_output(2)) OR (fsm_output(8)) OR (fsm_output(6));
  nor_1700_nl <= NOT((NOT (fsm_output(3))) OR (fsm_output(4)) OR (NOT (fsm_output(0)))
      OR (fsm_output(6)) OR (fsm_output(7)) OR (fsm_output(10)) OR (fsm_output(9))
      OR (fsm_output(1)));
  or_3616_nl <= (fsm_output(6)) OR (NOT((fsm_output(7)) AND (fsm_output(10)) AND
      (fsm_output(9)) AND (fsm_output(1))));
  or_3615_nl <= (NOT (fsm_output(6))) OR (fsm_output(7)) OR (NOT((fsm_output(10))
      AND (fsm_output(9)) AND (fsm_output(1))));
  mux_3944_nl <= MUX_s_1_2_2(or_3616_nl, or_3615_nl, fsm_output(0));
  or_3613_nl <= (fsm_output(0)) OR (fsm_output(6)) OR (fsm_output(7)) OR (fsm_output(10))
      OR (fsm_output(9)) OR (fsm_output(1));
  mux_3945_nl <= MUX_s_1_2_2(mux_3944_nl, or_3613_nl, fsm_output(4));
  nor_1701_nl <= NOT((fsm_output(3)) OR mux_3945_nl);
  mux_3946_nl <= MUX_s_1_2_2(nor_1700_nl, nor_1701_nl, fsm_output(5));
  nor_690_nl <= NOT((fsm_output(5)) OR (fsm_output(7)) OR (fsm_output(9)) OR (fsm_output(10)));
  mux_2663_nl <= MUX_s_1_2_2(nor_690_nl, mux_tmp_2659, and_526_cse);
  mux_2662_nl <= MUX_s_1_2_2(mux_tmp_2659, and_465_cse, fsm_output(1));
  mux_2664_nl <= MUX_s_1_2_2(mux_2663_nl, mux_2662_nl, fsm_output(3));
  mux_2661_nl <= MUX_s_1_2_2(mux_tmp_2659, and_465_cse, fsm_output(3));
  mux_2665_nl <= MUX_s_1_2_2(mux_2664_nl, mux_2661_nl, fsm_output(2));
  nand_170_nl <= NOT(CONV_SL_1_1(fsm_output(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1101")));
  mux_2660_nl <= MUX_s_1_2_2(mux_tmp_2659, and_465_cse, nand_170_nl);
  mux_2666_nl <= MUX_s_1_2_2(mux_2665_nl, mux_2660_nl, fsm_output(4));
  mux_2667_nl <= MUX_s_1_2_2(mux_2666_nl, and_756_cse, fsm_output(6));
  mux_2668_nl <= MUX_s_1_2_2(mux_2667_nl, and_757_cse, fsm_output(8));
  COMP_LOOP_or_8_nl <= (COMP_LOOP_COMP_LOOP_nor_itm AND and_dcpl_257) OR (COMP_LOOP_COMP_LOOP_and_14_itm
      AND and_279_m1c) OR (COMP_LOOP_COMP_LOOP_and_13_itm AND and_281_m1c) OR (COMP_LOOP_COMP_LOOP_and_12_itm
      AND and_284_m1c) OR (COMP_LOOP_COMP_LOOP_and_11_itm AND and_286_m1c) OR (COMP_LOOP_COMP_LOOP_and_10_itm
      AND and_288_m1c) OR (COMP_LOOP_COMP_LOOP_and_9_itm AND and_291_m1c) OR (COMP_LOOP_COMP_LOOP_and_8_itm
      AND and_292_m1c) OR (COMP_LOOP_COMP_LOOP_and_68_itm AND and_295_m1c) OR (COMP_LOOP_COMP_LOOP_and_6_itm
      AND and_297_m1c) OR (COMP_LOOP_COMP_LOOP_and_5_itm AND and_299_m1c) OR (COMP_LOOP_COMP_LOOP_and_4_itm
      AND and_302_m1c) OR (COMP_LOOP_COMP_LOOP_and_64_itm AND and_304_m1c) OR (COMP_LOOP_COMP_LOOP_and_2_itm
      AND and_307_m1c) OR (COMP_LOOP_COMP_LOOP_and_62_itm AND and_309_m1c) OR (COMP_LOOP_COMP_LOOP_and_305_itm
      AND and_311_m1c);
  COMP_LOOP_or_9_nl <= (COMP_LOOP_COMP_LOOP_and_305_itm AND and_dcpl_257) OR (COMP_LOOP_COMP_LOOP_nor_itm
      AND and_279_m1c) OR (COMP_LOOP_COMP_LOOP_and_14_itm AND and_281_m1c) OR (COMP_LOOP_COMP_LOOP_and_13_itm
      AND and_284_m1c) OR (COMP_LOOP_COMP_LOOP_and_12_itm AND and_286_m1c) OR (COMP_LOOP_COMP_LOOP_and_11_itm
      AND and_288_m1c) OR (COMP_LOOP_COMP_LOOP_and_10_itm AND and_291_m1c) OR (COMP_LOOP_COMP_LOOP_and_9_itm
      AND and_292_m1c) OR (COMP_LOOP_COMP_LOOP_and_8_itm AND and_295_m1c) OR (COMP_LOOP_COMP_LOOP_and_68_itm
      AND and_297_m1c) OR (COMP_LOOP_COMP_LOOP_and_6_itm AND and_299_m1c) OR (COMP_LOOP_COMP_LOOP_and_5_itm
      AND and_302_m1c) OR (COMP_LOOP_COMP_LOOP_and_4_itm AND and_304_m1c) OR (COMP_LOOP_COMP_LOOP_and_64_itm
      AND and_307_m1c) OR (COMP_LOOP_COMP_LOOP_and_2_itm AND and_309_m1c) OR (COMP_LOOP_COMP_LOOP_and_62_itm
      AND and_311_m1c);
  COMP_LOOP_or_10_nl <= (COMP_LOOP_COMP_LOOP_and_62_itm AND and_dcpl_257) OR (COMP_LOOP_COMP_LOOP_and_305_itm
      AND and_279_m1c) OR (COMP_LOOP_COMP_LOOP_nor_itm AND and_281_m1c) OR (COMP_LOOP_COMP_LOOP_and_14_itm
      AND and_284_m1c) OR (COMP_LOOP_COMP_LOOP_and_13_itm AND and_286_m1c) OR (COMP_LOOP_COMP_LOOP_and_12_itm
      AND and_288_m1c) OR (COMP_LOOP_COMP_LOOP_and_11_itm AND and_291_m1c) OR (COMP_LOOP_COMP_LOOP_and_10_itm
      AND and_292_m1c) OR (COMP_LOOP_COMP_LOOP_and_9_itm AND and_295_m1c) OR (COMP_LOOP_COMP_LOOP_and_8_itm
      AND and_297_m1c) OR (COMP_LOOP_COMP_LOOP_and_68_itm AND and_299_m1c) OR (COMP_LOOP_COMP_LOOP_and_6_itm
      AND and_302_m1c) OR (COMP_LOOP_COMP_LOOP_and_5_itm AND and_304_m1c) OR (COMP_LOOP_COMP_LOOP_and_4_itm
      AND and_307_m1c) OR (COMP_LOOP_COMP_LOOP_and_64_itm AND and_309_m1c) OR (COMP_LOOP_COMP_LOOP_and_2_itm
      AND and_311_m1c);
  COMP_LOOP_or_11_nl <= (COMP_LOOP_COMP_LOOP_and_2_itm AND and_dcpl_257) OR (COMP_LOOP_COMP_LOOP_and_62_itm
      AND and_279_m1c) OR (COMP_LOOP_COMP_LOOP_and_305_itm AND and_281_m1c) OR (COMP_LOOP_COMP_LOOP_nor_itm
      AND and_284_m1c) OR (COMP_LOOP_COMP_LOOP_and_14_itm AND and_286_m1c) OR (COMP_LOOP_COMP_LOOP_and_13_itm
      AND and_288_m1c) OR (COMP_LOOP_COMP_LOOP_and_12_itm AND and_291_m1c) OR (COMP_LOOP_COMP_LOOP_and_11_itm
      AND and_292_m1c) OR (COMP_LOOP_COMP_LOOP_and_10_itm AND and_295_m1c) OR (COMP_LOOP_COMP_LOOP_and_9_itm
      AND and_297_m1c) OR (COMP_LOOP_COMP_LOOP_and_8_itm AND and_299_m1c) OR (COMP_LOOP_COMP_LOOP_and_68_itm
      AND and_302_m1c) OR (COMP_LOOP_COMP_LOOP_and_6_itm AND and_304_m1c) OR (COMP_LOOP_COMP_LOOP_and_5_itm
      AND and_307_m1c) OR (COMP_LOOP_COMP_LOOP_and_4_itm AND and_309_m1c) OR (COMP_LOOP_COMP_LOOP_and_64_itm
      AND and_311_m1c);
  COMP_LOOP_or_12_nl <= (COMP_LOOP_COMP_LOOP_and_64_itm AND and_dcpl_257) OR (COMP_LOOP_COMP_LOOP_and_2_itm
      AND and_279_m1c) OR (COMP_LOOP_COMP_LOOP_and_62_itm AND and_281_m1c) OR (COMP_LOOP_COMP_LOOP_and_305_itm
      AND and_284_m1c) OR (COMP_LOOP_COMP_LOOP_nor_itm AND and_286_m1c) OR (COMP_LOOP_COMP_LOOP_and_14_itm
      AND and_288_m1c) OR (COMP_LOOP_COMP_LOOP_and_13_itm AND and_291_m1c) OR (COMP_LOOP_COMP_LOOP_and_12_itm
      AND and_292_m1c) OR (COMP_LOOP_COMP_LOOP_and_11_itm AND and_295_m1c) OR (COMP_LOOP_COMP_LOOP_and_10_itm
      AND and_297_m1c) OR (COMP_LOOP_COMP_LOOP_and_9_itm AND and_299_m1c) OR (COMP_LOOP_COMP_LOOP_and_8_itm
      AND and_302_m1c) OR (COMP_LOOP_COMP_LOOP_and_68_itm AND and_304_m1c) OR (COMP_LOOP_COMP_LOOP_and_6_itm
      AND and_307_m1c) OR (COMP_LOOP_COMP_LOOP_and_5_itm AND and_309_m1c) OR (COMP_LOOP_COMP_LOOP_and_4_itm
      AND and_311_m1c);
  COMP_LOOP_or_13_nl <= (COMP_LOOP_COMP_LOOP_and_4_itm AND and_dcpl_257) OR (COMP_LOOP_COMP_LOOP_and_64_itm
      AND and_279_m1c) OR (COMP_LOOP_COMP_LOOP_and_2_itm AND and_281_m1c) OR (COMP_LOOP_COMP_LOOP_and_62_itm
      AND and_284_m1c) OR (COMP_LOOP_COMP_LOOP_and_305_itm AND and_286_m1c) OR (COMP_LOOP_COMP_LOOP_nor_itm
      AND and_288_m1c) OR (COMP_LOOP_COMP_LOOP_and_14_itm AND and_291_m1c) OR (COMP_LOOP_COMP_LOOP_and_13_itm
      AND and_292_m1c) OR (COMP_LOOP_COMP_LOOP_and_12_itm AND and_295_m1c) OR (COMP_LOOP_COMP_LOOP_and_11_itm
      AND and_297_m1c) OR (COMP_LOOP_COMP_LOOP_and_10_itm AND and_299_m1c) OR (COMP_LOOP_COMP_LOOP_and_9_itm
      AND and_302_m1c) OR (COMP_LOOP_COMP_LOOP_and_8_itm AND and_304_m1c) OR (COMP_LOOP_COMP_LOOP_and_68_itm
      AND and_307_m1c) OR (COMP_LOOP_COMP_LOOP_and_6_itm AND and_309_m1c) OR (COMP_LOOP_COMP_LOOP_and_5_itm
      AND and_311_m1c);
  COMP_LOOP_or_14_nl <= (COMP_LOOP_COMP_LOOP_and_5_itm AND and_dcpl_257) OR (COMP_LOOP_COMP_LOOP_and_4_itm
      AND and_279_m1c) OR (COMP_LOOP_COMP_LOOP_and_64_itm AND and_281_m1c) OR (COMP_LOOP_COMP_LOOP_and_2_itm
      AND and_284_m1c) OR (COMP_LOOP_COMP_LOOP_and_62_itm AND and_286_m1c) OR (COMP_LOOP_COMP_LOOP_and_305_itm
      AND and_288_m1c) OR (COMP_LOOP_COMP_LOOP_nor_itm AND and_291_m1c) OR (COMP_LOOP_COMP_LOOP_and_14_itm
      AND and_292_m1c) OR (COMP_LOOP_COMP_LOOP_and_13_itm AND and_295_m1c) OR (COMP_LOOP_COMP_LOOP_and_12_itm
      AND and_297_m1c) OR (COMP_LOOP_COMP_LOOP_and_11_itm AND and_299_m1c) OR (COMP_LOOP_COMP_LOOP_and_10_itm
      AND and_302_m1c) OR (COMP_LOOP_COMP_LOOP_and_9_itm AND and_304_m1c) OR (COMP_LOOP_COMP_LOOP_and_8_itm
      AND and_307_m1c) OR (COMP_LOOP_COMP_LOOP_and_68_itm AND and_309_m1c) OR (COMP_LOOP_COMP_LOOP_and_6_itm
      AND and_311_m1c);
  COMP_LOOP_or_15_nl <= (COMP_LOOP_COMP_LOOP_and_6_itm AND and_dcpl_257) OR (COMP_LOOP_COMP_LOOP_and_5_itm
      AND and_279_m1c) OR (COMP_LOOP_COMP_LOOP_and_4_itm AND and_281_m1c) OR (COMP_LOOP_COMP_LOOP_and_64_itm
      AND and_284_m1c) OR (COMP_LOOP_COMP_LOOP_and_2_itm AND and_286_m1c) OR (COMP_LOOP_COMP_LOOP_and_62_itm
      AND and_288_m1c) OR (COMP_LOOP_COMP_LOOP_and_305_itm AND and_291_m1c) OR (COMP_LOOP_COMP_LOOP_nor_itm
      AND and_292_m1c) OR (COMP_LOOP_COMP_LOOP_and_14_itm AND and_295_m1c) OR (COMP_LOOP_COMP_LOOP_and_13_itm
      AND and_297_m1c) OR (COMP_LOOP_COMP_LOOP_and_12_itm AND and_299_m1c) OR (COMP_LOOP_COMP_LOOP_and_11_itm
      AND and_302_m1c) OR (COMP_LOOP_COMP_LOOP_and_10_itm AND and_304_m1c) OR (COMP_LOOP_COMP_LOOP_and_9_itm
      AND and_307_m1c) OR (COMP_LOOP_COMP_LOOP_and_8_itm AND and_309_m1c) OR (COMP_LOOP_COMP_LOOP_and_68_itm
      AND and_311_m1c);
  COMP_LOOP_or_16_nl <= (COMP_LOOP_COMP_LOOP_and_68_itm AND and_dcpl_257) OR (COMP_LOOP_COMP_LOOP_and_6_itm
      AND and_279_m1c) OR (COMP_LOOP_COMP_LOOP_and_5_itm AND and_281_m1c) OR (COMP_LOOP_COMP_LOOP_and_4_itm
      AND and_284_m1c) OR (COMP_LOOP_COMP_LOOP_and_64_itm AND and_286_m1c) OR (COMP_LOOP_COMP_LOOP_and_2_itm
      AND and_288_m1c) OR (COMP_LOOP_COMP_LOOP_and_62_itm AND and_291_m1c) OR (COMP_LOOP_COMP_LOOP_and_305_itm
      AND and_292_m1c) OR (COMP_LOOP_COMP_LOOP_nor_itm AND and_295_m1c) OR (COMP_LOOP_COMP_LOOP_and_14_itm
      AND and_297_m1c) OR (COMP_LOOP_COMP_LOOP_and_13_itm AND and_299_m1c) OR (COMP_LOOP_COMP_LOOP_and_12_itm
      AND and_302_m1c) OR (COMP_LOOP_COMP_LOOP_and_11_itm AND and_304_m1c) OR (COMP_LOOP_COMP_LOOP_and_10_itm
      AND and_307_m1c) OR (COMP_LOOP_COMP_LOOP_and_9_itm AND and_309_m1c) OR (COMP_LOOP_COMP_LOOP_and_8_itm
      AND and_311_m1c);
  COMP_LOOP_or_17_nl <= (COMP_LOOP_COMP_LOOP_and_8_itm AND and_dcpl_257) OR (COMP_LOOP_COMP_LOOP_and_68_itm
      AND and_279_m1c) OR (COMP_LOOP_COMP_LOOP_and_6_itm AND and_281_m1c) OR (COMP_LOOP_COMP_LOOP_and_5_itm
      AND and_284_m1c) OR (COMP_LOOP_COMP_LOOP_and_4_itm AND and_286_m1c) OR (COMP_LOOP_COMP_LOOP_and_64_itm
      AND and_288_m1c) OR (COMP_LOOP_COMP_LOOP_and_2_itm AND and_291_m1c) OR (COMP_LOOP_COMP_LOOP_and_62_itm
      AND and_292_m1c) OR (COMP_LOOP_COMP_LOOP_and_305_itm AND and_295_m1c) OR (COMP_LOOP_COMP_LOOP_nor_itm
      AND and_297_m1c) OR (COMP_LOOP_COMP_LOOP_and_14_itm AND and_299_m1c) OR (COMP_LOOP_COMP_LOOP_and_13_itm
      AND and_302_m1c) OR (COMP_LOOP_COMP_LOOP_and_12_itm AND and_304_m1c) OR (COMP_LOOP_COMP_LOOP_and_11_itm
      AND and_307_m1c) OR (COMP_LOOP_COMP_LOOP_and_10_itm AND and_309_m1c) OR (COMP_LOOP_COMP_LOOP_and_9_itm
      AND and_311_m1c);
  COMP_LOOP_or_18_nl <= (COMP_LOOP_COMP_LOOP_and_9_itm AND and_dcpl_257) OR (COMP_LOOP_COMP_LOOP_and_8_itm
      AND and_279_m1c) OR (COMP_LOOP_COMP_LOOP_and_68_itm AND and_281_m1c) OR (COMP_LOOP_COMP_LOOP_and_6_itm
      AND and_284_m1c) OR (COMP_LOOP_COMP_LOOP_and_5_itm AND and_286_m1c) OR (COMP_LOOP_COMP_LOOP_and_4_itm
      AND and_288_m1c) OR (COMP_LOOP_COMP_LOOP_and_64_itm AND and_291_m1c) OR (COMP_LOOP_COMP_LOOP_and_2_itm
      AND and_292_m1c) OR (COMP_LOOP_COMP_LOOP_and_62_itm AND and_295_m1c) OR (COMP_LOOP_COMP_LOOP_and_305_itm
      AND and_297_m1c) OR (COMP_LOOP_COMP_LOOP_nor_itm AND and_299_m1c) OR (COMP_LOOP_COMP_LOOP_and_14_itm
      AND and_302_m1c) OR (COMP_LOOP_COMP_LOOP_and_13_itm AND and_304_m1c) OR (COMP_LOOP_COMP_LOOP_and_12_itm
      AND and_307_m1c) OR (COMP_LOOP_COMP_LOOP_and_11_itm AND and_309_m1c) OR (COMP_LOOP_COMP_LOOP_and_10_itm
      AND and_311_m1c);
  COMP_LOOP_or_19_nl <= (COMP_LOOP_COMP_LOOP_and_10_itm AND and_dcpl_257) OR (COMP_LOOP_COMP_LOOP_and_9_itm
      AND and_279_m1c) OR (COMP_LOOP_COMP_LOOP_and_8_itm AND and_281_m1c) OR (COMP_LOOP_COMP_LOOP_and_68_itm
      AND and_284_m1c) OR (COMP_LOOP_COMP_LOOP_and_6_itm AND and_286_m1c) OR (COMP_LOOP_COMP_LOOP_and_5_itm
      AND and_288_m1c) OR (COMP_LOOP_COMP_LOOP_and_4_itm AND and_291_m1c) OR (COMP_LOOP_COMP_LOOP_and_64_itm
      AND and_292_m1c) OR (COMP_LOOP_COMP_LOOP_and_2_itm AND and_295_m1c) OR (COMP_LOOP_COMP_LOOP_and_62_itm
      AND and_297_m1c) OR (COMP_LOOP_COMP_LOOP_and_305_itm AND and_299_m1c) OR (COMP_LOOP_COMP_LOOP_nor_itm
      AND and_302_m1c) OR (COMP_LOOP_COMP_LOOP_and_14_itm AND and_304_m1c) OR (COMP_LOOP_COMP_LOOP_and_13_itm
      AND and_307_m1c) OR (COMP_LOOP_COMP_LOOP_and_12_itm AND and_309_m1c) OR (COMP_LOOP_COMP_LOOP_and_11_itm
      AND and_311_m1c);
  COMP_LOOP_or_20_nl <= (COMP_LOOP_COMP_LOOP_and_11_itm AND and_dcpl_257) OR (COMP_LOOP_COMP_LOOP_and_10_itm
      AND and_279_m1c) OR (COMP_LOOP_COMP_LOOP_and_9_itm AND and_281_m1c) OR (COMP_LOOP_COMP_LOOP_and_8_itm
      AND and_284_m1c) OR (COMP_LOOP_COMP_LOOP_and_68_itm AND and_286_m1c) OR (COMP_LOOP_COMP_LOOP_and_6_itm
      AND and_288_m1c) OR (COMP_LOOP_COMP_LOOP_and_5_itm AND and_291_m1c) OR (COMP_LOOP_COMP_LOOP_and_4_itm
      AND and_292_m1c) OR (COMP_LOOP_COMP_LOOP_and_64_itm AND and_295_m1c) OR (COMP_LOOP_COMP_LOOP_and_2_itm
      AND and_297_m1c) OR (COMP_LOOP_COMP_LOOP_and_62_itm AND and_299_m1c) OR (COMP_LOOP_COMP_LOOP_and_305_itm
      AND and_302_m1c) OR (COMP_LOOP_COMP_LOOP_nor_itm AND and_304_m1c) OR (COMP_LOOP_COMP_LOOP_and_14_itm
      AND and_307_m1c) OR (COMP_LOOP_COMP_LOOP_and_13_itm AND and_309_m1c) OR (COMP_LOOP_COMP_LOOP_and_12_itm
      AND and_311_m1c);
  COMP_LOOP_or_21_nl <= (COMP_LOOP_COMP_LOOP_and_12_itm AND and_dcpl_257) OR (COMP_LOOP_COMP_LOOP_and_11_itm
      AND and_279_m1c) OR (COMP_LOOP_COMP_LOOP_and_10_itm AND and_281_m1c) OR (COMP_LOOP_COMP_LOOP_and_9_itm
      AND and_284_m1c) OR (COMP_LOOP_COMP_LOOP_and_8_itm AND and_286_m1c) OR (COMP_LOOP_COMP_LOOP_and_68_itm
      AND and_288_m1c) OR (COMP_LOOP_COMP_LOOP_and_6_itm AND and_291_m1c) OR (COMP_LOOP_COMP_LOOP_and_5_itm
      AND and_292_m1c) OR (COMP_LOOP_COMP_LOOP_and_4_itm AND and_295_m1c) OR (COMP_LOOP_COMP_LOOP_and_64_itm
      AND and_297_m1c) OR (COMP_LOOP_COMP_LOOP_and_2_itm AND and_299_m1c) OR (COMP_LOOP_COMP_LOOP_and_62_itm
      AND and_302_m1c) OR (COMP_LOOP_COMP_LOOP_and_305_itm AND and_304_m1c) OR (COMP_LOOP_COMP_LOOP_nor_itm
      AND and_307_m1c) OR (COMP_LOOP_COMP_LOOP_and_14_itm AND and_309_m1c) OR (COMP_LOOP_COMP_LOOP_and_13_itm
      AND and_311_m1c);
  COMP_LOOP_or_22_nl <= (COMP_LOOP_COMP_LOOP_and_13_itm AND and_dcpl_257) OR (COMP_LOOP_COMP_LOOP_and_12_itm
      AND and_279_m1c) OR (COMP_LOOP_COMP_LOOP_and_11_itm AND and_281_m1c) OR (COMP_LOOP_COMP_LOOP_and_10_itm
      AND and_284_m1c) OR (COMP_LOOP_COMP_LOOP_and_9_itm AND and_286_m1c) OR (COMP_LOOP_COMP_LOOP_and_8_itm
      AND and_288_m1c) OR (COMP_LOOP_COMP_LOOP_and_68_itm AND and_291_m1c) OR (COMP_LOOP_COMP_LOOP_and_6_itm
      AND and_292_m1c) OR (COMP_LOOP_COMP_LOOP_and_5_itm AND and_295_m1c) OR (COMP_LOOP_COMP_LOOP_and_4_itm
      AND and_297_m1c) OR (COMP_LOOP_COMP_LOOP_and_64_itm AND and_299_m1c) OR (COMP_LOOP_COMP_LOOP_and_2_itm
      AND and_302_m1c) OR (COMP_LOOP_COMP_LOOP_and_62_itm AND and_304_m1c) OR (COMP_LOOP_COMP_LOOP_and_305_itm
      AND and_307_m1c) OR (COMP_LOOP_COMP_LOOP_nor_itm AND and_309_m1c) OR (COMP_LOOP_COMP_LOOP_and_14_itm
      AND and_311_m1c);
  COMP_LOOP_or_23_nl <= (COMP_LOOP_COMP_LOOP_and_14_itm AND and_dcpl_257) OR (COMP_LOOP_COMP_LOOP_and_13_itm
      AND and_279_m1c) OR (COMP_LOOP_COMP_LOOP_and_12_itm AND and_281_m1c) OR (COMP_LOOP_COMP_LOOP_and_11_itm
      AND and_284_m1c) OR (COMP_LOOP_COMP_LOOP_and_10_itm AND and_286_m1c) OR (COMP_LOOP_COMP_LOOP_and_9_itm
      AND and_288_m1c) OR (COMP_LOOP_COMP_LOOP_and_8_itm AND and_291_m1c) OR (COMP_LOOP_COMP_LOOP_and_68_itm
      AND and_292_m1c) OR (COMP_LOOP_COMP_LOOP_and_6_itm AND and_295_m1c) OR (COMP_LOOP_COMP_LOOP_and_5_itm
      AND and_297_m1c) OR (COMP_LOOP_COMP_LOOP_and_4_itm AND and_299_m1c) OR (COMP_LOOP_COMP_LOOP_and_64_itm
      AND and_302_m1c) OR (COMP_LOOP_COMP_LOOP_and_2_itm AND and_304_m1c) OR (COMP_LOOP_COMP_LOOP_and_62_itm
      AND and_307_m1c) OR (COMP_LOOP_COMP_LOOP_and_305_itm AND and_309_m1c) OR (COMP_LOOP_COMP_LOOP_nor_itm
      AND and_311_m1c);
  and_276_nl <= (fsm_output(7)) AND mux_tmp_2669;
  mux_2737_nl <= MUX_s_1_2_2(mux_tmp_2736, and_276_nl, fsm_output(1));
  nor_687_nl <= NOT((NOT (fsm_output(9))) OR (fsm_output(6)) OR (fsm_output(10)));
  mux_2734_nl <= MUX_s_1_2_2(nor_687_nl, mux_tmp_2669, fsm_output(7));
  mux_2735_nl <= MUX_s_1_2_2(mux_2734_nl, mux_tmp_2709, and_526_cse);
  mux_2738_nl <= MUX_s_1_2_2(mux_2737_nl, mux_2735_nl, fsm_output(2));
  mux_2739_nl <= MUX_s_1_2_2(mux_tmp_2736, mux_2738_nl, fsm_output(3));
  mux_2730_nl <= MUX_s_1_2_2(mux_tmp_2702, mux_tmp_2675, fsm_output(7));
  mux_2729_nl <= MUX_s_1_2_2(or_tmp_2604, mux_tmp_2675, fsm_output(7));
  mux_2731_nl <= MUX_s_1_2_2(mux_2730_nl, mux_2729_nl, or_3388_cse);
  or_2666_nl <= (NOT(and_526_cse OR (fsm_output(7)))) OR (fsm_output(9));
  mux_2728_nl <= MUX_s_1_2_2((fsm_output(6)), or_tmp_167, or_2666_nl);
  mux_2732_nl <= MUX_s_1_2_2(mux_2731_nl, mux_2728_nl, fsm_output(2));
  and_454_nl <= (fsm_output(2)) AND (fsm_output(0)) AND (fsm_output(1)) AND (fsm_output(7));
  mux_2727_nl <= MUX_s_1_2_2(mux_tmp_2675, mux_tmp_2693, and_454_nl);
  mux_2733_nl <= MUX_s_1_2_2(mux_2732_nl, mux_2727_nl, fsm_output(3));
  mux_2740_nl <= MUX_s_1_2_2(mux_2739_nl, mux_2733_nl, fsm_output(8));
  mux_2725_nl <= MUX_s_1_2_2((NOT mux_2698_itm), mux_tmp_2675, fsm_output(7));
  mux_2721_nl <= MUX_s_1_2_2(mux_tmp_2675, mux_544_cse, fsm_output(7));
  mux_2722_nl <= MUX_s_1_2_2(mux_tmp_2690, mux_2721_nl, or_3388_cse);
  mux_2723_nl <= MUX_s_1_2_2(mux_tmp_2690, mux_2722_nl, fsm_output(2));
  mux_2717_nl <= MUX_s_1_2_2((NOT or_tmp_167), or_352_cse, fsm_output(9));
  mux_2718_nl <= MUX_s_1_2_2(mux_tmp_2693, mux_2717_nl, fsm_output(7));
  mux_2719_nl <= MUX_s_1_2_2(mux_2718_nl, mux_tmp_2715, and_526_cse);
  mux_2716_nl <= MUX_s_1_2_2(mux_tmp_2715, mux_tmp_2672, fsm_output(1));
  mux_2720_nl <= MUX_s_1_2_2(mux_2719_nl, mux_2716_nl, fsm_output(2));
  mux_2724_nl <= MUX_s_1_2_2(mux_2723_nl, mux_2720_nl, fsm_output(3));
  mux_2726_nl <= MUX_s_1_2_2(mux_2725_nl, mux_2724_nl, fsm_output(8));
  mux_2741_nl <= MUX_s_1_2_2(mux_2740_nl, mux_2726_nl, fsm_output(5));
  mux_2710_nl <= MUX_s_1_2_2(mux_tmp_2709, mux_tmp_2706, fsm_output(1));
  mux_2707_nl <= MUX_s_1_2_2(mux_tmp_2706, mux_tmp_2703, and_526_cse);
  mux_2711_nl <= MUX_s_1_2_2(mux_2710_nl, mux_2707_nl, fsm_output(2));
  mux_2704_nl <= MUX_s_1_2_2(mux_tmp_2703, mux_tmp_2700, fsm_output(1));
  mux_2699_nl <= MUX_s_1_2_2((NOT mux_2698_itm), or_tmp_167, fsm_output(7));
  mux_2701_nl <= MUX_s_1_2_2(mux_tmp_2700, mux_2699_nl, or_3388_cse);
  mux_2705_nl <= MUX_s_1_2_2(mux_2704_nl, mux_2701_nl, fsm_output(2));
  mux_2712_nl <= MUX_s_1_2_2(mux_2711_nl, mux_2705_nl, fsm_output(3));
  mux_2694_nl <= MUX_s_1_2_2(mux_tmp_2675, mux_tmp_2693, fsm_output(7));
  mux_2695_nl <= MUX_s_1_2_2(mux_2694_nl, mux_tmp_2691, fsm_output(1));
  mux_2692_nl <= MUX_s_1_2_2(mux_tmp_2691, mux_tmp_2690, or_3388_cse);
  mux_2696_nl <= MUX_s_1_2_2(mux_2695_nl, mux_2692_nl, fsm_output(2));
  mux_2697_nl <= MUX_s_1_2_2(mux_2696_nl, mux_tmp_2690, fsm_output(3));
  mux_2713_nl <= MUX_s_1_2_2(mux_2712_nl, mux_2697_nl, fsm_output(8));
  mux_2684_nl <= MUX_s_1_2_2(nor_tmp_48, (fsm_output(6)), fsm_output(9));
  mux_2685_nl <= MUX_s_1_2_2((NOT mux_2684_nl), mux_tmp_2675, fsm_output(7));
  mux_2686_nl <= MUX_s_1_2_2(mux_2685_nl, mux_tmp_2682, and_526_cse);
  mux_2680_nl <= MUX_s_1_2_2(not_tmp_500, mux_tmp_2675, fsm_output(7));
  mux_2683_nl <= MUX_s_1_2_2(mux_tmp_2682, mux_2680_nl, fsm_output(1));
  mux_2687_nl <= MUX_s_1_2_2(mux_2686_nl, mux_2683_nl, fsm_output(2));
  or_2658_nl <= (fsm_output(0)) OR (fsm_output(1)) OR (fsm_output(7));
  mux_2678_nl <= MUX_s_1_2_2(not_tmp_500, mux_tmp_2675, or_2658_nl);
  mux_2674_nl <= MUX_s_1_2_2((fsm_output(6)), or_tmp_167, and_458_cse);
  mux_2679_nl <= MUX_s_1_2_2(mux_2678_nl, mux_2674_nl, fsm_output(2));
  mux_2688_nl <= MUX_s_1_2_2(mux_2687_nl, mux_2679_nl, fsm_output(3));
  mux_2671_nl <= MUX_s_1_2_2(mux_544_cse, mux_tmp_2669, fsm_output(7));
  mux_2673_nl <= MUX_s_1_2_2(mux_tmp_2672, mux_2671_nl, and_459_cse);
  mux_2689_nl <= MUX_s_1_2_2(mux_2688_nl, mux_2673_nl, fsm_output(8));
  mux_2714_nl <= MUX_s_1_2_2(mux_2713_nl, mux_2689_nl, fsm_output(5));
  and_312_nl <= and_dcpl_236 AND and_dcpl_127;
  COMP_LOOP_or_29_nl <= ((NOT (modulo_result_rem_cmp_z(63))) AND and_317_m1c) OR
      (NOT(mux_2840_itm OR (modulo_result_rem_cmp_z(63))));
  COMP_LOOP_or_30_nl <= ((modulo_result_rem_cmp_z(63)) AND and_317_m1c) OR ((NOT
      mux_2840_itm) AND (modulo_result_rem_cmp_z(63)));
  COMP_LOOP_and_277_nl <= COMP_LOOP_COMP_LOOP_nor_1_itm AND mux_2771_m1c;
  COMP_LOOP_COMP_LOOP_and_932_nl <= (COMP_LOOP_acc_10_cse_12_1_1_sva(0)) AND COMP_LOOP_nor_11_itm
      AND mux_2771_m1c;
  COMP_LOOP_COMP_LOOP_and_934_nl <= (COMP_LOOP_acc_10_cse_12_1_1_sva(1)) AND COMP_LOOP_nor_12_itm
      AND mux_2771_m1c;
  COMP_LOOP_and_1_nl <= COMP_LOOP_COMP_LOOP_and_137_itm AND mux_2771_m1c;
  COMP_LOOP_COMP_LOOP_and_936_nl <= (COMP_LOOP_acc_10_cse_12_1_1_sva(2)) AND COMP_LOOP_nor_134_itm
      AND mux_2771_m1c;
  COMP_LOOP_and_2_nl <= COMP_LOOP_COMP_LOOP_and_139_itm AND mux_2771_m1c;
  COMP_LOOP_and_3_nl <= COMP_LOOP_COMP_LOOP_and_140_itm AND mux_2771_m1c;
  COMP_LOOP_and_4_nl <= COMP_LOOP_COMP_LOOP_and_141_itm AND mux_2771_m1c;
  COMP_LOOP_COMP_LOOP_and_930_nl <= (COMP_LOOP_acc_10_cse_12_1_1_sva(3)) AND COMP_LOOP_nor_137_itm
      AND mux_2771_m1c;
  COMP_LOOP_and_5_nl <= COMP_LOOP_COMP_LOOP_and_143_itm AND mux_2771_m1c;
  COMP_LOOP_and_6_nl <= COMP_LOOP_COMP_LOOP_and_144_itm AND mux_2771_m1c;
  COMP_LOOP_and_7_nl <= COMP_LOOP_COMP_LOOP_and_145_itm AND mux_2771_m1c;
  COMP_LOOP_and_8_nl <= COMP_LOOP_COMP_LOOP_and_146_itm AND mux_2771_m1c;
  COMP_LOOP_and_9_nl <= COMP_LOOP_COMP_LOOP_and_147_itm AND mux_2771_m1c;
  COMP_LOOP_and_10_nl <= COMP_LOOP_COMP_LOOP_and_148_itm AND mux_2771_m1c;
  COMP_LOOP_and_11_nl <= COMP_LOOP_COMP_LOOP_and_149_itm AND mux_2771_m1c;
  nand_2_nl <= NOT((fsm_output(5)) AND mux_125_cse);
  mux_126_nl <= MUX_s_1_2_2(nand_2_nl, or_tmp_68, fsm_output(2));
  or_92_nl <= (NOT (fsm_output(2))) OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR
      (fsm_output(3)) OR (NOT (fsm_output(8))) OR (fsm_output(6)) OR (fsm_output(10));
  mux_127_nl <= MUX_s_1_2_2(mux_126_nl, or_92_nl, fsm_output(9));
  nand_3_nl <= NOT((fsm_output(4)) AND (NOT mux_127_nl));
  or_91_nl <= (fsm_output(2)) OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR mux_tmp_119;
  or_89_nl <= (NOT (fsm_output(2))) OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR
      (fsm_output(3)) OR (fsm_output(8)) OR (NOT (fsm_output(6))) OR (fsm_output(10));
  mux_123_nl <= MUX_s_1_2_2(or_91_nl, or_89_nl, fsm_output(9));
  or_88_nl <= (fsm_output(9)) OR (NOT((fsm_output(2)) AND (fsm_output(5)) AND (fsm_output(7))
      AND (fsm_output(3)) AND (fsm_output(8)) AND (fsm_output(6)) AND (fsm_output(10))));
  mux_124_nl <= MUX_s_1_2_2(mux_123_nl, or_88_nl, fsm_output(4));
  mux_128_nl <= MUX_s_1_2_2(nand_3_nl, mux_124_nl, fsm_output(1));
  or_87_nl <= (fsm_output(2)) OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR (NOT
      (fsm_output(3))) OR (fsm_output(8)) OR not_tmp_49;
  or_85_nl <= (NOT (fsm_output(2))) OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR
      mux_tmp_119;
  mux_120_nl <= MUX_s_1_2_2(or_87_nl, or_85_nl, fsm_output(9));
  or_81_nl <= (fsm_output(9)) OR (fsm_output(2)) OR (fsm_output(5)) OR (NOT (fsm_output(7)))
      OR (fsm_output(3)) OR (NOT (fsm_output(8))) OR (fsm_output(6)) OR (fsm_output(10));
  mux_121_nl <= MUX_s_1_2_2(mux_120_nl, or_81_nl, fsm_output(4));
  or_79_nl <= (NOT (fsm_output(2))) OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR
      (fsm_output(3)) OR (NOT (fsm_output(8))) OR (fsm_output(6)) OR (NOT (fsm_output(10)));
  nand_373_nl <= NOT((fsm_output(5)) AND (fsm_output(7)) AND (fsm_output(3)) AND
      (fsm_output(8)) AND (fsm_output(6)) AND (NOT (fsm_output(10))));
  mux_116_nl <= MUX_s_1_2_2(nand_373_nl, or_tmp_68, fsm_output(2));
  mux_117_nl <= MUX_s_1_2_2(or_79_nl, mux_116_nl, fsm_output(9));
  mux_118_nl <= MUX_s_1_2_2(or_80_cse, mux_117_nl, fsm_output(4));
  mux_122_nl <= MUX_s_1_2_2(mux_121_nl, mux_118_nl, fsm_output(1));
  mux_129_nl <= MUX_s_1_2_2(mux_128_nl, mux_122_nl, fsm_output(0));
  mux_2975_nl <= MUX_s_1_2_2(mux_2203_cse, mux_tmp_2159, fsm_output(6));
  mux_2976_nl <= MUX_s_1_2_2(mux_2975_nl, mux_tmp_2920, fsm_output(0));
  mux_2973_nl <= MUX_s_1_2_2(or_tmp_2280, or_tmp_2729, fsm_output(6));
  mux_2972_nl <= MUX_s_1_2_2(or_tmp_2731, or_tmp_2729, fsm_output(6));
  mux_2974_nl <= MUX_s_1_2_2(mux_2973_nl, mux_2972_nl, fsm_output(0));
  mux_2977_nl <= MUX_s_1_2_2(mux_2976_nl, mux_2974_nl, fsm_output(8));
  mux_2971_nl <= MUX_s_1_2_2(mux_tmp_2879, or_tmp_2734, fsm_output(8));
  mux_2978_nl <= MUX_s_1_2_2(mux_2977_nl, mux_2971_nl, fsm_output(3));
  mux_2967_nl <= MUX_s_1_2_2(or_tmp_2749, mux_tmp_2912, fsm_output(6));
  mux_2968_nl <= MUX_s_1_2_2(mux_2967_nl, nand_tmp_71, fsm_output(0));
  mux_2969_nl <= MUX_s_1_2_2(mux_2968_nl, or_3532_cse, fsm_output(8));
  mux_2963_nl <= MUX_s_1_2_2((NOT (fsm_output(10))), or_tmp_2276, fsm_output(9));
  mux_2964_nl <= MUX_s_1_2_2(mux_2963_nl, or_tmp_2731, fsm_output(6));
  mux_2965_nl <= MUX_s_1_2_2(mux_2964_nl, mux_tmp_2906, fsm_output(0));
  mux_2966_nl <= MUX_s_1_2_2(or_tmp_2740, mux_2965_nl, fsm_output(8));
  mux_2970_nl <= MUX_s_1_2_2(mux_2969_nl, mux_2966_nl, fsm_output(3));
  mux_2979_nl <= MUX_s_1_2_2(mux_2978_nl, mux_2970_nl, fsm_output(5));
  or_2810_nl <= (fsm_output(6)) OR mux_tmp_2848;
  mux_2960_nl <= MUX_s_1_2_2(nand_tmp_69, or_2810_nl, fsm_output(8));
  nand_72_nl <= NOT((fsm_output(6)) AND (NOT mux_tmp_2895));
  mux_2959_nl <= MUX_s_1_2_2(nand_72_nl, or_tmp_2743, fsm_output(8));
  mux_2961_nl <= MUX_s_1_2_2(mux_2960_nl, mux_2959_nl, fsm_output(3));
  mux_2956_nl <= MUX_s_1_2_2(mux_tmp_2867, mux_tmp_2890, fsm_output(0));
  mux_2955_nl <= MUX_s_1_2_2(mux_tmp_2862, mux_tmp_2888, fsm_output(0));
  mux_2957_nl <= MUX_s_1_2_2(mux_2956_nl, mux_2955_nl, fsm_output(8));
  mux_2953_nl <= MUX_s_1_2_2(mux_tmp_2850, mux_tmp_2886, fsm_output(0));
  mux_2954_nl <= MUX_s_1_2_2(mux_tmp_2878, mux_2953_nl, fsm_output(8));
  mux_2958_nl <= MUX_s_1_2_2(mux_2957_nl, mux_2954_nl, fsm_output(3));
  mux_2962_nl <= MUX_s_1_2_2(mux_2961_nl, mux_2958_nl, fsm_output(5));
  mux_2980_nl <= MUX_s_1_2_2(mux_2979_nl, mux_2962_nl, fsm_output(4));
  or_2809_nl <= (fsm_output(6)) OR mux_tmp_2851;
  mux_2948_nl <= MUX_s_1_2_2(or_2809_nl, or_tmp_2734, fsm_output(0));
  mux_2949_nl <= MUX_s_1_2_2(mux_tmp_2880, mux_2948_nl, fsm_output(8));
  mux_2946_nl <= MUX_s_1_2_2(mux_tmp_2916, mux_tmp_2876, fsm_output(0));
  mux_2947_nl <= MUX_s_1_2_2(mux_2946_nl, or_tmp_2734, fsm_output(8));
  mux_2950_nl <= MUX_s_1_2_2(mux_2949_nl, mux_2947_nl, fsm_output(3));
  mux_2944_nl <= MUX_s_1_2_2(nand_tmp_70, mux_tmp_2910, fsm_output(8));
  mux_2942_nl <= MUX_s_1_2_2(or_tmp_258, mux_tmp_2159, fsm_output(6));
  mux_2943_nl <= MUX_s_1_2_2(or_tmp_2740, mux_2942_nl, fsm_output(8));
  mux_2945_nl <= MUX_s_1_2_2(mux_2944_nl, mux_2943_nl, fsm_output(3));
  mux_2951_nl <= MUX_s_1_2_2(mux_2950_nl, mux_2945_nl, fsm_output(5));
  mux_2938_nl <= MUX_s_1_2_2(nand_tmp_69, nand_tmp_67, fsm_output(0));
  mux_2936_nl <= MUX_s_1_2_2(or_tmp_2731, or_tmp_2749, fsm_output(6));
  mux_2937_nl <= MUX_s_1_2_2(or_tmp_2745, mux_2936_nl, fsm_output(0));
  mux_2939_nl <= MUX_s_1_2_2(mux_2938_nl, mux_2937_nl, fsm_output(8));
  mux_2933_nl <= MUX_s_1_2_2(or_tmp_2746, mux_tmp_2856, fsm_output(6));
  mux_2934_nl <= MUX_s_1_2_2(nand_tmp_68, mux_2933_nl, fsm_output(0));
  mux_2935_nl <= MUX_s_1_2_2(mux_2934_nl, or_3532_cse, fsm_output(8));
  mux_2940_nl <= MUX_s_1_2_2(mux_2939_nl, mux_2935_nl, fsm_output(3));
  mux_2930_nl <= MUX_s_1_2_2(mux_tmp_2159, or_tmp_2736, fsm_output(6));
  mux_2931_nl <= MUX_s_1_2_2(mux_2930_nl, mux_tmp_2888, fsm_output(8));
  mux_2927_nl <= MUX_s_1_2_2((NOT (fsm_output(7))), mux_2926_cse, fsm_output(9));
  or_2807_nl <= (fsm_output(6)) OR mux_2927_nl;
  mux_2928_nl <= MUX_s_1_2_2(or_2807_nl, or_tmp_2734, fsm_output(0));
  mux_2929_nl <= MUX_s_1_2_2(mux_2928_nl, mux_tmp_2844, fsm_output(8));
  mux_2932_nl <= MUX_s_1_2_2(mux_2931_nl, mux_2929_nl, fsm_output(3));
  mux_2941_nl <= MUX_s_1_2_2(mux_2940_nl, mux_2932_nl, fsm_output(5));
  mux_2952_nl <= MUX_s_1_2_2(mux_2951_nl, mux_2941_nl, fsm_output(4));
  mux_2981_nl <= MUX_s_1_2_2(mux_2980_nl, mux_2952_nl, fsm_output(2));
  mux_2921_nl <= MUX_s_1_2_2(mux_tmp_2920, or_tmp_2734, fsm_output(8));
  mux_2917_nl <= MUX_s_1_2_2(mux_tmp_2856, mux_tmp_2851, fsm_output(6));
  mux_2918_nl <= MUX_s_1_2_2(mux_2917_nl, mux_tmp_2916, fsm_output(0));
  mux_2919_nl <= MUX_s_1_2_2(mux_2918_nl, or_tmp_2734, fsm_output(8));
  mux_2922_nl <= MUX_s_1_2_2(mux_2921_nl, mux_2919_nl, fsm_output(3));
  mux_2913_nl <= MUX_s_1_2_2(nand_tmp_71, nand_tmp_70, fsm_output(0));
  mux_2911_nl <= MUX_s_1_2_2(or_3532_cse, mux_tmp_2910, fsm_output(0));
  mux_2914_nl <= MUX_s_1_2_2(mux_2913_nl, mux_2911_nl, fsm_output(8));
  mux_2905_nl <= MUX_s_1_2_2(or_tmp_258, mux_tmp_2851, fsm_output(6));
  mux_2907_nl <= MUX_s_1_2_2(mux_tmp_2906, mux_2905_nl, fsm_output(0));
  mux_2908_nl <= MUX_s_1_2_2(or_tmp_2740, mux_2907_nl, fsm_output(8));
  mux_2915_nl <= MUX_s_1_2_2(mux_2914_nl, mux_2908_nl, fsm_output(3));
  mux_2923_nl <= MUX_s_1_2_2(mux_2922_nl, mux_2915_nl, fsm_output(5));
  mux_2899_nl <= MUX_s_1_2_2(or_tmp_2742, or_tmp_2746, fsm_output(6));
  mux_2900_nl <= MUX_s_1_2_2(mux_2899_nl, or_tmp_2745, fsm_output(0));
  mux_2902_nl <= MUX_s_1_2_2(nand_tmp_69, mux_2900_nl, fsm_output(8));
  mux_2896_nl <= MUX_s_1_2_2(or_tmp_2739, mux_tmp_2895, fsm_output(6));
  mux_2897_nl <= MUX_s_1_2_2(mux_2896_nl, nand_tmp_68, fsm_output(0));
  mux_2894_nl <= MUX_s_1_2_2(or_tmp_2743, or_3532_cse, fsm_output(0));
  mux_2898_nl <= MUX_s_1_2_2(mux_2897_nl, mux_2894_nl, fsm_output(8));
  mux_2903_nl <= MUX_s_1_2_2(mux_2902_nl, mux_2898_nl, fsm_output(3));
  mux_2889_nl <= MUX_s_1_2_2(or_tmp_2731, or_tmp_2281, fsm_output(6));
  mux_2891_nl <= MUX_s_1_2_2(mux_tmp_2890, mux_2889_nl, fsm_output(0));
  mux_2892_nl <= MUX_s_1_2_2(mux_2891_nl, mux_tmp_2888, fsm_output(8));
  mux_2887_nl <= MUX_s_1_2_2(or_tmp_2734, mux_tmp_2886, fsm_output(8));
  mux_2893_nl <= MUX_s_1_2_2(mux_2892_nl, mux_2887_nl, fsm_output(3));
  mux_2904_nl <= MUX_s_1_2_2(mux_2903_nl, mux_2893_nl, fsm_output(5));
  mux_2924_nl <= MUX_s_1_2_2(mux_2923_nl, mux_2904_nl, fsm_output(4));
  mux_2881_nl <= MUX_s_1_2_2(mux_tmp_2880, mux_tmp_2879, fsm_output(0));
  mux_2882_nl <= MUX_s_1_2_2(mux_2881_nl, mux_tmp_2878, fsm_output(8));
  mux_2873_nl <= MUX_s_1_2_2(mux_tmp_2848, or_tmp_2739, fsm_output(6));
  mux_2874_nl <= MUX_s_1_2_2(or_tmp_2734, mux_2873_nl, fsm_output(0));
  mux_2877_nl <= MUX_s_1_2_2(mux_tmp_2876, mux_2874_nl, fsm_output(8));
  mux_2883_nl <= MUX_s_1_2_2(mux_2882_nl, mux_2877_nl, fsm_output(3));
  mux_2869_nl <= MUX_s_1_2_2((NOT or_tmp_2280), or_tmp_2276, fsm_output(9));
  mux_2870_nl <= MUX_s_1_2_2(mux_2869_nl, or_tmp_2280, fsm_output(6));
  mux_2871_nl <= MUX_s_1_2_2(or_tmp_2740, mux_2870_nl, fsm_output(8));
  mux_2864_nl <= MUX_s_1_2_2(or_tmp_2276, mux_tmp_2863, fsm_output(6));
  mux_2865_nl <= MUX_s_1_2_2(mux_2864_nl, mux_tmp_2862, fsm_output(0));
  mux_2868_nl <= MUX_s_1_2_2(mux_tmp_2867, mux_2865_nl, fsm_output(8));
  mux_2872_nl <= MUX_s_1_2_2(mux_2871_nl, mux_2868_nl, fsm_output(3));
  mux_2884_nl <= MUX_s_1_2_2(mux_2883_nl, mux_2872_nl, fsm_output(5));
  or_2797_nl <= (fsm_output(6)) OR or_tmp_2731;
  mux_2859_nl <= MUX_s_1_2_2(nand_tmp_67, or_2797_nl, fsm_output(8));
  nand_66_nl <= NOT((fsm_output(6)) AND (NOT mux_tmp_2856));
  mux_2857_nl <= MUX_s_1_2_2(nand_66_nl, or_3532_cse, fsm_output(8));
  mux_2860_nl <= MUX_s_1_2_2(mux_2859_nl, mux_2857_nl, fsm_output(3));
  mux_2852_nl <= MUX_s_1_2_2(mux_tmp_2851, or_tmp_2736, fsm_output(6));
  mux_2853_nl <= MUX_s_1_2_2(mux_2852_nl, or_tmp_2734, fsm_output(0));
  mux_2854_nl <= MUX_s_1_2_2(mux_2853_nl, mux_tmp_2850, fsm_output(8));
  mux_2842_nl <= MUX_s_1_2_2(or_tmp_2729, mux_tmp_2841, fsm_output(6));
  mux_2845_nl <= MUX_s_1_2_2(mux_tmp_2844, mux_2842_nl, fsm_output(0));
  mux_2847_nl <= MUX_s_1_2_2(or_tmp_2734, mux_2845_nl, fsm_output(8));
  mux_2855_nl <= MUX_s_1_2_2(mux_2854_nl, mux_2847_nl, fsm_output(3));
  mux_2861_nl <= MUX_s_1_2_2(mux_2860_nl, mux_2855_nl, fsm_output(5));
  mux_2885_nl <= MUX_s_1_2_2(mux_2884_nl, mux_2861_nl, fsm_output(4));
  mux_2925_nl <= MUX_s_1_2_2(mux_2924_nl, mux_2885_nl, fsm_output(2));
  COMP_LOOP_COMP_LOOP_and_17_nl <= CONV_SL_1_1(z_out_2_12_1(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0011"));
  COMP_LOOP_1_acc_8_nl <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_10_lpi_4_dfm) -
      SIGNED(COMP_LOOP_10_mul_mut), 64));
  nor_631_nl <= NOT((NOT (fsm_output(3))) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(1)))
      OR (fsm_output(9)) OR (fsm_output(2)) OR (fsm_output(6)) OR (fsm_output(10)));
  mux_3284_nl <= MUX_s_1_2_2(or_2921_cse, mux_3935_cse, fsm_output(0));
  nor_632_nl <= NOT((fsm_output(3)) OR mux_3284_nl);
  mux_3285_nl <= MUX_s_1_2_2(nor_631_nl, nor_632_nl, fsm_output(8));
  and_417_nl <= (fsm_output(8)) AND (fsm_output(3)) AND (NOT mux_3245_cse);
  mux_3286_nl <= MUX_s_1_2_2(mux_3285_nl, and_417_nl, fsm_output(5));
  or_2958_nl <= (fsm_output(9)) OR (NOT (fsm_output(2))) OR (fsm_output(6)) OR (fsm_output(10));
  or_2957_nl <= (NOT (fsm_output(9))) OR (NOT (fsm_output(2))) OR (fsm_output(6))
      OR (fsm_output(10));
  mux_3279_nl <= MUX_s_1_2_2(or_2958_nl, or_2957_nl, fsm_output(1));
  or_2959_nl <= (fsm_output(0)) OR mux_3279_nl;
  or_2954_nl <= (fsm_output(1)) OR (fsm_output(9)) OR (fsm_output(2)) OR (fsm_output(6))
      OR (NOT (fsm_output(10)));
  mux_3278_nl <= MUX_s_1_2_2(or_2912_cse, or_2954_nl, fsm_output(0));
  mux_3280_nl <= MUX_s_1_2_2(or_2959_nl, mux_3278_nl, fsm_output(3));
  nor_633_nl <= NOT((NOT (fsm_output(5))) OR (fsm_output(8)) OR mux_3280_nl);
  mux_3287_nl <= MUX_s_1_2_2(mux_3286_nl, nor_633_nl, fsm_output(4));
  and_418_nl <= (fsm_output(8)) AND (fsm_output(3)) AND (fsm_output(0)) AND (fsm_output(1))
      AND (NOT (fsm_output(9))) AND (fsm_output(2)) AND (fsm_output(6)) AND (NOT
      (fsm_output(10)));
  nor_634_nl <= NOT((fsm_output(8)) OR (fsm_output(3)) OR (fsm_output(0)) OR (fsm_output(1))
      OR (fsm_output(9)) OR (fsm_output(2)) OR (fsm_output(6)) OR (NOT (fsm_output(10))));
  mux_3276_nl <= MUX_s_1_2_2(and_418_nl, nor_634_nl, fsm_output(5));
  nand_92_nl <= NOT((fsm_output(3)) AND (NOT mux_3254_cse));
  or_2943_nl <= (fsm_output(1)) OR (fsm_output(9)) OR nand_367_cse;
  mux_3273_nl <= MUX_s_1_2_2(or_2905_cse, or_2943_nl, fsm_output(0));
  or_2945_nl <= (fsm_output(3)) OR mux_3273_nl;
  mux_3275_nl <= MUX_s_1_2_2(nand_92_nl, or_2945_nl, fsm_output(8));
  nor_635_nl <= NOT((fsm_output(5)) OR mux_3275_nl);
  mux_3277_nl <= MUX_s_1_2_2(mux_3276_nl, nor_635_nl, fsm_output(4));
  mux_3288_nl <= MUX_s_1_2_2(mux_3287_nl, mux_3277_nl, fsm_output(7));
  COMP_LOOP_COMP_LOOP_and_10_nl <= CONV_SL_1_1(VEC_LOOP_j_sva_11_0(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1011"));
  COMP_LOOP_1_acc_nl <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED((z_out_1(5 DOWNTO 0))
      & STD_LOGIC_VECTOR'( "0000")) + SIGNED('1' & (NOT (STAGE_LOOP_lshift_psp_sva(9
      DOWNTO 1)))) + SIGNED'( "0000000001"), 10));
  or_2647_nl <= CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00"));
  mux_2642_nl <= MUX_s_1_2_2(nor_609_cse, and_757_cse, or_2647_nl);
  mux_3330_nl <= MUX_s_1_2_2(mux_tmp_3329, mux_2642_nl, or_3388_cse);
  mux_3331_nl <= MUX_s_1_2_2(mux_3330_nl, mux_2643_cse, fsm_output(3));
  or_3032_nl <= (fsm_output(1)) OR (fsm_output(6));
  mux_3326_nl <= MUX_s_1_2_2(mux_tmp_2640, and_756_cse, or_3032_nl);
  and_410_nl <= ((NOT((NOT (fsm_output(0))) OR (NOT (fsm_output(1))) OR (fsm_output(6))))
      OR (fsm_output(7))) AND CONV_SL_1_1(fsm_output(10 DOWNTO 9)=STD_LOGIC_VECTOR'("11"));
  mux_3327_nl <= MUX_s_1_2_2(mux_3326_nl, and_410_nl, fsm_output(3));
  mux_3332_nl <= MUX_s_1_2_2(mux_3331_nl, mux_3327_nl, fsm_output(4));
  and_411_nl <= ((NOT((NOT (fsm_output(3))) OR (fsm_output(6)))) OR (fsm_output(7)))
      AND CONV_SL_1_1(fsm_output(10 DOWNTO 9)=STD_LOGIC_VECTOR'("11"));
  mux_3325_nl <= MUX_s_1_2_2(mux_2643_cse, and_411_nl, fsm_output(4));
  mux_3333_nl <= MUX_s_1_2_2(mux_3332_nl, mux_3325_nl, fsm_output(2));
  mux_3334_nl <= MUX_s_1_2_2(mux_tmp_3329, mux_3333_nl, fsm_output(5));
  or_3037_nl <= (fsm_output(3)) OR (fsm_output(1)) OR (fsm_output(2)) OR (fsm_output(9));
  mux_3337_nl <= MUX_s_1_2_2((fsm_output(9)), or_3037_nl, and_407_cse);
  and_408_nl <= (fsm_output(0)) AND (fsm_output(1)) AND (fsm_output(2)) AND (fsm_output(9));
  or_3036_nl <= CONV_SL_1_1(fsm_output(5 DOWNTO 3)/=STD_LOGIC_VECTOR'("000"));
  mux_3336_nl <= MUX_s_1_2_2(and_408_nl, (fsm_output(9)), or_3036_nl);
  mux_3338_nl <= MUX_s_1_2_2((NOT mux_3337_nl), mux_3336_nl, fsm_output(7));
  mux_3339_nl <= MUX_s_1_2_2(mux_3338_nl, and_458_cse, fsm_output(6));
  mux_3340_nl <= MUX_s_1_2_2(mux_3339_nl, (fsm_output(9)), fsm_output(8));
  mux_3346_nl <= MUX_s_1_2_2(mux_tmp_3341, nor_tmp_457, fsm_output(3));
  mux_3347_nl <= MUX_s_1_2_2(not_tmp_90, mux_3346_nl, fsm_output(4));
  mux_3344_nl <= MUX_s_1_2_2(not_tmp_90, nor_tmp_457, fsm_output(4));
  mux_3345_nl <= MUX_s_1_2_2(mux_3344_nl, mux_tmp_3343, fsm_output(0));
  mux_3348_nl <= MUX_s_1_2_2(mux_3347_nl, mux_3345_nl, fsm_output(1));
  mux_3349_nl <= MUX_s_1_2_2(mux_3348_nl, mux_tmp_3343, fsm_output(2));
  mux_3350_nl <= MUX_s_1_2_2(not_tmp_90, mux_3349_nl, fsm_output(5));
  nor_623_nl <= NOT((fsm_output(5)) OR (fsm_output(8)));
  mux_3351_nl <= MUX_s_1_2_2(nor_623_nl, (fsm_output(8)), fsm_output(6));
  mux_3353_nl <= MUX_s_1_2_2(mux_648_cse, mux_3351_nl, or_3039_cse);
  mux_3354_nl <= MUX_s_1_2_2(mux_648_cse, mux_3353_nl, fsm_output(4));
  mux_3355_nl <= MUX_s_1_2_2(mux_3354_nl, (fsm_output(8)), fsm_output(7));
  and_401_nl <= (fsm_output(0)) AND (fsm_output(7)) AND (fsm_output(8));
  mux_3356_nl <= MUX_s_1_2_2(not_tmp_133, and_401_nl, fsm_output(3));
  and_402_nl <= (fsm_output(3)) AND (fsm_output(7)) AND (fsm_output(8));
  mux_3357_nl <= MUX_s_1_2_2(mux_3356_nl, and_402_nl, or_2368_cse);
  mux_3358_nl <= MUX_s_1_2_2(not_tmp_133, mux_3357_nl, and_407_cse);
  mux_3359_nl <= MUX_s_1_2_2(mux_3358_nl, and_404_cse, fsm_output(6));
  or_3045_nl <= CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")) OR
      mux_tmp_3361;
  mux_3362_nl <= MUX_s_1_2_2(or_3079_cse, or_3045_nl, fsm_output(4));
  mux_3360_nl <= MUX_s_1_2_2(or_3079_cse, or_3074_cse, fsm_output(4));
  mux_3363_nl <= MUX_s_1_2_2(mux_3362_nl, mux_3360_nl, fsm_output(1));
  mux_3364_nl <= MUX_s_1_2_2(mux_3363_nl, (NOT or_3074_cse), fsm_output(9));
  or_3048_nl <= (or_3039_cse AND (fsm_output(4))) OR (fsm_output(9));
  mux_3365_nl <= MUX_s_1_2_2((fsm_output(9)), or_3048_nl, fsm_output(5));
  nor_621_nl <= NOT((fsm_output(7)) OR mux_3365_nl);
  and_334_nl <= (fsm_output(7)) AND (fsm_output(5)) AND (and_459_cse OR (fsm_output(4)))
      AND (fsm_output(9));
  mux_3366_nl <= MUX_s_1_2_2(nor_621_nl, and_334_nl, fsm_output(6));
  mux_3367_nl <= MUX_s_1_2_2(mux_3366_nl, (fsm_output(9)), fsm_output(8));
  nor_619_nl <= NOT(CONV_SL_1_1(fsm_output(9 DOWNTO 8)/=STD_LOGIC_VECTOR'("00")));
  nor_620_nl <= NOT((fsm_output(3)) OR (fsm_output(2)) OR (fsm_output(1)) OR (fsm_output(8))
      OR (fsm_output(9)));
  mux_3370_nl <= MUX_s_1_2_2(nor_619_nl, nor_620_nl, and_407_cse);
  and_30_nl <= (fsm_output(8)) AND (fsm_output(2)) AND or_3388_cse AND (fsm_output(9));
  mux_3368_nl <= MUX_s_1_2_2(and_30_nl, nor_tmp_82, fsm_output(3));
  and_337_nl <= (fsm_output(4)) AND mux_3368_nl;
  mux_3369_nl <= MUX_s_1_2_2(and_337_nl, nor_tmp_82, fsm_output(5));
  mux_3371_nl <= MUX_s_1_2_2(mux_3370_nl, mux_3369_nl, fsm_output(6));
  mux_3372_nl <= MUX_s_1_2_2(mux_3371_nl, nor_tmp_82, fsm_output(7));
  nor_1596_nl <= NOT(CONV_SL_1_1(fsm_output(9 DOWNTO 7)/=STD_LOGIC_VECTOR'("000")));
  nor_1597_nl <= NOT((fsm_output(3)) OR (fsm_output(1)) OR (fsm_output(7)) OR (fsm_output(8))
      OR (fsm_output(9)));
  and_749_nl <= (fsm_output(3)) AND (fsm_output(7)) AND (fsm_output(8)) AND (fsm_output(9));
  mux_3373_nl <= MUX_s_1_2_2(nor_1597_nl, and_749_nl, fsm_output(2));
  mux_3374_nl <= MUX_s_1_2_2(nor_1596_nl, mux_3373_nl, and_407_cse);
  and_750_nl <= CONV_SL_1_1(fsm_output(9 DOWNTO 7)=STD_LOGIC_VECTOR'("111"));
  mux_3375_nl <= MUX_s_1_2_2(mux_3374_nl, and_750_nl, fsm_output(6));
  or_3060_nl <= (NOT(CONV_SL_1_1(fsm_output(9 DOWNTO 6)/=STD_LOGIC_VECTOR'("0000"))))
      OR (fsm_output(10));
  mux_3379_nl <= MUX_s_1_2_2(mux_tmp_3378, or_3060_nl, fsm_output(4));
  or_3058_nl <= (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(7)) OR (fsm_output(8))
      OR (fsm_output(9));
  mux_3376_nl <= MUX_s_1_2_2((NOT (fsm_output(10))), (fsm_output(10)), or_3058_nl);
  mux_3377_nl <= MUX_s_1_2_2(mux_3376_nl, or_tmp_2988, fsm_output(0));
  mux_3380_nl <= MUX_s_1_2_2(mux_3379_nl, mux_3377_nl, fsm_output(1));
  mux_3381_nl <= MUX_s_1_2_2(mux_3380_nl, or_tmp_2988, or_2644_cse);
  or_3065_nl <= (fsm_output(1)) OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(10));
  mux_3384_nl <= MUX_s_1_2_2((fsm_output(10)), or_3065_nl, and_407_cse);
  and_394_nl <= or_2368_cse AND (fsm_output(3)) AND (fsm_output(10));
  mux_3383_nl <= MUX_s_1_2_2(and_394_nl, (fsm_output(10)), or_3063_cse);
  mux_3385_nl <= MUX_s_1_2_2((NOT mux_3384_nl), mux_3383_nl, fsm_output(7));
  mux_3386_nl <= MUX_s_1_2_2(mux_3385_nl, and_395_cse, fsm_output(6));
  nor_615_nl <= NOT((fsm_output(7)) OR (fsm_output(10)));
  mux_3388_nl <= MUX_s_1_2_2(nor_615_nl, and_395_cse, fsm_output(6));
  mux_3389_nl <= MUX_s_1_2_2(not_tmp_647, mux_3388_nl, fsm_output(0));
  and_391_nl <= (fsm_output(6)) AND (fsm_output(7)) AND (fsm_output(10));
  mux_3390_nl <= MUX_s_1_2_2(mux_3389_nl, and_391_nl, or_3039_cse);
  mux_3391_nl <= MUX_s_1_2_2(not_tmp_647, mux_3390_nl, and_407_cse);
  nor_613_nl <= NOT((fsm_output(8)) OR (fsm_output(10)));
  nor_614_nl <= NOT((fsm_output(1)) OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(8))
      OR (fsm_output(10)));
  mux_3394_nl <= MUX_s_1_2_2(nor_613_nl, nor_614_nl, and_407_cse);
  and_388_nl <= (fsm_output(4)) AND (fsm_output(3)) AND (fsm_output(8)) AND (fsm_output(10));
  mux_3393_nl <= MUX_s_1_2_2(and_388_nl, nor_tmp_405, fsm_output(5));
  mux_3395_nl <= MUX_s_1_2_2(mux_3394_nl, mux_3393_nl, fsm_output(6));
  mux_3396_nl <= MUX_s_1_2_2(mux_3395_nl, nor_tmp_405, fsm_output(7));
  nor_611_nl <= NOT((fsm_output(7)) OR (fsm_output(8)) OR (fsm_output(10)));
  nor_612_nl <= NOT((fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(7)) OR (fsm_output(8))
      OR (fsm_output(10)));
  and_384_nl <= (fsm_output(2)) AND (fsm_output(3)) AND (fsm_output(0)) AND (fsm_output(7))
      AND (fsm_output(8)) AND (fsm_output(10));
  mux_3398_nl <= MUX_s_1_2_2(nor_612_nl, and_384_nl, fsm_output(1));
  mux_3399_nl <= MUX_s_1_2_2(nor_611_nl, mux_3398_nl, and_407_cse);
  and_386_nl <= (fsm_output(7)) AND (fsm_output(8)) AND (fsm_output(10));
  mux_3400_nl <= MUX_s_1_2_2(mux_3399_nl, and_386_nl, fsm_output(6));
  or_3078_nl <= (or_3039_cse AND (fsm_output(5))) OR CONV_SL_1_1(fsm_output(8 DOWNTO
      6)/=STD_LOGIC_VECTOR'("000"));
  mux_3403_nl <= MUX_s_1_2_2(or_3079_cse, or_3078_nl, fsm_output(4));
  nor_1680_nl <= NOT((fsm_output(10)) OR mux_3403_nl);
  or_3076_nl <= ((and_529_cse OR (fsm_output(3))) AND (fsm_output(5))) OR CONV_SL_1_1(fsm_output(8
      DOWNTO 6)/=STD_LOGIC_VECTOR'("000"));
  mux_3402_nl <= MUX_s_1_2_2(or_3076_nl, or_3074_cse, fsm_output(4));
  and_1162_nl <= (fsm_output(10)) AND mux_3402_nl;
  nor_610_nl <= NOT((fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(1)) OR (fsm_output(9))
      OR (fsm_output(10)));
  mux_3406_nl <= MUX_s_1_2_2(nor_609_cse, nor_610_nl, and_407_cse);
  and_341_nl <= CONV_SL_1_1(fsm_output(3 DOWNTO 2)=STD_LOGIC_VECTOR'("11")) AND or_3388_cse
      AND CONV_SL_1_1(fsm_output(10 DOWNTO 9)=STD_LOGIC_VECTOR'("11"));
  mux_3405_nl <= MUX_s_1_2_2(and_341_nl, and_757_cse, or_3063_cse);
  mux_3407_nl <= MUX_s_1_2_2(mux_3406_nl, mux_3405_nl, fsm_output(7));
  mux_3408_nl <= MUX_s_1_2_2(mux_3407_nl, and_756_cse, fsm_output(6));
  operator_64_false_1_mux_2_nl <= MUX_v_12_2_2((STD_LOGIC_VECTOR'( "0000001") & (NOT
      COMP_LOOP_k_9_4_sva_4_0)), VEC_LOOP_j_sva_11_0, and_dcpl_332);
  operator_64_false_1_mux_3_nl <= MUX_v_10_2_2(STD_LOGIC_VECTOR'( "0000000001"),
      STAGE_LOOP_lshift_psp_sva, and_dcpl_332);
  z_out <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(operator_64_false_1_mux_2_nl),
      13) + CONV_UNSIGNED(UNSIGNED(operator_64_false_1_mux_3_nl), 13), 13));
  COMP_LOOP_COMP_LOOP_or_72_nl <= (NOT(and_dcpl_342 OR and_dcpl_356)) OR and_dcpl_350
      OR and_dcpl_359;
  COMP_LOOP_COMP_LOOP_or_73_nl <= (NOT((operator_66_true_div_cmp_z(63)) OR and_dcpl_342
      OR and_dcpl_356)) OR and_dcpl_350;
  COMP_LOOP_mux1h_575_nl <= MUX1HOT_v_63_4_2((STD_LOGIC_VECTOR'( "000000000000000000000000000000000000000000000000000000")
      & (VEC_LOOP_j_sva_11_0(11 DOWNTO 3))), (NOT (operator_64_false_acc_mut_63_0(62
      DOWNTO 0))), (STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000")
      & COMP_LOOP_k_9_4_sva_4_0), (NOT (operator_66_true_div_cmp_z(62 DOWNTO 0))),
      STD_LOGIC_VECTOR'( and_dcpl_342 & and_dcpl_350 & and_dcpl_356 & and_dcpl_359));
  COMP_LOOP_nor_695_nl <= NOT(and_dcpl_350 OR and_dcpl_356 OR and_dcpl_359);
  COMP_LOOP_COMP_LOOP_and_938_nl <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), COMP_LOOP_k_9_4_sva_4_0,
      COMP_LOOP_nor_695_nl);
  z_out_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_COMP_LOOP_or_72_nl
      & COMP_LOOP_COMP_LOOP_or_73_nl & COMP_LOOP_mux1h_575_nl) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_COMP_LOOP_and_938_nl
      & '1'), 6), 65), 65));
  COMP_LOOP_mux1h_576_nl <= MUX1HOT_v_7_4_2(((z_out_7(5 DOWNTO 0)) & (STAGE_LOOP_lshift_psp_sva(3))),
      (z_out_5(9 DOWNTO 3)), (z_out_4(9 DOWNTO 3)), z_out_7, STD_LOGIC_VECTOR'( and_824_ssc
      & COMP_LOOP_or_54_ssc & COMP_LOOP_or_55_ssc & and_872_ssc));
  COMP_LOOP_or_69_nl <= and_824_ssc OR and_872_ssc;
  COMP_LOOP_mux1h_577_nl <= MUX1HOT_v_3_3_2((STAGE_LOOP_lshift_psp_sva(2 DOWNTO 0)),
      (z_out_5(2 DOWNTO 0)), (z_out_4(2 DOWNTO 0)), STD_LOGIC_VECTOR'( COMP_LOOP_or_69_nl
      & COMP_LOOP_or_54_ssc & COMP_LOOP_or_55_ssc));
  COMP_LOOP_acc_105_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_sva_11_0),
      12), 13) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_mux1h_576_nl & COMP_LOOP_mux1h_577_nl),
      10), 13), 13));
  z_out_2_12_1 <= COMP_LOOP_acc_105_nl(12 DOWNTO 1);
  COMP_LOOP_COMP_LOOP_or_74_nl <= (VEC_LOOP_j_sva_11_0(11)) OR and_dcpl_460 OR and_dcpl_468
      OR and_dcpl_475 OR and_dcpl_481 OR and_dcpl_486 OR and_dcpl_495 OR and_dcpl_500
      OR and_dcpl_503 OR and_dcpl_507 OR and_dcpl_510 OR and_dcpl_513;
  COMP_LOOP_COMP_LOOP_mux_18_nl <= MUX_v_9_2_2((VEC_LOOP_j_sva_11_0(10 DOWNTO 2)),
      (NOT (STAGE_LOOP_lshift_psp_sva(9 DOWNTO 1))), COMP_LOOP_or_61_itm);
  COMP_LOOP_or_70_nl <= (NOT and_dcpl_453) OR and_dcpl_460 OR and_dcpl_468 OR and_dcpl_475
      OR and_dcpl_481 OR and_dcpl_486 OR and_dcpl_495 OR and_dcpl_500 OR and_dcpl_503
      OR and_dcpl_507 OR and_dcpl_510 OR and_dcpl_513;
  COMP_LOOP_COMP_LOOP_mux_19_nl <= MUX_v_5_2_2((STD_LOGIC_VECTOR'( "00") & (COMP_LOOP_k_9_4_sva_4_0(4
      DOWNTO 2))), COMP_LOOP_k_9_4_sva_4_0, COMP_LOOP_or_61_itm);
  COMP_LOOP_COMP_LOOP_or_75_nl <= ((COMP_LOOP_k_9_4_sva_4_0(1)) AND (NOT(and_dcpl_460
      OR and_dcpl_468 OR and_dcpl_475 OR and_dcpl_481 OR and_dcpl_486))) OR and_dcpl_495
      OR and_dcpl_500 OR and_dcpl_503 OR and_dcpl_507 OR and_dcpl_510 OR and_dcpl_513;
  COMP_LOOP_COMP_LOOP_or_76_nl <= ((COMP_LOOP_k_9_4_sva_4_0(0)) AND (NOT(and_dcpl_460
      OR and_dcpl_468 OR and_dcpl_495 OR and_dcpl_500 OR and_dcpl_503))) OR and_dcpl_475
      OR and_dcpl_481 OR and_dcpl_486 OR and_dcpl_507 OR and_dcpl_510 OR and_dcpl_513;
  COMP_LOOP_COMP_LOOP_or_77_nl <= (NOT(and_dcpl_453 OR and_dcpl_460 OR and_dcpl_475
      OR and_dcpl_481 OR and_dcpl_495 OR and_dcpl_500 OR and_dcpl_507 OR and_dcpl_510))
      OR and_dcpl_468 OR and_dcpl_486 OR and_dcpl_503 OR and_dcpl_513;
  COMP_LOOP_COMP_LOOP_or_78_nl <= (NOT(and_dcpl_468 OR and_dcpl_475 OR and_dcpl_486
      OR and_dcpl_495 OR and_dcpl_503 OR and_dcpl_507 OR and_dcpl_513)) OR and_dcpl_453
      OR and_dcpl_460 OR and_dcpl_481 OR and_dcpl_500 OR and_dcpl_510;
  acc_3_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_COMP_LOOP_or_74_nl
      & COMP_LOOP_COMP_LOOP_mux_18_nl & COMP_LOOP_or_70_nl) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_COMP_LOOP_mux_19_nl
      & COMP_LOOP_COMP_LOOP_or_75_nl & COMP_LOOP_COMP_LOOP_or_76_nl & COMP_LOOP_COMP_LOOP_or_77_nl
      & COMP_LOOP_COMP_LOOP_or_78_nl & '1'), 10), 11), 11));
  z_out_3 <= acc_3_nl(10 DOWNTO 1);
  COMP_LOOP_mux_82_nl <= MUX_v_10_2_2((VEC_LOOP_j_sva_11_0(11 DOWNTO 2)), STAGE_LOOP_lshift_psp_sva,
      COMP_LOOP_or_24_itm);
  COMP_LOOP_COMP_LOOP_mux_20_nl <= MUX_v_5_2_2((STD_LOGIC_VECTOR'( "00") & (COMP_LOOP_k_9_4_sva_4_0(4
      DOWNTO 2))), COMP_LOOP_k_9_4_sva_4_0, COMP_LOOP_or_24_itm);
  COMP_LOOP_COMP_LOOP_or_79_nl <= ((COMP_LOOP_k_9_4_sva_4_0(1)) AND (NOT(and_dcpl_531
      OR and_dcpl_540))) OR and_dcpl_544 OR and_dcpl_553 OR and_dcpl_557 OR and_dcpl_561;
  COMP_LOOP_COMP_LOOP_or_80_nl <= ((COMP_LOOP_k_9_4_sva_4_0(0)) AND (NOT(and_dcpl_544
      OR and_dcpl_553))) OR and_dcpl_531 OR and_dcpl_540 OR and_dcpl_557 OR and_dcpl_561;
  COMP_LOOP_COMP_LOOP_or_81_nl <= (NOT(and_dcpl_531 OR and_dcpl_544 OR and_dcpl_557
      OR and_dcpl_561)) OR and_978_ssc OR and_dcpl_540 OR and_dcpl_553;
  COMP_LOOP_COMP_LOOP_or_82_nl <= (NOT(and_dcpl_531 OR and_dcpl_557)) OR and_978_ssc
      OR and_dcpl_540 OR and_dcpl_544 OR and_dcpl_553 OR and_dcpl_561;
  z_out_4 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_mux_82_nl) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_COMP_LOOP_mux_20_nl
      & COMP_LOOP_COMP_LOOP_or_79_nl & COMP_LOOP_COMP_LOOP_or_80_nl & COMP_LOOP_COMP_LOOP_or_81_nl
      & COMP_LOOP_COMP_LOOP_or_82_nl), 9), 10), 10));
  and_1178_nl <= and_dcpl_569 AND and_dcpl_567 AND and_827_cse AND and_825_cse;
  and_1179_nl <= and_dcpl_569 AND and_dcpl_383 AND and_835_cse AND (NOT (fsm_output(6)))
      AND (NOT (fsm_output(0)));
  and_1180_nl <= and_dcpl_472 AND (NOT (fsm_output(10))) AND and_dcpl_114 AND (fsm_output(8))
      AND and_dcpl_371 AND (fsm_output(1)) AND (NOT (fsm_output(6))) AND (fsm_output(0));
  and_1181_nl <= and_dcpl_594 AND and_dcpl_114 AND (NOT (fsm_output(8))) AND (fsm_output(4))
      AND (NOT (fsm_output(7))) AND (NOT (fsm_output(1))) AND and_825_cse;
  and_1182_nl <= and_dcpl_594 AND and_dcpl_567 AND and_827_cse AND and_815_cse;
  and_1183_nl <= and_dcpl_568 AND (fsm_output(10)) AND and_dcpl_338 AND and_835_cse
      AND and_815_cse;
  and_1184_nl <= and_dcpl_472 AND (fsm_output(10)) AND and_dcpl_383 AND (fsm_output(4))
      AND (fsm_output(7)) AND (NOT (fsm_output(1))) AND and_815_cse;
  COMP_LOOP_mux1h_578_nl <= MUX1HOT_v_4_7_2(STD_LOGIC_VECTOR'( "0001"), STD_LOGIC_VECTOR'(
      "0010"), STD_LOGIC_VECTOR'( "0011"), STD_LOGIC_VECTOR'( "0101"), STD_LOGIC_VECTOR'(
      "0110"), STD_LOGIC_VECTOR'( "1010"), STD_LOGIC_VECTOR'( "1110"), STD_LOGIC_VECTOR'(
      and_1178_nl & and_1179_nl & and_1180_nl & and_1181_nl & and_1182_nl & and_1183_nl
      & and_1184_nl));
  and_1185_nl <= (NOT (fsm_output(2))) AND (fsm_output(9)) AND (fsm_output(10)) AND
      and_dcpl_338 AND and_dcpl_344 AND (fsm_output(1)) AND and_825_cse;
  COMP_LOOP_or_71_nl <= MUX_v_4_2_2(COMP_LOOP_mux1h_578_nl, STD_LOGIC_VECTOR'("1111"),
      and_1185_nl);
  z_out_5 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(STAGE_LOOP_lshift_psp_sva) +
      CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0 & COMP_LOOP_or_71_nl),
      9), 10), 10));
  COMP_LOOP_COMP_LOOP_or_83_nl <= ((p_sva(63)) AND COMP_LOOP_nor_633_itm) OR not_tmp_838
      OR and_dcpl_650;
  COMP_LOOP_COMP_LOOP_or_84_nl <= ((p_sva(62)) AND COMP_LOOP_nor_633_itm) OR not_tmp_838
      OR and_dcpl_650;
  COMP_LOOP_COMP_LOOP_or_85_nl <= ((p_sva(61)) AND COMP_LOOP_nor_633_itm) OR not_tmp_838
      OR and_dcpl_650;
  COMP_LOOP_COMP_LOOP_or_86_nl <= ((p_sva(60)) AND COMP_LOOP_nor_633_itm) OR not_tmp_838
      OR and_dcpl_650;
  COMP_LOOP_COMP_LOOP_or_87_nl <= ((p_sva(59)) AND COMP_LOOP_nor_633_itm) OR not_tmp_838
      OR and_dcpl_650;
  COMP_LOOP_COMP_LOOP_or_88_nl <= ((p_sva(58)) AND COMP_LOOP_nor_633_itm) OR not_tmp_838
      OR and_dcpl_650;
  COMP_LOOP_COMP_LOOP_or_89_nl <= ((p_sva(57)) AND COMP_LOOP_nor_633_itm) OR not_tmp_838
      OR and_dcpl_650;
  COMP_LOOP_COMP_LOOP_or_90_nl <= ((p_sva(56)) AND COMP_LOOP_nor_633_itm) OR not_tmp_838
      OR and_dcpl_650;
  COMP_LOOP_COMP_LOOP_or_91_nl <= ((p_sva(55)) AND COMP_LOOP_nor_633_itm) OR not_tmp_838
      OR and_dcpl_650;
  COMP_LOOP_COMP_LOOP_or_92_nl <= ((p_sva(54)) AND COMP_LOOP_nor_633_itm) OR not_tmp_838
      OR and_dcpl_650;
  COMP_LOOP_COMP_LOOP_or_93_nl <= ((p_sva(53)) AND COMP_LOOP_nor_633_itm) OR not_tmp_838
      OR and_dcpl_650;
  COMP_LOOP_COMP_LOOP_or_94_nl <= ((p_sva(52)) AND COMP_LOOP_nor_633_itm) OR not_tmp_838
      OR and_dcpl_650;
  COMP_LOOP_COMP_LOOP_or_95_nl <= ((p_sva(51)) AND COMP_LOOP_nor_633_itm) OR not_tmp_838
      OR and_dcpl_650;
  COMP_LOOP_COMP_LOOP_or_96_nl <= ((p_sva(50)) AND COMP_LOOP_nor_633_itm) OR not_tmp_838
      OR and_dcpl_650;
  COMP_LOOP_COMP_LOOP_or_97_nl <= ((p_sva(49)) AND COMP_LOOP_nor_633_itm) OR not_tmp_838
      OR and_dcpl_650;
  COMP_LOOP_COMP_LOOP_or_98_nl <= ((p_sva(48)) AND COMP_LOOP_nor_633_itm) OR not_tmp_838
      OR and_dcpl_650;
  COMP_LOOP_COMP_LOOP_or_99_nl <= ((p_sva(47)) AND COMP_LOOP_nor_633_itm) OR not_tmp_838
      OR and_dcpl_650;
  COMP_LOOP_COMP_LOOP_or_100_nl <= ((p_sva(46)) AND COMP_LOOP_nor_633_itm) OR not_tmp_838
      OR and_dcpl_650;
  COMP_LOOP_COMP_LOOP_or_101_nl <= ((p_sva(45)) AND COMP_LOOP_nor_633_itm) OR not_tmp_838
      OR and_dcpl_650;
  COMP_LOOP_COMP_LOOP_or_102_nl <= ((p_sva(44)) AND COMP_LOOP_nor_633_itm) OR not_tmp_838
      OR and_dcpl_650;
  COMP_LOOP_COMP_LOOP_or_103_nl <= ((p_sva(43)) AND COMP_LOOP_nor_633_itm) OR not_tmp_838
      OR and_dcpl_650;
  COMP_LOOP_COMP_LOOP_or_104_nl <= ((p_sva(42)) AND COMP_LOOP_nor_633_itm) OR not_tmp_838
      OR and_dcpl_650;
  COMP_LOOP_COMP_LOOP_or_105_nl <= ((p_sva(41)) AND COMP_LOOP_nor_633_itm) OR not_tmp_838
      OR and_dcpl_650;
  COMP_LOOP_COMP_LOOP_or_106_nl <= ((p_sva(40)) AND COMP_LOOP_nor_633_itm) OR not_tmp_838
      OR and_dcpl_650;
  COMP_LOOP_COMP_LOOP_or_107_nl <= ((p_sva(39)) AND COMP_LOOP_nor_633_itm) OR not_tmp_838
      OR and_dcpl_650;
  COMP_LOOP_COMP_LOOP_or_108_nl <= ((p_sva(38)) AND COMP_LOOP_nor_633_itm) OR not_tmp_838
      OR and_dcpl_650;
  COMP_LOOP_COMP_LOOP_or_109_nl <= ((p_sva(37)) AND COMP_LOOP_nor_633_itm) OR not_tmp_838
      OR and_dcpl_650;
  COMP_LOOP_COMP_LOOP_or_110_nl <= ((p_sva(36)) AND COMP_LOOP_nor_633_itm) OR not_tmp_838
      OR and_dcpl_650;
  COMP_LOOP_COMP_LOOP_or_111_nl <= ((p_sva(35)) AND COMP_LOOP_nor_633_itm) OR not_tmp_838
      OR and_dcpl_650;
  COMP_LOOP_COMP_LOOP_or_112_nl <= ((p_sva(34)) AND COMP_LOOP_nor_633_itm) OR not_tmp_838
      OR and_dcpl_650;
  COMP_LOOP_COMP_LOOP_or_113_nl <= ((p_sva(33)) AND COMP_LOOP_nor_633_itm) OR not_tmp_838
      OR and_dcpl_650;
  COMP_LOOP_COMP_LOOP_or_114_nl <= ((p_sva(32)) AND COMP_LOOP_nor_633_itm) OR not_tmp_838
      OR and_dcpl_650;
  COMP_LOOP_COMP_LOOP_or_115_nl <= ((p_sva(31)) AND COMP_LOOP_nor_633_itm) OR not_tmp_838
      OR and_dcpl_650;
  COMP_LOOP_COMP_LOOP_or_116_nl <= ((p_sva(30)) AND COMP_LOOP_nor_633_itm) OR not_tmp_838
      OR and_dcpl_650;
  COMP_LOOP_COMP_LOOP_or_117_nl <= ((p_sva(29)) AND COMP_LOOP_nor_633_itm) OR not_tmp_838
      OR and_dcpl_650;
  COMP_LOOP_COMP_LOOP_or_118_nl <= ((p_sva(28)) AND COMP_LOOP_nor_633_itm) OR not_tmp_838
      OR and_dcpl_650;
  COMP_LOOP_COMP_LOOP_or_119_nl <= ((p_sva(27)) AND COMP_LOOP_nor_633_itm) OR not_tmp_838
      OR and_dcpl_650;
  COMP_LOOP_COMP_LOOP_or_120_nl <= ((p_sva(26)) AND COMP_LOOP_nor_633_itm) OR not_tmp_838
      OR and_dcpl_650;
  COMP_LOOP_COMP_LOOP_or_121_nl <= ((p_sva(25)) AND COMP_LOOP_nor_633_itm) OR not_tmp_838
      OR and_dcpl_650;
  COMP_LOOP_COMP_LOOP_or_122_nl <= ((p_sva(24)) AND COMP_LOOP_nor_633_itm) OR not_tmp_838
      OR and_dcpl_650;
  COMP_LOOP_COMP_LOOP_or_123_nl <= ((p_sva(23)) AND COMP_LOOP_nor_633_itm) OR not_tmp_838
      OR and_dcpl_650;
  COMP_LOOP_COMP_LOOP_or_124_nl <= ((p_sva(22)) AND COMP_LOOP_nor_633_itm) OR not_tmp_838
      OR and_dcpl_650;
  COMP_LOOP_COMP_LOOP_or_125_nl <= ((p_sva(21)) AND COMP_LOOP_nor_633_itm) OR not_tmp_838
      OR and_dcpl_650;
  COMP_LOOP_COMP_LOOP_or_126_nl <= ((p_sva(20)) AND COMP_LOOP_nor_633_itm) OR not_tmp_838
      OR and_dcpl_650;
  COMP_LOOP_COMP_LOOP_or_127_nl <= ((p_sva(19)) AND COMP_LOOP_nor_633_itm) OR not_tmp_838
      OR and_dcpl_650;
  COMP_LOOP_COMP_LOOP_or_128_nl <= ((p_sva(18)) AND COMP_LOOP_nor_633_itm) OR not_tmp_838
      OR and_dcpl_650;
  COMP_LOOP_COMP_LOOP_or_129_nl <= ((p_sva(17)) AND COMP_LOOP_nor_633_itm) OR not_tmp_838
      OR and_dcpl_650;
  COMP_LOOP_COMP_LOOP_or_130_nl <= ((p_sva(16)) AND COMP_LOOP_nor_633_itm) OR not_tmp_838
      OR and_dcpl_650;
  COMP_LOOP_COMP_LOOP_or_131_nl <= ((p_sva(15)) AND COMP_LOOP_nor_633_itm) OR not_tmp_838
      OR and_dcpl_650;
  COMP_LOOP_COMP_LOOP_or_132_nl <= ((p_sva(14)) AND COMP_LOOP_nor_633_itm) OR not_tmp_838
      OR and_dcpl_650;
  COMP_LOOP_COMP_LOOP_or_133_nl <= ((p_sva(13)) AND COMP_LOOP_nor_633_itm) OR not_tmp_838
      OR and_dcpl_650;
  COMP_LOOP_COMP_LOOP_or_134_nl <= ((p_sva(12)) AND COMP_LOOP_nor_633_itm) OR not_tmp_838
      OR and_dcpl_650;
  COMP_LOOP_mux_83_nl <= MUX_v_4_2_2((VEC_LOOP_j_sva_11_0(11 DOWNTO 8)), (p_sva(11
      DOWNTO 8)), and_dcpl_647);
  COMP_LOOP_and_398_nl <= MUX_v_4_2_2(STD_LOGIC_VECTOR'("0000"), COMP_LOOP_mux_83_nl,
      COMP_LOOP_nor_685_itm);
  COMP_LOOP_or_72_nl <= not_tmp_838 OR and_dcpl_650;
  COMP_LOOP_COMP_LOOP_or_135_nl <= MUX_v_4_2_2(COMP_LOOP_and_398_nl, STD_LOGIC_VECTOR'("1111"),
      COMP_LOOP_or_72_nl);
  COMP_LOOP_mux1h_579_nl <= MUX1HOT_s_1_4_2((VEC_LOOP_j_sva_11_0(7)), (NOT modExp_exp_1_7_1_sva),
      (p_sva(7)), (NOT COMP_LOOP_nor_134_itm), STD_LOGIC_VECTOR'( and_dcpl_628 &
      not_tmp_838 & and_dcpl_647 & and_dcpl_650));
  COMP_LOOP_or_73_nl <= COMP_LOOP_mux1h_579_nl OR and_dcpl_636 OR and_dcpl_642;
  COMP_LOOP_mux1h_580_nl <= MUX1HOT_v_7_5_2((VEC_LOOP_j_sva_11_0(6 DOWNTO 0)), (NOT
      (STAGE_LOOP_lshift_psp_sva(9 DOWNTO 3))), STD_LOGIC_VECTOR'( (NOT modExp_exp_1_6_1_sva)
      & (NOT modExp_exp_1_5_1_sva) & (NOT modExp_exp_1_4_1_sva) & (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      & (NOT COMP_LOOP_nor_137_itm) & (NOT COMP_LOOP_nor_134_itm) & (NOT COMP_LOOP_nor_12_itm)),
      (p_sva(6 DOWNTO 0)), STD_LOGIC_VECTOR'( (NOT modExp_exp_1_7_1_sva) & (NOT modExp_exp_1_6_1_sva)
      & (NOT modExp_exp_1_5_1_sva) & (NOT modExp_exp_1_4_1_sva) & (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      & (NOT COMP_LOOP_nor_137_itm) & (NOT COMP_LOOP_nor_12_itm)), STD_LOGIC_VECTOR'(
      and_dcpl_628 & COMP_LOOP_or_65_itm & not_tmp_838 & and_dcpl_647 & and_dcpl_650));
  COMP_LOOP_or_74_nl <= (NOT(and_dcpl_628 OR not_tmp_838 OR and_dcpl_647 OR and_dcpl_650))
      OR and_dcpl_636 OR and_dcpl_642;
  COMP_LOOP_COMP_LOOP_or_136_nl <= (NOT(and_dcpl_628 OR and_dcpl_636 OR and_dcpl_642
      OR not_tmp_838 OR and_dcpl_650)) OR and_dcpl_647;
  COMP_LOOP_COMP_LOOP_or_137_nl <= ((COMP_LOOP_k_9_4_sva_4_0(4)) AND COMP_LOOP_nor_687_itm)
      OR and_dcpl_647;
  COMP_LOOP_COMP_LOOP_or_138_nl <= ((COMP_LOOP_k_9_4_sva_4_0(3)) AND COMP_LOOP_nor_687_itm)
      OR and_dcpl_647;
  COMP_LOOP_COMP_LOOP_mux_21_nl <= MUX_v_3_2_2((COMP_LOOP_k_9_4_sva_4_0(2 DOWNTO
      0)), (COMP_LOOP_k_9_4_sva_4_0(4 DOWNTO 2)), COMP_LOOP_or_65_itm);
  COMP_LOOP_nor_706_nl <= NOT(not_tmp_838 OR and_dcpl_650);
  COMP_LOOP_and_401_nl <= MUX_v_3_2_2(STD_LOGIC_VECTOR'("000"), COMP_LOOP_COMP_LOOP_mux_21_nl,
      COMP_LOOP_nor_706_nl);
  COMP_LOOP_or_75_nl <= MUX_v_3_2_2(COMP_LOOP_and_401_nl, STD_LOGIC_VECTOR'("111"),
      and_dcpl_647);
  COMP_LOOP_nor_707_nl <= NOT(and_dcpl_628 OR not_tmp_838 OR and_dcpl_650);
  COMP_LOOP_and_402_nl <= MUX_v_2_2_2(STD_LOGIC_VECTOR'("00"), (COMP_LOOP_k_9_4_sva_4_0(1
      DOWNTO 0)), COMP_LOOP_nor_707_nl);
  COMP_LOOP_COMP_LOOP_or_139_nl <= MUX_v_2_2_2(COMP_LOOP_and_402_nl, STD_LOGIC_VECTOR'("11"),
      and_dcpl_647);
  COMP_LOOP_COMP_LOOP_or_140_nl <= (NOT(and_dcpl_636 OR not_tmp_838 OR and_dcpl_650))
      OR and_dcpl_628 OR and_dcpl_642 OR and_dcpl_647;
  COMP_LOOP_COMP_LOOP_or_141_nl <= COMP_LOOP_nor_685_itm OR and_dcpl_628 OR not_tmp_838
      OR and_dcpl_647 OR and_dcpl_650;
  acc_6_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_COMP_LOOP_or_83_nl
      & COMP_LOOP_COMP_LOOP_or_84_nl & COMP_LOOP_COMP_LOOP_or_85_nl & COMP_LOOP_COMP_LOOP_or_86_nl
      & COMP_LOOP_COMP_LOOP_or_87_nl & COMP_LOOP_COMP_LOOP_or_88_nl & COMP_LOOP_COMP_LOOP_or_89_nl
      & COMP_LOOP_COMP_LOOP_or_90_nl & COMP_LOOP_COMP_LOOP_or_91_nl & COMP_LOOP_COMP_LOOP_or_92_nl
      & COMP_LOOP_COMP_LOOP_or_93_nl & COMP_LOOP_COMP_LOOP_or_94_nl & COMP_LOOP_COMP_LOOP_or_95_nl
      & COMP_LOOP_COMP_LOOP_or_96_nl & COMP_LOOP_COMP_LOOP_or_97_nl & COMP_LOOP_COMP_LOOP_or_98_nl
      & COMP_LOOP_COMP_LOOP_or_99_nl & COMP_LOOP_COMP_LOOP_or_100_nl & COMP_LOOP_COMP_LOOP_or_101_nl
      & COMP_LOOP_COMP_LOOP_or_102_nl & COMP_LOOP_COMP_LOOP_or_103_nl & COMP_LOOP_COMP_LOOP_or_104_nl
      & COMP_LOOP_COMP_LOOP_or_105_nl & COMP_LOOP_COMP_LOOP_or_106_nl & COMP_LOOP_COMP_LOOP_or_107_nl
      & COMP_LOOP_COMP_LOOP_or_108_nl & COMP_LOOP_COMP_LOOP_or_109_nl & COMP_LOOP_COMP_LOOP_or_110_nl
      & COMP_LOOP_COMP_LOOP_or_111_nl & COMP_LOOP_COMP_LOOP_or_112_nl & COMP_LOOP_COMP_LOOP_or_113_nl
      & COMP_LOOP_COMP_LOOP_or_114_nl & COMP_LOOP_COMP_LOOP_or_115_nl & COMP_LOOP_COMP_LOOP_or_116_nl
      & COMP_LOOP_COMP_LOOP_or_117_nl & COMP_LOOP_COMP_LOOP_or_118_nl & COMP_LOOP_COMP_LOOP_or_119_nl
      & COMP_LOOP_COMP_LOOP_or_120_nl & COMP_LOOP_COMP_LOOP_or_121_nl & COMP_LOOP_COMP_LOOP_or_122_nl
      & COMP_LOOP_COMP_LOOP_or_123_nl & COMP_LOOP_COMP_LOOP_or_124_nl & COMP_LOOP_COMP_LOOP_or_125_nl
      & COMP_LOOP_COMP_LOOP_or_126_nl & COMP_LOOP_COMP_LOOP_or_127_nl & COMP_LOOP_COMP_LOOP_or_128_nl
      & COMP_LOOP_COMP_LOOP_or_129_nl & COMP_LOOP_COMP_LOOP_or_130_nl & COMP_LOOP_COMP_LOOP_or_131_nl
      & COMP_LOOP_COMP_LOOP_or_132_nl & COMP_LOOP_COMP_LOOP_or_133_nl & COMP_LOOP_COMP_LOOP_or_134_nl
      & COMP_LOOP_COMP_LOOP_or_135_nl & COMP_LOOP_or_73_nl & COMP_LOOP_mux1h_580_nl
      & COMP_LOOP_or_74_nl), 65), 66) + CONV_UNSIGNED(CONV_SIGNED(SIGNED(COMP_LOOP_COMP_LOOP_or_136_nl
      & COMP_LOOP_COMP_LOOP_or_137_nl & COMP_LOOP_COMP_LOOP_or_138_nl & COMP_LOOP_or_75_nl
      & COMP_LOOP_COMP_LOOP_or_139_nl & COMP_LOOP_COMP_LOOP_or_140_nl & COMP_LOOP_COMP_LOOP_or_141_nl
      & '1'), 11), 66), 66));
  z_out_6 <= acc_6_nl(65 DOWNTO 1);
  COMP_LOOP_COMP_LOOP_or_142_nl <= ((STAGE_LOOP_lshift_psp_sva(9)) AND (NOT(and_dcpl_669
      OR and_dcpl_678))) OR and_dcpl_660;
  COMP_LOOP_mux1h_581_nl <= MUX1HOT_v_6_4_2((NOT (STAGE_LOOP_lshift_psp_sva(9 DOWNTO
      4))), ('1' & (NOT (STAGE_LOOP_lshift_psp_sva(9 DOWNTO 5)))), (STAGE_LOOP_lshift_psp_sva(9
      DOWNTO 4)), (STAGE_LOOP_lshift_psp_sva(8 DOWNTO 3)), STD_LOGIC_VECTOR'( and_dcpl_660
      & and_dcpl_669 & and_dcpl_678 & and_dcpl_686));
  COMP_LOOP_or_76_nl <= (NOT(and_dcpl_678 OR and_dcpl_686)) OR and_dcpl_660 OR and_dcpl_669;
  COMP_LOOP_or_77_nl <= and_dcpl_669 OR and_dcpl_678;
  COMP_LOOP_COMP_LOOP_mux_22_nl <= MUX_v_5_2_2(COMP_LOOP_k_9_4_sva_4_0, ('0' & (COMP_LOOP_k_9_4_sva_4_0(4
      DOWNTO 1))), COMP_LOOP_or_77_nl);
  COMP_LOOP_COMP_LOOP_or_143_nl <= ((COMP_LOOP_k_9_4_sva_4_0(0)) AND (NOT and_dcpl_660))
      OR and_dcpl_686;
  acc_7_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_COMP_LOOP_or_142_nl
      & COMP_LOOP_mux1h_581_nl & COMP_LOOP_or_76_nl) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_COMP_LOOP_mux_22_nl
      & COMP_LOOP_COMP_LOOP_or_143_nl & '1'), 7), 8), 8));
  z_out_7 <= acc_7_nl(7 DOWNTO 1);
  mux_3950_nl <= MUX_s_1_2_2(or_tmp_3307, or_tmp_3326, fsm_output(0));
  or_3639_nl <= (NOT (fsm_output(8))) OR (fsm_output(6)) OR mux_3950_nl;
  or_3640_nl <= (fsm_output(8)) OR (fsm_output(6)) OR (NOT (fsm_output(0))) OR (fsm_output(9))
      OR (fsm_output(10)) OR (NOT (fsm_output(1))) OR (fsm_output(2));
  mux_3949_nl <= MUX_s_1_2_2(or_3639_nl, or_3640_nl, fsm_output(3));
  nor_1711_nl <= NOT((fsm_output(4)) OR mux_3949_nl);
  mux_3952_nl <= MUX_s_1_2_2(or_tmp_3326, or_tmp_3312, fsm_output(0));
  and_1186_nl <= (fsm_output(3)) AND (fsm_output(8)) AND (fsm_output(6)) AND (NOT
      mux_3952_nl);
  or_3641_nl <= (fsm_output(10)) OR (fsm_output(1)) OR (NOT (fsm_output(2)));
  or_3642_nl <= (fsm_output(10)) OR (NOT and_529_cse);
  mux_3954_nl <= MUX_s_1_2_2(or_3641_nl, or_3642_nl, fsm_output(9));
  nor_1712_nl <= NOT((fsm_output(8)) OR (fsm_output(6)) OR (fsm_output(0)) OR mux_3954_nl);
  nand_428_nl <= NOT((fsm_output(9)) AND (fsm_output(10)) AND (NOT (fsm_output(1)))
      AND (fsm_output(2)));
  or_3643_nl <= (fsm_output(9)) OR (NOT (fsm_output(10))) OR (fsm_output(1)) OR (fsm_output(2));
  mux_3955_nl <= MUX_s_1_2_2(nand_428_nl, or_3643_nl, fsm_output(0));
  nor_1713_nl <= NOT((fsm_output(8)) OR (fsm_output(6)) OR mux_3955_nl);
  mux_3953_nl <= MUX_s_1_2_2(nor_1712_nl, nor_1713_nl, fsm_output(3));
  mux_3951_nl <= MUX_s_1_2_2(and_1186_nl, mux_3953_nl, fsm_output(4));
  mux_3948_nl <= MUX_s_1_2_2(nor_1711_nl, mux_3951_nl, fsm_output(5));
  and_1187_nl <= (fsm_output(3)) AND (fsm_output(8)) AND (fsm_output(6)) AND (fsm_output(0))
      AND (NOT (fsm_output(9))) AND (NOT (fsm_output(10))) AND and_529_cse;
  or_3644_nl <= (fsm_output(9)) OR (NOT (fsm_output(10))) OR (fsm_output(1)) OR (NOT
      (fsm_output(2)));
  mux_3959_nl <= MUX_s_1_2_2(or_tmp_3312, or_3644_nl, fsm_output(0));
  and_1188_nl <= (fsm_output(8)) AND (fsm_output(6)) AND (NOT mux_3959_nl);
  or_3645_nl <= (fsm_output(9)) OR (fsm_output(10)) OR (NOT (fsm_output(1))) OR (fsm_output(2));
  mux_3960_nl <= MUX_s_1_2_2(or_3645_nl, or_tmp_3307, fsm_output(0));
  nor_1714_nl <= NOT((fsm_output(8)) OR (fsm_output(6)) OR mux_3960_nl);
  mux_3958_nl <= MUX_s_1_2_2(and_1188_nl, nor_1714_nl, fsm_output(3));
  mux_3957_nl <= MUX_s_1_2_2(and_1187_nl, mux_3958_nl, fsm_output(4));
  mux_3956_nl <= MUX_s_1_2_2(mux_3957_nl, nor_1657_cse, fsm_output(5));
  mux_3947_nl <= MUX_s_1_2_2(mux_3948_nl, mux_3956_nl, fsm_output(7));
  modExp_while_if_mux_1_nl <= MUX_v_64_2_2(modExp_result_sva, COMP_LOOP_10_mul_mut,
      mux_3947_nl);
  z_out_8 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(SIGNED'( SIGNED(modExp_while_if_mux_1_nl)
      * SIGNED(COMP_LOOP_10_mul_mut)), 64));
END v44;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    vec_rsc_0_0_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    vec_rsc_0_0_da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_0_wea : OUT STD_LOGIC;
    vec_rsc_0_0_qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_0_lz : OUT STD_LOGIC;
    vec_rsc_0_1_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    vec_rsc_0_1_da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_1_wea : OUT STD_LOGIC;
    vec_rsc_0_1_qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_1_lz : OUT STD_LOGIC;
    vec_rsc_0_2_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    vec_rsc_0_2_da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_2_wea : OUT STD_LOGIC;
    vec_rsc_0_2_qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_2_lz : OUT STD_LOGIC;
    vec_rsc_0_3_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    vec_rsc_0_3_da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_3_wea : OUT STD_LOGIC;
    vec_rsc_0_3_qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_3_lz : OUT STD_LOGIC;
    vec_rsc_0_4_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    vec_rsc_0_4_da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_4_wea : OUT STD_LOGIC;
    vec_rsc_0_4_qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_4_lz : OUT STD_LOGIC;
    vec_rsc_0_5_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    vec_rsc_0_5_da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_5_wea : OUT STD_LOGIC;
    vec_rsc_0_5_qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_5_lz : OUT STD_LOGIC;
    vec_rsc_0_6_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    vec_rsc_0_6_da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_6_wea : OUT STD_LOGIC;
    vec_rsc_0_6_qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_6_lz : OUT STD_LOGIC;
    vec_rsc_0_7_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    vec_rsc_0_7_da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_7_wea : OUT STD_LOGIC;
    vec_rsc_0_7_qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_7_lz : OUT STD_LOGIC;
    vec_rsc_0_8_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    vec_rsc_0_8_da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_8_wea : OUT STD_LOGIC;
    vec_rsc_0_8_qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_8_lz : OUT STD_LOGIC;
    vec_rsc_0_9_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    vec_rsc_0_9_da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_9_wea : OUT STD_LOGIC;
    vec_rsc_0_9_qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_9_lz : OUT STD_LOGIC;
    vec_rsc_0_10_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    vec_rsc_0_10_da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_10_wea : OUT STD_LOGIC;
    vec_rsc_0_10_qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_10_lz : OUT STD_LOGIC;
    vec_rsc_0_11_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    vec_rsc_0_11_da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_11_wea : OUT STD_LOGIC;
    vec_rsc_0_11_qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_11_lz : OUT STD_LOGIC;
    vec_rsc_0_12_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    vec_rsc_0_12_da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_12_wea : OUT STD_LOGIC;
    vec_rsc_0_12_qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_12_lz : OUT STD_LOGIC;
    vec_rsc_0_13_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    vec_rsc_0_13_da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_13_wea : OUT STD_LOGIC;
    vec_rsc_0_13_qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_13_lz : OUT STD_LOGIC;
    vec_rsc_0_14_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    vec_rsc_0_14_da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_14_wea : OUT STD_LOGIC;
    vec_rsc_0_14_qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_14_lz : OUT STD_LOGIC;
    vec_rsc_0_15_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    vec_rsc_0_15_da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_15_wea : OUT STD_LOGIC;
    vec_rsc_0_15_qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_15_lz : OUT STD_LOGIC;
    p_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    p_rsc_triosy_lz : OUT STD_LOGIC;
    r_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    r_rsc_triosy_lz : OUT STD_LOGIC
  );
END inPlaceNTT_DIT;

ARCHITECTURE v44 OF inPlaceNTT_DIT IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';

  -- Interconnect Declarations
  SIGNAL vec_rsc_0_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_1_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_2_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_3_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_4_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_5_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_6_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_7_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_8_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_9_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_10_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_11_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_12_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_13_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_14_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_15_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_0_i_adra_d_iff : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_da_d_iff : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_wea_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_1_i_wea_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_2_i_wea_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_3_i_wea_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_4_i_wea_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_5_i_wea_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_6_i_wea_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_7_i_wea_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_8_i_wea_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_9_i_wea_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_10_i_wea_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_11_i_wea_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_12_i_wea_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_13_i_wea_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_14_i_wea_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_15_i_wea_d_iff : STD_LOGIC;

  COMPONENT inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_4_8_64_256_256_64_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_0_i_qa : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_da : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  COMPONENT inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_5_8_64_256_256_64_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_1_i_qa : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_da : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  COMPONENT inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_6_8_64_256_256_64_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_2_i_qa : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_da : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  COMPONENT inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_7_8_64_256_256_64_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_3_i_qa : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_da : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  COMPONENT inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_8_8_64_256_256_64_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_4_i_qa : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_da : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  COMPONENT inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_9_8_64_256_256_64_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_5_i_qa : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_da : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  COMPONENT inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_10_8_64_256_256_64_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_6_i_qa : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_da : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  COMPONENT inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_11_8_64_256_256_64_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_7_i_qa : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_da : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  COMPONENT inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_12_8_64_256_256_64_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_8_i_qa : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_8_i_da : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_8_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL vec_rsc_0_8_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL vec_rsc_0_8_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_8_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  COMPONENT inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_13_8_64_256_256_64_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_9_i_qa : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_9_i_da : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_9_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL vec_rsc_0_9_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL vec_rsc_0_9_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_9_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  COMPONENT inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_14_8_64_256_256_64_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_10_i_qa : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_10_i_da : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_10_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL vec_rsc_0_10_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL vec_rsc_0_10_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_10_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  COMPONENT inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_15_8_64_256_256_64_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_11_i_qa : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_11_i_da : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_11_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL vec_rsc_0_11_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL vec_rsc_0_11_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_11_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  COMPONENT inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_16_8_64_256_256_64_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_12_i_qa : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_12_i_da : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_12_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL vec_rsc_0_12_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL vec_rsc_0_12_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_12_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  COMPONENT inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_17_8_64_256_256_64_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_13_i_qa : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_13_i_da : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_13_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL vec_rsc_0_13_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL vec_rsc_0_13_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_13_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  COMPONENT inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_18_8_64_256_256_64_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_14_i_qa : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_14_i_da : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_14_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL vec_rsc_0_14_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL vec_rsc_0_14_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_14_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  COMPONENT inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_19_8_64_256_256_64_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_15_i_qa : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_15_i_da : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_15_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL vec_rsc_0_15_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL vec_rsc_0_15_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_15_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  COMPONENT inPlaceNTT_DIT_core
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      vec_rsc_triosy_0_0_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_1_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_2_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_3_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_4_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_5_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_6_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_7_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_8_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_9_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_10_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_11_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_12_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_13_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_14_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_15_lz : OUT STD_LOGIC;
      p_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      p_rsc_triosy_lz : OUT STD_LOGIC;
      r_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      r_rsc_triosy_lz : OUT STD_LOGIC;
      vec_rsc_0_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_1_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_2_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_3_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_4_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_5_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_6_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_7_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_8_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_9_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_10_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_11_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_12_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_13_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_14_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_15_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_0_i_adra_d_pff : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      vec_rsc_0_0_i_da_d_pff : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_0_i_wea_d_pff : OUT STD_LOGIC;
      vec_rsc_0_1_i_wea_d_pff : OUT STD_LOGIC;
      vec_rsc_0_2_i_wea_d_pff : OUT STD_LOGIC;
      vec_rsc_0_3_i_wea_d_pff : OUT STD_LOGIC;
      vec_rsc_0_4_i_wea_d_pff : OUT STD_LOGIC;
      vec_rsc_0_5_i_wea_d_pff : OUT STD_LOGIC;
      vec_rsc_0_6_i_wea_d_pff : OUT STD_LOGIC;
      vec_rsc_0_7_i_wea_d_pff : OUT STD_LOGIC;
      vec_rsc_0_8_i_wea_d_pff : OUT STD_LOGIC;
      vec_rsc_0_9_i_wea_d_pff : OUT STD_LOGIC;
      vec_rsc_0_10_i_wea_d_pff : OUT STD_LOGIC;
      vec_rsc_0_11_i_wea_d_pff : OUT STD_LOGIC;
      vec_rsc_0_12_i_wea_d_pff : OUT STD_LOGIC;
      vec_rsc_0_13_i_wea_d_pff : OUT STD_LOGIC;
      vec_rsc_0_14_i_wea_d_pff : OUT STD_LOGIC;
      vec_rsc_0_15_i_wea_d_pff : OUT STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIT_core_inst_p_rsc_dat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIT_core_inst_r_rsc_dat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIT_core_inst_vec_rsc_0_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIT_core_inst_vec_rsc_0_1_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIT_core_inst_vec_rsc_0_2_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIT_core_inst_vec_rsc_0_3_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIT_core_inst_vec_rsc_0_4_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIT_core_inst_vec_rsc_0_5_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIT_core_inst_vec_rsc_0_6_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIT_core_inst_vec_rsc_0_7_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIT_core_inst_vec_rsc_0_8_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIT_core_inst_vec_rsc_0_9_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIT_core_inst_vec_rsc_0_10_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIT_core_inst_vec_rsc_0_11_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIT_core_inst_vec_rsc_0_12_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIT_core_inst_vec_rsc_0_13_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIT_core_inst_vec_rsc_0_14_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIT_core_inst_vec_rsc_0_15_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIT_core_inst_vec_rsc_0_0_i_adra_d_pff : STD_LOGIC_VECTOR (7
      DOWNTO 0);
  SIGNAL inPlaceNTT_DIT_core_inst_vec_rsc_0_0_i_da_d_pff : STD_LOGIC_VECTOR (63 DOWNTO
      0);

BEGIN
  vec_rsc_0_0_i : inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_4_8_64_256_256_64_1_gen
    PORT MAP(
      qa => vec_rsc_0_0_i_qa,
      wea => vec_rsc_0_0_wea,
      da => vec_rsc_0_0_i_da,
      adra => vec_rsc_0_0_i_adra,
      adra_d => vec_rsc_0_0_i_adra_d,
      da_d => vec_rsc_0_0_i_da_d,
      qa_d => vec_rsc_0_0_i_qa_d_1,
      wea_d => vec_rsc_0_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_0_0_i_wea_d_iff
    );
  vec_rsc_0_0_i_qa <= vec_rsc_0_0_qa;
  vec_rsc_0_0_da <= vec_rsc_0_0_i_da;
  vec_rsc_0_0_adra <= vec_rsc_0_0_i_adra;
  vec_rsc_0_0_i_adra_d <= vec_rsc_0_0_i_adra_d_iff;
  vec_rsc_0_0_i_da_d <= vec_rsc_0_0_i_da_d_iff;
  vec_rsc_0_0_i_qa_d <= vec_rsc_0_0_i_qa_d_1;

  vec_rsc_0_1_i : inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_5_8_64_256_256_64_1_gen
    PORT MAP(
      qa => vec_rsc_0_1_i_qa,
      wea => vec_rsc_0_1_wea,
      da => vec_rsc_0_1_i_da,
      adra => vec_rsc_0_1_i_adra,
      adra_d => vec_rsc_0_1_i_adra_d,
      da_d => vec_rsc_0_1_i_da_d,
      qa_d => vec_rsc_0_1_i_qa_d_1,
      wea_d => vec_rsc_0_1_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_0_1_i_wea_d_iff
    );
  vec_rsc_0_1_i_qa <= vec_rsc_0_1_qa;
  vec_rsc_0_1_da <= vec_rsc_0_1_i_da;
  vec_rsc_0_1_adra <= vec_rsc_0_1_i_adra;
  vec_rsc_0_1_i_adra_d <= vec_rsc_0_0_i_adra_d_iff;
  vec_rsc_0_1_i_da_d <= vec_rsc_0_0_i_da_d_iff;
  vec_rsc_0_1_i_qa_d <= vec_rsc_0_1_i_qa_d_1;

  vec_rsc_0_2_i : inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_6_8_64_256_256_64_1_gen
    PORT MAP(
      qa => vec_rsc_0_2_i_qa,
      wea => vec_rsc_0_2_wea,
      da => vec_rsc_0_2_i_da,
      adra => vec_rsc_0_2_i_adra,
      adra_d => vec_rsc_0_2_i_adra_d,
      da_d => vec_rsc_0_2_i_da_d,
      qa_d => vec_rsc_0_2_i_qa_d_1,
      wea_d => vec_rsc_0_2_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_0_2_i_wea_d_iff
    );
  vec_rsc_0_2_i_qa <= vec_rsc_0_2_qa;
  vec_rsc_0_2_da <= vec_rsc_0_2_i_da;
  vec_rsc_0_2_adra <= vec_rsc_0_2_i_adra;
  vec_rsc_0_2_i_adra_d <= vec_rsc_0_0_i_adra_d_iff;
  vec_rsc_0_2_i_da_d <= vec_rsc_0_0_i_da_d_iff;
  vec_rsc_0_2_i_qa_d <= vec_rsc_0_2_i_qa_d_1;

  vec_rsc_0_3_i : inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_7_8_64_256_256_64_1_gen
    PORT MAP(
      qa => vec_rsc_0_3_i_qa,
      wea => vec_rsc_0_3_wea,
      da => vec_rsc_0_3_i_da,
      adra => vec_rsc_0_3_i_adra,
      adra_d => vec_rsc_0_3_i_adra_d,
      da_d => vec_rsc_0_3_i_da_d,
      qa_d => vec_rsc_0_3_i_qa_d_1,
      wea_d => vec_rsc_0_3_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_0_3_i_wea_d_iff
    );
  vec_rsc_0_3_i_qa <= vec_rsc_0_3_qa;
  vec_rsc_0_3_da <= vec_rsc_0_3_i_da;
  vec_rsc_0_3_adra <= vec_rsc_0_3_i_adra;
  vec_rsc_0_3_i_adra_d <= vec_rsc_0_0_i_adra_d_iff;
  vec_rsc_0_3_i_da_d <= vec_rsc_0_0_i_da_d_iff;
  vec_rsc_0_3_i_qa_d <= vec_rsc_0_3_i_qa_d_1;

  vec_rsc_0_4_i : inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_8_8_64_256_256_64_1_gen
    PORT MAP(
      qa => vec_rsc_0_4_i_qa,
      wea => vec_rsc_0_4_wea,
      da => vec_rsc_0_4_i_da,
      adra => vec_rsc_0_4_i_adra,
      adra_d => vec_rsc_0_4_i_adra_d,
      da_d => vec_rsc_0_4_i_da_d,
      qa_d => vec_rsc_0_4_i_qa_d_1,
      wea_d => vec_rsc_0_4_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_0_4_i_wea_d_iff
    );
  vec_rsc_0_4_i_qa <= vec_rsc_0_4_qa;
  vec_rsc_0_4_da <= vec_rsc_0_4_i_da;
  vec_rsc_0_4_adra <= vec_rsc_0_4_i_adra;
  vec_rsc_0_4_i_adra_d <= vec_rsc_0_0_i_adra_d_iff;
  vec_rsc_0_4_i_da_d <= vec_rsc_0_0_i_da_d_iff;
  vec_rsc_0_4_i_qa_d <= vec_rsc_0_4_i_qa_d_1;

  vec_rsc_0_5_i : inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_9_8_64_256_256_64_1_gen
    PORT MAP(
      qa => vec_rsc_0_5_i_qa,
      wea => vec_rsc_0_5_wea,
      da => vec_rsc_0_5_i_da,
      adra => vec_rsc_0_5_i_adra,
      adra_d => vec_rsc_0_5_i_adra_d,
      da_d => vec_rsc_0_5_i_da_d,
      qa_d => vec_rsc_0_5_i_qa_d_1,
      wea_d => vec_rsc_0_5_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_0_5_i_wea_d_iff
    );
  vec_rsc_0_5_i_qa <= vec_rsc_0_5_qa;
  vec_rsc_0_5_da <= vec_rsc_0_5_i_da;
  vec_rsc_0_5_adra <= vec_rsc_0_5_i_adra;
  vec_rsc_0_5_i_adra_d <= vec_rsc_0_0_i_adra_d_iff;
  vec_rsc_0_5_i_da_d <= vec_rsc_0_0_i_da_d_iff;
  vec_rsc_0_5_i_qa_d <= vec_rsc_0_5_i_qa_d_1;

  vec_rsc_0_6_i : inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_10_8_64_256_256_64_1_gen
    PORT MAP(
      qa => vec_rsc_0_6_i_qa,
      wea => vec_rsc_0_6_wea,
      da => vec_rsc_0_6_i_da,
      adra => vec_rsc_0_6_i_adra,
      adra_d => vec_rsc_0_6_i_adra_d,
      da_d => vec_rsc_0_6_i_da_d,
      qa_d => vec_rsc_0_6_i_qa_d_1,
      wea_d => vec_rsc_0_6_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_0_6_i_wea_d_iff
    );
  vec_rsc_0_6_i_qa <= vec_rsc_0_6_qa;
  vec_rsc_0_6_da <= vec_rsc_0_6_i_da;
  vec_rsc_0_6_adra <= vec_rsc_0_6_i_adra;
  vec_rsc_0_6_i_adra_d <= vec_rsc_0_0_i_adra_d_iff;
  vec_rsc_0_6_i_da_d <= vec_rsc_0_0_i_da_d_iff;
  vec_rsc_0_6_i_qa_d <= vec_rsc_0_6_i_qa_d_1;

  vec_rsc_0_7_i : inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_11_8_64_256_256_64_1_gen
    PORT MAP(
      qa => vec_rsc_0_7_i_qa,
      wea => vec_rsc_0_7_wea,
      da => vec_rsc_0_7_i_da,
      adra => vec_rsc_0_7_i_adra,
      adra_d => vec_rsc_0_7_i_adra_d,
      da_d => vec_rsc_0_7_i_da_d,
      qa_d => vec_rsc_0_7_i_qa_d_1,
      wea_d => vec_rsc_0_7_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_0_7_i_wea_d_iff
    );
  vec_rsc_0_7_i_qa <= vec_rsc_0_7_qa;
  vec_rsc_0_7_da <= vec_rsc_0_7_i_da;
  vec_rsc_0_7_adra <= vec_rsc_0_7_i_adra;
  vec_rsc_0_7_i_adra_d <= vec_rsc_0_0_i_adra_d_iff;
  vec_rsc_0_7_i_da_d <= vec_rsc_0_0_i_da_d_iff;
  vec_rsc_0_7_i_qa_d <= vec_rsc_0_7_i_qa_d_1;

  vec_rsc_0_8_i : inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_12_8_64_256_256_64_1_gen
    PORT MAP(
      qa => vec_rsc_0_8_i_qa,
      wea => vec_rsc_0_8_wea,
      da => vec_rsc_0_8_i_da,
      adra => vec_rsc_0_8_i_adra,
      adra_d => vec_rsc_0_8_i_adra_d,
      da_d => vec_rsc_0_8_i_da_d,
      qa_d => vec_rsc_0_8_i_qa_d_1,
      wea_d => vec_rsc_0_8_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_0_8_i_wea_d_iff
    );
  vec_rsc_0_8_i_qa <= vec_rsc_0_8_qa;
  vec_rsc_0_8_da <= vec_rsc_0_8_i_da;
  vec_rsc_0_8_adra <= vec_rsc_0_8_i_adra;
  vec_rsc_0_8_i_adra_d <= vec_rsc_0_0_i_adra_d_iff;
  vec_rsc_0_8_i_da_d <= vec_rsc_0_0_i_da_d_iff;
  vec_rsc_0_8_i_qa_d <= vec_rsc_0_8_i_qa_d_1;

  vec_rsc_0_9_i : inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_13_8_64_256_256_64_1_gen
    PORT MAP(
      qa => vec_rsc_0_9_i_qa,
      wea => vec_rsc_0_9_wea,
      da => vec_rsc_0_9_i_da,
      adra => vec_rsc_0_9_i_adra,
      adra_d => vec_rsc_0_9_i_adra_d,
      da_d => vec_rsc_0_9_i_da_d,
      qa_d => vec_rsc_0_9_i_qa_d_1,
      wea_d => vec_rsc_0_9_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_0_9_i_wea_d_iff
    );
  vec_rsc_0_9_i_qa <= vec_rsc_0_9_qa;
  vec_rsc_0_9_da <= vec_rsc_0_9_i_da;
  vec_rsc_0_9_adra <= vec_rsc_0_9_i_adra;
  vec_rsc_0_9_i_adra_d <= vec_rsc_0_0_i_adra_d_iff;
  vec_rsc_0_9_i_da_d <= vec_rsc_0_0_i_da_d_iff;
  vec_rsc_0_9_i_qa_d <= vec_rsc_0_9_i_qa_d_1;

  vec_rsc_0_10_i : inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_14_8_64_256_256_64_1_gen
    PORT MAP(
      qa => vec_rsc_0_10_i_qa,
      wea => vec_rsc_0_10_wea,
      da => vec_rsc_0_10_i_da,
      adra => vec_rsc_0_10_i_adra,
      adra_d => vec_rsc_0_10_i_adra_d,
      da_d => vec_rsc_0_10_i_da_d,
      qa_d => vec_rsc_0_10_i_qa_d_1,
      wea_d => vec_rsc_0_10_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_0_10_i_wea_d_iff
    );
  vec_rsc_0_10_i_qa <= vec_rsc_0_10_qa;
  vec_rsc_0_10_da <= vec_rsc_0_10_i_da;
  vec_rsc_0_10_adra <= vec_rsc_0_10_i_adra;
  vec_rsc_0_10_i_adra_d <= vec_rsc_0_0_i_adra_d_iff;
  vec_rsc_0_10_i_da_d <= vec_rsc_0_0_i_da_d_iff;
  vec_rsc_0_10_i_qa_d <= vec_rsc_0_10_i_qa_d_1;

  vec_rsc_0_11_i : inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_15_8_64_256_256_64_1_gen
    PORT MAP(
      qa => vec_rsc_0_11_i_qa,
      wea => vec_rsc_0_11_wea,
      da => vec_rsc_0_11_i_da,
      adra => vec_rsc_0_11_i_adra,
      adra_d => vec_rsc_0_11_i_adra_d,
      da_d => vec_rsc_0_11_i_da_d,
      qa_d => vec_rsc_0_11_i_qa_d_1,
      wea_d => vec_rsc_0_11_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_0_11_i_wea_d_iff
    );
  vec_rsc_0_11_i_qa <= vec_rsc_0_11_qa;
  vec_rsc_0_11_da <= vec_rsc_0_11_i_da;
  vec_rsc_0_11_adra <= vec_rsc_0_11_i_adra;
  vec_rsc_0_11_i_adra_d <= vec_rsc_0_0_i_adra_d_iff;
  vec_rsc_0_11_i_da_d <= vec_rsc_0_0_i_da_d_iff;
  vec_rsc_0_11_i_qa_d <= vec_rsc_0_11_i_qa_d_1;

  vec_rsc_0_12_i : inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_16_8_64_256_256_64_1_gen
    PORT MAP(
      qa => vec_rsc_0_12_i_qa,
      wea => vec_rsc_0_12_wea,
      da => vec_rsc_0_12_i_da,
      adra => vec_rsc_0_12_i_adra,
      adra_d => vec_rsc_0_12_i_adra_d,
      da_d => vec_rsc_0_12_i_da_d,
      qa_d => vec_rsc_0_12_i_qa_d_1,
      wea_d => vec_rsc_0_12_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_0_12_i_wea_d_iff
    );
  vec_rsc_0_12_i_qa <= vec_rsc_0_12_qa;
  vec_rsc_0_12_da <= vec_rsc_0_12_i_da;
  vec_rsc_0_12_adra <= vec_rsc_0_12_i_adra;
  vec_rsc_0_12_i_adra_d <= vec_rsc_0_0_i_adra_d_iff;
  vec_rsc_0_12_i_da_d <= vec_rsc_0_0_i_da_d_iff;
  vec_rsc_0_12_i_qa_d <= vec_rsc_0_12_i_qa_d_1;

  vec_rsc_0_13_i : inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_17_8_64_256_256_64_1_gen
    PORT MAP(
      qa => vec_rsc_0_13_i_qa,
      wea => vec_rsc_0_13_wea,
      da => vec_rsc_0_13_i_da,
      adra => vec_rsc_0_13_i_adra,
      adra_d => vec_rsc_0_13_i_adra_d,
      da_d => vec_rsc_0_13_i_da_d,
      qa_d => vec_rsc_0_13_i_qa_d_1,
      wea_d => vec_rsc_0_13_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_0_13_i_wea_d_iff
    );
  vec_rsc_0_13_i_qa <= vec_rsc_0_13_qa;
  vec_rsc_0_13_da <= vec_rsc_0_13_i_da;
  vec_rsc_0_13_adra <= vec_rsc_0_13_i_adra;
  vec_rsc_0_13_i_adra_d <= vec_rsc_0_0_i_adra_d_iff;
  vec_rsc_0_13_i_da_d <= vec_rsc_0_0_i_da_d_iff;
  vec_rsc_0_13_i_qa_d <= vec_rsc_0_13_i_qa_d_1;

  vec_rsc_0_14_i : inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_18_8_64_256_256_64_1_gen
    PORT MAP(
      qa => vec_rsc_0_14_i_qa,
      wea => vec_rsc_0_14_wea,
      da => vec_rsc_0_14_i_da,
      adra => vec_rsc_0_14_i_adra,
      adra_d => vec_rsc_0_14_i_adra_d,
      da_d => vec_rsc_0_14_i_da_d,
      qa_d => vec_rsc_0_14_i_qa_d_1,
      wea_d => vec_rsc_0_14_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_0_14_i_wea_d_iff
    );
  vec_rsc_0_14_i_qa <= vec_rsc_0_14_qa;
  vec_rsc_0_14_da <= vec_rsc_0_14_i_da;
  vec_rsc_0_14_adra <= vec_rsc_0_14_i_adra;
  vec_rsc_0_14_i_adra_d <= vec_rsc_0_0_i_adra_d_iff;
  vec_rsc_0_14_i_da_d <= vec_rsc_0_0_i_da_d_iff;
  vec_rsc_0_14_i_qa_d <= vec_rsc_0_14_i_qa_d_1;

  vec_rsc_0_15_i : inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_19_8_64_256_256_64_1_gen
    PORT MAP(
      qa => vec_rsc_0_15_i_qa,
      wea => vec_rsc_0_15_wea,
      da => vec_rsc_0_15_i_da,
      adra => vec_rsc_0_15_i_adra,
      adra_d => vec_rsc_0_15_i_adra_d,
      da_d => vec_rsc_0_15_i_da_d,
      qa_d => vec_rsc_0_15_i_qa_d_1,
      wea_d => vec_rsc_0_15_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_0_15_i_wea_d_iff
    );
  vec_rsc_0_15_i_qa <= vec_rsc_0_15_qa;
  vec_rsc_0_15_da <= vec_rsc_0_15_i_da;
  vec_rsc_0_15_adra <= vec_rsc_0_15_i_adra;
  vec_rsc_0_15_i_adra_d <= vec_rsc_0_0_i_adra_d_iff;
  vec_rsc_0_15_i_da_d <= vec_rsc_0_0_i_da_d_iff;
  vec_rsc_0_15_i_qa_d <= vec_rsc_0_15_i_qa_d_1;

  inPlaceNTT_DIT_core_inst : inPlaceNTT_DIT_core
    PORT MAP(
      clk => clk,
      rst => rst,
      vec_rsc_triosy_0_0_lz => vec_rsc_triosy_0_0_lz,
      vec_rsc_triosy_0_1_lz => vec_rsc_triosy_0_1_lz,
      vec_rsc_triosy_0_2_lz => vec_rsc_triosy_0_2_lz,
      vec_rsc_triosy_0_3_lz => vec_rsc_triosy_0_3_lz,
      vec_rsc_triosy_0_4_lz => vec_rsc_triosy_0_4_lz,
      vec_rsc_triosy_0_5_lz => vec_rsc_triosy_0_5_lz,
      vec_rsc_triosy_0_6_lz => vec_rsc_triosy_0_6_lz,
      vec_rsc_triosy_0_7_lz => vec_rsc_triosy_0_7_lz,
      vec_rsc_triosy_0_8_lz => vec_rsc_triosy_0_8_lz,
      vec_rsc_triosy_0_9_lz => vec_rsc_triosy_0_9_lz,
      vec_rsc_triosy_0_10_lz => vec_rsc_triosy_0_10_lz,
      vec_rsc_triosy_0_11_lz => vec_rsc_triosy_0_11_lz,
      vec_rsc_triosy_0_12_lz => vec_rsc_triosy_0_12_lz,
      vec_rsc_triosy_0_13_lz => vec_rsc_triosy_0_13_lz,
      vec_rsc_triosy_0_14_lz => vec_rsc_triosy_0_14_lz,
      vec_rsc_triosy_0_15_lz => vec_rsc_triosy_0_15_lz,
      p_rsc_dat => inPlaceNTT_DIT_core_inst_p_rsc_dat,
      p_rsc_triosy_lz => p_rsc_triosy_lz,
      r_rsc_dat => inPlaceNTT_DIT_core_inst_r_rsc_dat,
      r_rsc_triosy_lz => r_rsc_triosy_lz,
      vec_rsc_0_0_i_qa_d => inPlaceNTT_DIT_core_inst_vec_rsc_0_0_i_qa_d,
      vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_1_i_qa_d => inPlaceNTT_DIT_core_inst_vec_rsc_0_1_i_qa_d,
      vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_2_i_qa_d => inPlaceNTT_DIT_core_inst_vec_rsc_0_2_i_qa_d,
      vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_3_i_qa_d => inPlaceNTT_DIT_core_inst_vec_rsc_0_3_i_qa_d,
      vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_4_i_qa_d => inPlaceNTT_DIT_core_inst_vec_rsc_0_4_i_qa_d,
      vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_5_i_qa_d => inPlaceNTT_DIT_core_inst_vec_rsc_0_5_i_qa_d,
      vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_6_i_qa_d => inPlaceNTT_DIT_core_inst_vec_rsc_0_6_i_qa_d,
      vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_7_i_qa_d => inPlaceNTT_DIT_core_inst_vec_rsc_0_7_i_qa_d,
      vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_8_i_qa_d => inPlaceNTT_DIT_core_inst_vec_rsc_0_8_i_qa_d,
      vec_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_9_i_qa_d => inPlaceNTT_DIT_core_inst_vec_rsc_0_9_i_qa_d,
      vec_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_10_i_qa_d => inPlaceNTT_DIT_core_inst_vec_rsc_0_10_i_qa_d,
      vec_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_11_i_qa_d => inPlaceNTT_DIT_core_inst_vec_rsc_0_11_i_qa_d,
      vec_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_12_i_qa_d => inPlaceNTT_DIT_core_inst_vec_rsc_0_12_i_qa_d,
      vec_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_13_i_qa_d => inPlaceNTT_DIT_core_inst_vec_rsc_0_13_i_qa_d,
      vec_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_14_i_qa_d => inPlaceNTT_DIT_core_inst_vec_rsc_0_14_i_qa_d,
      vec_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_15_i_qa_d => inPlaceNTT_DIT_core_inst_vec_rsc_0_15_i_qa_d,
      vec_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_0_i_adra_d_pff => inPlaceNTT_DIT_core_inst_vec_rsc_0_0_i_adra_d_pff,
      vec_rsc_0_0_i_da_d_pff => inPlaceNTT_DIT_core_inst_vec_rsc_0_0_i_da_d_pff,
      vec_rsc_0_0_i_wea_d_pff => vec_rsc_0_0_i_wea_d_iff,
      vec_rsc_0_1_i_wea_d_pff => vec_rsc_0_1_i_wea_d_iff,
      vec_rsc_0_2_i_wea_d_pff => vec_rsc_0_2_i_wea_d_iff,
      vec_rsc_0_3_i_wea_d_pff => vec_rsc_0_3_i_wea_d_iff,
      vec_rsc_0_4_i_wea_d_pff => vec_rsc_0_4_i_wea_d_iff,
      vec_rsc_0_5_i_wea_d_pff => vec_rsc_0_5_i_wea_d_iff,
      vec_rsc_0_6_i_wea_d_pff => vec_rsc_0_6_i_wea_d_iff,
      vec_rsc_0_7_i_wea_d_pff => vec_rsc_0_7_i_wea_d_iff,
      vec_rsc_0_8_i_wea_d_pff => vec_rsc_0_8_i_wea_d_iff,
      vec_rsc_0_9_i_wea_d_pff => vec_rsc_0_9_i_wea_d_iff,
      vec_rsc_0_10_i_wea_d_pff => vec_rsc_0_10_i_wea_d_iff,
      vec_rsc_0_11_i_wea_d_pff => vec_rsc_0_11_i_wea_d_iff,
      vec_rsc_0_12_i_wea_d_pff => vec_rsc_0_12_i_wea_d_iff,
      vec_rsc_0_13_i_wea_d_pff => vec_rsc_0_13_i_wea_d_iff,
      vec_rsc_0_14_i_wea_d_pff => vec_rsc_0_14_i_wea_d_iff,
      vec_rsc_0_15_i_wea_d_pff => vec_rsc_0_15_i_wea_d_iff
    );
  inPlaceNTT_DIT_core_inst_p_rsc_dat <= p_rsc_dat;
  inPlaceNTT_DIT_core_inst_r_rsc_dat <= r_rsc_dat;
  inPlaceNTT_DIT_core_inst_vec_rsc_0_0_i_qa_d <= vec_rsc_0_0_i_qa_d;
  inPlaceNTT_DIT_core_inst_vec_rsc_0_1_i_qa_d <= vec_rsc_0_1_i_qa_d;
  inPlaceNTT_DIT_core_inst_vec_rsc_0_2_i_qa_d <= vec_rsc_0_2_i_qa_d;
  inPlaceNTT_DIT_core_inst_vec_rsc_0_3_i_qa_d <= vec_rsc_0_3_i_qa_d;
  inPlaceNTT_DIT_core_inst_vec_rsc_0_4_i_qa_d <= vec_rsc_0_4_i_qa_d;
  inPlaceNTT_DIT_core_inst_vec_rsc_0_5_i_qa_d <= vec_rsc_0_5_i_qa_d;
  inPlaceNTT_DIT_core_inst_vec_rsc_0_6_i_qa_d <= vec_rsc_0_6_i_qa_d;
  inPlaceNTT_DIT_core_inst_vec_rsc_0_7_i_qa_d <= vec_rsc_0_7_i_qa_d;
  inPlaceNTT_DIT_core_inst_vec_rsc_0_8_i_qa_d <= vec_rsc_0_8_i_qa_d;
  inPlaceNTT_DIT_core_inst_vec_rsc_0_9_i_qa_d <= vec_rsc_0_9_i_qa_d;
  inPlaceNTT_DIT_core_inst_vec_rsc_0_10_i_qa_d <= vec_rsc_0_10_i_qa_d;
  inPlaceNTT_DIT_core_inst_vec_rsc_0_11_i_qa_d <= vec_rsc_0_11_i_qa_d;
  inPlaceNTT_DIT_core_inst_vec_rsc_0_12_i_qa_d <= vec_rsc_0_12_i_qa_d;
  inPlaceNTT_DIT_core_inst_vec_rsc_0_13_i_qa_d <= vec_rsc_0_13_i_qa_d;
  inPlaceNTT_DIT_core_inst_vec_rsc_0_14_i_qa_d <= vec_rsc_0_14_i_qa_d;
  inPlaceNTT_DIT_core_inst_vec_rsc_0_15_i_qa_d <= vec_rsc_0_15_i_qa_d;
  vec_rsc_0_0_i_adra_d_iff <= inPlaceNTT_DIT_core_inst_vec_rsc_0_0_i_adra_d_pff;
  vec_rsc_0_0_i_da_d_iff <= inPlaceNTT_DIT_core_inst_vec_rsc_0_0_i_da_d_pff;

END v44;



