
//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_io_sync_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_io_sync_v2 (ld, lz);
    parameter valid = 0;

    input  ld;
    output lz;

    wire   lz;

    assign lz = ld;

endmodule


//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_out_dreg_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_out_dreg_v2 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input    [width-1:0] d;
  output   [width-1:0] z;

  wire     [width-1:0] z;

  assign z = d;

endmodule

//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_rem_beh.v 
module mgc_rem(a,b,z);
   parameter width_a = 8;
   parameter width_b = 8;
   parameter signd = 1;
   input [width_a-1:0] a;
   input [width_b-1:0] b; 
   output [width_b-1:0] z;  
   reg  [width_b-1:0] z;

   always@(a or b)
     begin
	if(signd)
	  rem_s(a,b,z);
	else
          rem_u(a,b,z);
     end


//-----------------------------------------------------------------
//     -- Vectorized Overloaded Arithmetic Operators
//-----------------------------------------------------------------
   
   function [width_a-1:0] fabs_l; 
      input [width_a-1:0] arg1;
      begin
         case(arg1[width_a-1])
            1'b1:
               fabs_l = {(width_a){1'b0}} - arg1;
            default: // was: 1'b0:
               fabs_l = arg1;
         endcase
      end
   endfunction
   
   function [width_b-1:0] fabs_r; 
      input [width_b-1:0] arg1;
      begin
         case (arg1[width_b-1])
            1'b1:
               fabs_r =  {(width_b){1'b0}} - arg1;
            default: // was: 1'b0:
               fabs_r = arg1;
         endcase
      end
   endfunction

   function [width_b:0] minus;
     input [width_b:0] in1;
     input [width_b:0] in2;
     reg [width_b+1:0] tmp;
     begin
       tmp = in1 - in2;
       minus = tmp[width_b:0];
     end
   endfunction

   
   task divmod;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      output [width_b-1:0] rmod;
      
      parameter llen = width_a;
      parameter rlen = width_b;
      reg [(llen+rlen)-1:0] lbuf;
      reg [rlen:0] diff;
	  integer i;
      begin
	 lbuf = {(llen+rlen){1'b0}};
//64'b0;
	 lbuf[llen-1:0] = l;
	 for(i=width_a-1;i>=0;i=i-1)
	   begin
              diff = minus(lbuf[(llen+rlen)-1:llen-1], {1'b0,r});
	      rdiv[i] = ~diff[rlen];
	      if(diff[rlen] == 0)
		lbuf[(llen+rlen)-1:llen-1] = diff;
	      lbuf[(llen+rlen)-1:1] = lbuf[(llen+rlen)-2:0];
	   end
	 rmod = lbuf[(llen+rlen)-1:llen];
      end
   endtask
      

   task div_u;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(l, r, rdiv, rmod);
      end
   endtask
   
   task mod_u;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_b-1:0] rmod;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(l, r, rdiv, rmod);
      end
   endtask

   task rem_u; 
      input [width_a-1:0] l;
      input [width_b-1:0] r;    
      output [width_b-1:0] rmod;
      begin
	 mod_u(l,r,rmod);
      end
   endtask // rem_u

   task div_s;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(fabs_l(l), fabs_r(r),rdiv,rmod);
	 if(l[width_a-1] != r[width_b-1])
	   rdiv = {(width_a){1'b0}} - rdiv;
      end
   endtask

   task mod_s;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_b-1:0] rmod;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      reg [width_b-1:0] rnul;
      reg [width_b:0] rmod_t;
      begin
         rnul = {width_b{1'b0}};
	 divmod(fabs_l(l), fabs_r(r), rdiv, rmod);
         if (l[width_a-1])
	   rmod = {(width_b){1'b0}} - rmod;
	 if((rmod != rnul) && (l[width_a-1] != r[width_b-1]))
            begin
               rmod_t = r + rmod;
               rmod = rmod_t[width_b-1:0];
            end
      end
   endtask // mod_s
   
   task rem_s; 
      input [width_a-1:0] l;
      input [width_b-1:0] r;    
      output [width_b-1:0] rmod;   
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(fabs_l(l),fabs_r(r),rdiv,rmod);
	 if(l[width_a-1])
	   rmod = {(width_b){1'b0}} - rmod;
      end
   endtask

  endmodule

//------> ../td_ccore_solutions/modulo_dev_bb61c76201db0c9669a47462bb7d006361ff_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5c/896140 Production Release
//  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
// 
//  Generated by:   yl7897@newnano.poly.edu
//  Generated date: Tue Jul 20 15:24:30 2021
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    modulo_dev_core
// ------------------------------------------------------------------


module modulo_dev_core (
  base_rsc_dat, m_rsc_dat, return_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk,
      ccs_ccore_srst, ccs_ccore_en
);
  input [63:0] base_rsc_dat;
  input [63:0] m_rsc_dat;
  output [63:0] return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_srst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [63:0] base_rsci_idat;
  wire [63:0] m_rsci_idat;
  reg [63:0] return_rsci_d;
  wire ccs_ccore_start_rsci_idat;
  wire [64:0] rem_13_cmp_z;
  wire [64:0] rem_13_cmp_1_z;
  wire [64:0] rem_13_cmp_2_z;
  wire [64:0] rem_13_cmp_3_z;
  wire [64:0] rem_13_cmp_4_z;
  wire [64:0] rem_13_cmp_5_z;
  wire [64:0] rem_13_cmp_6_z;
  wire [64:0] rem_13_cmp_7_z;
  wire [64:0] rem_13_cmp_8_z;
  wire [64:0] rem_13_cmp_9_z;
  wire [64:0] rem_13_cmp_10_z;
  wire [64:0] rem_13_cmp_11_z;
  reg [63:0] rem_13_cmp_b_63_0;
  reg [63:0] rem_13_cmp_1_b_63_0;
  reg [63:0] rem_13_cmp_2_b_63_0;
  reg [63:0] rem_13_cmp_3_b_63_0;
  reg [63:0] rem_13_cmp_4_b_63_0;
  reg [63:0] rem_13_cmp_5_b_63_0;
  reg [63:0] rem_13_cmp_6_b_63_0;
  reg [63:0] rem_13_cmp_7_b_63_0;
  reg [63:0] rem_13_cmp_8_b_63_0;
  reg [63:0] rem_13_cmp_9_b_63_0;
  reg [63:0] rem_13_cmp_10_b_63_0;
  reg [63:0] rem_13_cmp_11_b_63_0;
  reg [63:0] rem_13_cmp_a_63_0;
  reg [63:0] rem_13_cmp_1_a_63_0;
  reg [63:0] rem_13_cmp_2_a_63_0;
  reg [63:0] rem_13_cmp_3_a_63_0;
  reg [63:0] rem_13_cmp_4_a_63_0;
  reg [63:0] rem_13_cmp_5_a_63_0;
  reg [63:0] rem_13_cmp_6_a_63_0;
  reg [63:0] rem_13_cmp_7_a_63_0;
  reg [63:0] rem_13_cmp_8_a_63_0;
  reg [63:0] rem_13_cmp_9_a_63_0;
  reg [63:0] rem_13_cmp_10_a_63_0;
  reg [63:0] rem_13_cmp_11_a_63_0;
  wire [1:0] acc_tmp;
  wire [2:0] nl_acc_tmp;
  wire [3:0] acc_1_tmp;
  wire [4:0] nl_acc_1_tmp;
  wire and_dcpl_1;
  wire and_dcpl_2;
  wire and_dcpl_3;
  wire and_dcpl_4;
  wire and_dcpl_6;
  wire and_dcpl_8;
  wire and_dcpl_9;
  wire and_dcpl_11;
  wire and_dcpl_13;
  wire and_dcpl_18;
  wire and_dcpl_23;
  wire and_dcpl_28;
  wire and_dcpl_29;
  wire and_dcpl_30;
  wire and_dcpl_31;
  wire and_dcpl_33;
  wire and_dcpl_35;
  wire and_dcpl_36;
  wire and_dcpl_38;
  wire and_dcpl_40;
  wire and_dcpl_45;
  wire and_dcpl_50;
  wire and_dcpl_55;
  wire and_dcpl_56;
  wire and_dcpl_57;
  wire and_dcpl_58;
  wire and_dcpl_60;
  wire and_dcpl_62;
  wire and_dcpl_63;
  wire and_dcpl_65;
  wire and_dcpl_67;
  wire and_dcpl_72;
  wire and_dcpl_77;
  wire and_dcpl_82;
  wire and_dcpl_83;
  wire and_dcpl_84;
  wire and_dcpl_85;
  wire and_dcpl_87;
  wire and_dcpl_89;
  wire and_dcpl_90;
  wire and_dcpl_92;
  wire and_dcpl_94;
  wire and_dcpl_99;
  wire and_dcpl_104;
  wire and_dcpl_109;
  wire and_dcpl_110;
  wire and_dcpl_111;
  wire and_dcpl_112;
  wire and_dcpl_114;
  wire and_dcpl_115;
  wire and_dcpl_117;
  wire and_dcpl_119;
  wire and_dcpl_121;
  wire and_dcpl_126;
  wire and_dcpl_129;
  wire and_dcpl_136;
  wire and_dcpl_137;
  wire and_dcpl_138;
  wire and_dcpl_139;
  wire and_dcpl_141;
  wire and_dcpl_143;
  wire and_dcpl_144;
  wire and_dcpl_146;
  wire and_dcpl_148;
  wire and_dcpl_153;
  wire and_dcpl_158;
  wire and_dcpl_163;
  wire and_dcpl_164;
  wire and_dcpl_165;
  wire and_dcpl_166;
  wire and_dcpl_168;
  wire and_dcpl_170;
  wire and_dcpl_171;
  wire and_dcpl_173;
  wire and_dcpl_175;
  wire and_dcpl_180;
  wire and_dcpl_185;
  wire and_dcpl_190;
  wire and_dcpl_191;
  wire and_dcpl_192;
  wire and_dcpl_193;
  wire and_dcpl_195;
  wire and_dcpl_197;
  wire and_dcpl_198;
  wire and_dcpl_200;
  wire and_dcpl_202;
  wire and_dcpl_207;
  wire and_dcpl_212;
  wire and_dcpl_217;
  wire and_dcpl_218;
  wire and_dcpl_219;
  wire and_dcpl_220;
  wire and_dcpl_222;
  wire and_dcpl_224;
  wire and_dcpl_225;
  wire and_dcpl_227;
  wire and_dcpl_229;
  wire and_dcpl_234;
  wire and_dcpl_239;
  wire and_dcpl_244;
  wire and_dcpl_245;
  wire and_dcpl_246;
  wire and_dcpl_247;
  wire and_dcpl_249;
  wire and_dcpl_251;
  wire and_dcpl_252;
  wire and_dcpl_254;
  wire and_dcpl_256;
  wire and_dcpl_261;
  wire and_dcpl_266;
  wire and_dcpl_271;
  wire and_dcpl_272;
  wire and_dcpl_274;
  wire and_dcpl_276;
  wire and_dcpl_278;
  wire and_dcpl_280;
  wire and_dcpl_285;
  wire and_dcpl_291;
  wire and_dcpl_292;
  wire and_dcpl_293;
  wire and_dcpl_294;
  wire and_dcpl_295;
  wire and_dcpl_296;
  wire and_dcpl_298;
  wire not_tmp_54;
  wire or_tmp_2;
  wire and_dcpl_300;
  wire and_dcpl_301;
  wire and_dcpl_302;
  wire and_dcpl_304;
  wire and_tmp;
  wire and_dcpl_306;
  wire and_dcpl_307;
  wire and_dcpl_308;
  wire and_dcpl_310;
  wire and_tmp_2;
  wire and_dcpl_312;
  wire and_dcpl_313;
  wire and_dcpl_314;
  wire and_dcpl_316;
  wire and_tmp_5;
  wire and_dcpl_318;
  wire and_tmp_9;
  wire and_dcpl_324;
  wire and_tmp_13;
  wire and_dcpl_330;
  wire mux_tmp_19;
  wire and_tmp_17;
  wire and_dcpl_336;
  wire mux_tmp_22;
  wire mux_tmp_23;
  wire and_tmp_21;
  wire and_dcpl_342;
  wire mux_tmp_26;
  wire mux_tmp_27;
  wire mux_tmp_28;
  wire and_tmp_25;
  wire and_dcpl_348;
  wire and_tmp_35;
  wire and_dcpl_355;
  wire and_dcpl_356;
  wire and_dcpl_358;
  wire or_tmp_80;
  wire and_dcpl_360;
  wire and_dcpl_362;
  wire mux_tmp_32;
  wire and_dcpl_364;
  wire and_dcpl_366;
  wire mux_tmp_34;
  wire mux_tmp_35;
  wire and_dcpl_368;
  wire and_dcpl_370;
  wire mux_tmp_37;
  wire mux_tmp_38;
  wire mux_tmp_39;
  wire and_dcpl_372;
  wire mux_tmp_41;
  wire mux_tmp_42;
  wire mux_tmp_43;
  wire mux_tmp_44;
  wire and_dcpl_376;
  wire mux_tmp_46;
  wire mux_tmp_47;
  wire mux_tmp_48;
  wire mux_tmp_49;
  wire mux_tmp_50;
  wire and_dcpl_379;
  wire mux_tmp_52;
  wire mux_tmp_53;
  wire mux_tmp_54;
  wire mux_tmp_55;
  wire mux_tmp_56;
  wire mux_tmp_57;
  wire and_dcpl_382;
  wire mux_tmp_59;
  wire mux_tmp_60;
  wire mux_tmp_61;
  wire mux_tmp_62;
  wire mux_tmp_63;
  wire mux_tmp_64;
  wire mux_tmp_65;
  wire and_dcpl_385;
  wire mux_tmp_67;
  wire mux_tmp_68;
  wire mux_tmp_69;
  wire mux_tmp_70;
  wire mux_tmp_71;
  wire mux_tmp_72;
  wire mux_tmp_73;
  wire mux_tmp_74;
  wire and_dcpl_388;
  wire and_tmp_44;
  wire mux_tmp_76;
  wire and_dcpl_393;
  wire and_dcpl_394;
  wire and_dcpl_395;
  wire or_tmp_185;
  wire and_dcpl_397;
  wire and_dcpl_398;
  wire and_tmp_45;
  wire and_dcpl_400;
  wire and_dcpl_401;
  wire and_tmp_47;
  wire and_dcpl_403;
  wire and_dcpl_404;
  wire and_tmp_50;
  wire and_dcpl_406;
  wire and_tmp_54;
  wire and_dcpl_409;
  wire and_tmp_58;
  wire and_dcpl_413;
  wire mux_tmp_84;
  wire and_tmp_62;
  wire and_dcpl_417;
  wire mux_tmp_87;
  wire mux_tmp_88;
  wire and_tmp_66;
  wire and_dcpl_421;
  wire mux_tmp_91;
  wire mux_tmp_92;
  wire mux_tmp_93;
  wire and_tmp_70;
  wire and_dcpl_425;
  wire and_tmp_80;
  wire and_dcpl_430;
  wire and_dcpl_431;
  wire or_tmp_263;
  wire and_dcpl_433;
  wire mux_tmp_97;
  wire and_dcpl_435;
  wire mux_tmp_99;
  wire mux_tmp_100;
  wire and_dcpl_437;
  wire mux_tmp_102;
  wire mux_tmp_103;
  wire mux_tmp_104;
  wire and_dcpl_439;
  wire mux_tmp_106;
  wire mux_tmp_107;
  wire mux_tmp_108;
  wire mux_tmp_109;
  wire and_dcpl_442;
  wire mux_tmp_111;
  wire mux_tmp_112;
  wire mux_tmp_113;
  wire mux_tmp_114;
  wire mux_tmp_115;
  wire and_dcpl_445;
  wire mux_tmp_117;
  wire mux_tmp_118;
  wire mux_tmp_119;
  wire mux_tmp_120;
  wire mux_tmp_121;
  wire mux_tmp_122;
  wire and_dcpl_448;
  wire mux_tmp_124;
  wire mux_tmp_125;
  wire mux_tmp_126;
  wire mux_tmp_127;
  wire mux_tmp_128;
  wire mux_tmp_129;
  wire mux_tmp_130;
  wire and_dcpl_451;
  wire mux_tmp_132;
  wire mux_tmp_133;
  wire mux_tmp_134;
  wire mux_tmp_135;
  wire mux_tmp_136;
  wire mux_tmp_137;
  wire mux_tmp_138;
  wire mux_tmp_139;
  wire and_dcpl_454;
  wire and_tmp_89;
  wire mux_tmp_141;
  wire and_dcpl_460;
  wire and_dcpl_461;
  wire and_dcpl_462;
  wire and_dcpl_463;
  wire not_tmp_332;
  wire or_tmp_368;
  wire and_dcpl_465;
  wire and_dcpl_466;
  wire and_dcpl_467;
  wire and_tmp_90;
  wire and_dcpl_469;
  wire and_dcpl_470;
  wire and_dcpl_471;
  wire and_tmp_92;
  wire and_dcpl_473;
  wire and_dcpl_474;
  wire and_dcpl_475;
  wire and_tmp_95;
  wire and_dcpl_477;
  wire and_tmp_99;
  wire and_dcpl_480;
  wire and_tmp_103;
  wire and_dcpl_483;
  wire mux_tmp_149;
  wire and_tmp_107;
  wire and_dcpl_486;
  wire mux_tmp_152;
  wire mux_tmp_153;
  wire and_tmp_111;
  wire and_dcpl_489;
  wire mux_tmp_156;
  wire mux_tmp_157;
  wire mux_tmp_158;
  wire and_tmp_115;
  wire and_dcpl_492;
  wire and_tmp_125;
  wire and_dcpl_498;
  wire or_tmp_446;
  wire and_dcpl_500;
  wire mux_tmp_162;
  wire and_dcpl_502;
  wire mux_tmp_164;
  wire mux_tmp_165;
  wire and_dcpl_504;
  wire mux_tmp_167;
  wire mux_tmp_168;
  wire mux_tmp_169;
  wire and_dcpl_506;
  wire mux_tmp_171;
  wire mux_tmp_172;
  wire mux_tmp_173;
  wire mux_tmp_174;
  wire and_dcpl_508;
  wire mux_tmp_176;
  wire mux_tmp_177;
  wire mux_tmp_178;
  wire mux_tmp_179;
  wire mux_tmp_180;
  wire and_dcpl_510;
  wire mux_tmp_182;
  wire mux_tmp_183;
  wire mux_tmp_184;
  wire mux_tmp_185;
  wire mux_tmp_186;
  wire mux_tmp_187;
  wire and_dcpl_512;
  wire mux_tmp_189;
  wire mux_tmp_190;
  wire mux_tmp_191;
  wire mux_tmp_192;
  wire mux_tmp_193;
  wire mux_tmp_194;
  wire mux_tmp_195;
  wire and_dcpl_514;
  wire mux_tmp_197;
  wire mux_tmp_198;
  wire mux_tmp_199;
  wire mux_tmp_200;
  wire mux_tmp_201;
  wire mux_tmp_202;
  wire mux_tmp_203;
  wire mux_tmp_204;
  wire and_dcpl_516;
  wire and_tmp_134;
  wire mux_tmp_206;
  wire and_dcpl_520;
  wire and_dcpl_521;
  wire or_tmp_551;
  wire and_dcpl_523;
  wire and_dcpl_524;
  wire and_tmp_135;
  wire and_dcpl_526;
  wire and_dcpl_527;
  wire and_tmp_137;
  wire and_dcpl_529;
  wire and_dcpl_530;
  wire and_tmp_140;
  wire and_dcpl_532;
  wire and_tmp_144;
  wire and_dcpl_534;
  wire and_tmp_148;
  wire and_dcpl_536;
  wire mux_tmp_214;
  wire and_tmp_152;
  wire and_dcpl_538;
  wire mux_tmp_217;
  wire mux_tmp_218;
  wire and_tmp_156;
  wire and_dcpl_540;
  wire mux_tmp_221;
  wire mux_tmp_222;
  wire mux_tmp_223;
  wire and_tmp_160;
  wire and_dcpl_542;
  wire and_tmp_170;
  wire and_dcpl_546;
  wire or_tmp_629;
  wire and_dcpl_548;
  wire mux_tmp_227;
  wire and_dcpl_550;
  wire mux_tmp_229;
  wire mux_tmp_230;
  wire and_dcpl_552;
  wire mux_tmp_232;
  wire mux_tmp_233;
  wire mux_tmp_234;
  wire and_dcpl_554;
  wire mux_tmp_236;
  wire mux_tmp_237;
  wire mux_tmp_238;
  wire mux_tmp_239;
  wire and_dcpl_556;
  wire mux_tmp_241;
  wire mux_tmp_242;
  wire mux_tmp_243;
  wire mux_tmp_244;
  wire mux_tmp_245;
  wire and_dcpl_558;
  wire mux_tmp_247;
  wire mux_tmp_248;
  wire mux_tmp_249;
  wire mux_tmp_250;
  wire mux_tmp_251;
  wire mux_tmp_252;
  wire and_dcpl_560;
  wire mux_tmp_254;
  wire mux_tmp_255;
  wire mux_tmp_256;
  wire mux_tmp_257;
  wire mux_tmp_258;
  wire mux_tmp_259;
  wire mux_tmp_260;
  wire and_dcpl_562;
  wire mux_tmp_262;
  wire mux_tmp_263;
  wire mux_tmp_264;
  wire mux_tmp_265;
  wire mux_tmp_266;
  wire mux_tmp_267;
  wire mux_tmp_268;
  wire mux_tmp_269;
  wire and_dcpl_564;
  wire and_tmp_179;
  wire mux_tmp_271;
  wire and_dcpl_568;
  wire and_dcpl_569;
  wire and_dcpl_570;
  wire and_dcpl_571;
  wire or_tmp_733;
  wire and_dcpl_573;
  wire and_dcpl_574;
  wire and_dcpl_575;
  wire and_tmp_180;
  wire and_dcpl_577;
  wire and_dcpl_578;
  wire and_dcpl_579;
  wire and_tmp_182;
  wire and_dcpl_581;
  wire and_dcpl_582;
  wire and_dcpl_583;
  wire and_tmp_185;
  wire and_dcpl_585;
  wire and_tmp_189;
  wire and_dcpl_589;
  wire and_tmp_193;
  wire and_dcpl_593;
  wire mux_tmp_279;
  wire and_tmp_197;
  wire and_dcpl_597;
  wire mux_tmp_282;
  wire mux_tmp_283;
  wire and_tmp_201;
  wire and_dcpl_601;
  wire mux_tmp_286;
  wire mux_tmp_287;
  wire mux_tmp_288;
  wire and_tmp_205;
  wire and_dcpl_605;
  wire or_tmp_808;
  wire mux_tmp_291;
  wire mux_tmp_292;
  wire mux_tmp_293;
  wire mux_tmp_294;
  wire mux_tmp_295;
  wire mux_tmp_296;
  wire mux_tmp_297;
  wire mux_tmp_298;
  wire and_tmp_206;
  wire and_dcpl_610;
  wire or_tmp_820;
  wire and_dcpl_612;
  wire mux_tmp_301;
  wire and_dcpl_614;
  wire mux_tmp_303;
  wire mux_tmp_304;
  wire and_dcpl_616;
  wire mux_tmp_306;
  wire mux_tmp_307;
  wire mux_tmp_308;
  wire and_dcpl_618;
  wire mux_tmp_310;
  wire mux_tmp_311;
  wire mux_tmp_312;
  wire mux_tmp_313;
  wire and_dcpl_622;
  wire mux_tmp_315;
  wire mux_tmp_316;
  wire mux_tmp_317;
  wire mux_tmp_318;
  wire mux_tmp_319;
  wire and_dcpl_625;
  wire mux_tmp_321;
  wire mux_tmp_322;
  wire mux_tmp_323;
  wire mux_tmp_324;
  wire mux_tmp_325;
  wire mux_tmp_326;
  wire and_dcpl_628;
  wire mux_tmp_328;
  wire mux_tmp_329;
  wire mux_tmp_330;
  wire mux_tmp_331;
  wire mux_tmp_332;
  wire mux_tmp_333;
  wire mux_tmp_334;
  wire and_dcpl_631;
  wire mux_tmp_336;
  wire mux_tmp_337;
  wire mux_tmp_338;
  wire mux_tmp_339;
  wire mux_tmp_340;
  wire mux_tmp_341;
  wire mux_tmp_342;
  wire mux_tmp_343;
  wire and_dcpl_634;
  wire or_tmp_921;
  wire mux_tmp_345;
  wire mux_tmp_346;
  wire mux_tmp_347;
  wire mux_tmp_348;
  wire mux_tmp_349;
  wire mux_tmp_350;
  wire mux_tmp_351;
  wire mux_tmp_352;
  wire mux_tmp_353;
  wire mux_tmp_354;
  wire and_dcpl_638;
  wire and_dcpl_639;
  wire or_tmp_934;
  wire and_dcpl_641;
  wire and_dcpl_642;
  wire and_tmp_207;
  wire and_dcpl_644;
  wire and_dcpl_645;
  wire and_tmp_209;
  wire and_dcpl_647;
  wire and_dcpl_648;
  wire and_tmp_212;
  wire and_dcpl_650;
  wire and_tmp_216;
  wire and_dcpl_653;
  wire and_tmp_220;
  wire and_dcpl_657;
  wire mux_tmp_362;
  wire and_tmp_224;
  wire and_dcpl_661;
  wire mux_tmp_365;
  wire mux_tmp_366;
  wire and_tmp_228;
  wire and_dcpl_665;
  wire mux_tmp_369;
  wire mux_tmp_370;
  wire mux_tmp_371;
  wire and_tmp_232;
  wire and_dcpl_669;
  wire or_tmp_1009;
  wire mux_tmp_374;
  wire mux_tmp_375;
  wire mux_tmp_376;
  wire mux_tmp_377;
  wire mux_tmp_378;
  wire mux_tmp_379;
  wire mux_tmp_380;
  wire mux_tmp_381;
  wire and_tmp_233;
  wire and_dcpl_673;
  wire or_tmp_1021;
  wire and_dcpl_675;
  wire mux_tmp_384;
  wire and_dcpl_677;
  wire mux_tmp_386;
  wire mux_tmp_387;
  wire and_dcpl_679;
  wire mux_tmp_389;
  wire mux_tmp_390;
  wire mux_tmp_391;
  wire and_dcpl_681;
  wire mux_tmp_393;
  wire mux_tmp_394;
  wire mux_tmp_395;
  wire mux_tmp_396;
  wire and_dcpl_684;
  wire mux_tmp_398;
  wire mux_tmp_399;
  wire mux_tmp_400;
  wire mux_tmp_401;
  wire mux_tmp_402;
  wire and_dcpl_687;
  wire mux_tmp_404;
  wire mux_tmp_405;
  wire mux_tmp_406;
  wire mux_tmp_407;
  wire mux_tmp_408;
  wire mux_tmp_409;
  wire and_dcpl_690;
  wire mux_tmp_411;
  wire mux_tmp_412;
  wire mux_tmp_413;
  wire mux_tmp_414;
  wire mux_tmp_415;
  wire mux_tmp_416;
  wire mux_tmp_417;
  wire and_dcpl_693;
  wire mux_tmp_419;
  wire mux_tmp_420;
  wire mux_tmp_421;
  wire mux_tmp_422;
  wire mux_tmp_423;
  wire mux_tmp_424;
  wire mux_tmp_425;
  wire mux_tmp_426;
  wire and_dcpl_696;
  wire or_tmp_1122;
  wire mux_tmp_428;
  wire mux_tmp_429;
  wire mux_tmp_430;
  wire mux_tmp_431;
  wire mux_tmp_432;
  wire mux_tmp_433;
  wire mux_tmp_434;
  wire mux_tmp_435;
  wire mux_tmp_436;
  wire mux_tmp_437;
  reg [1:0] rem_12cyc_st_10_1_0;
  reg [1:0] rem_12cyc_st_10_3_2;
  reg [1:0] rem_12cyc_st_9_1_0;
  reg [1:0] rem_12cyc_st_9_3_2;
  reg [1:0] rem_12cyc_st_8_1_0;
  reg [1:0] rem_12cyc_st_8_3_2;
  reg [1:0] rem_12cyc_st_7_1_0;
  reg [1:0] rem_12cyc_st_7_3_2;
  reg [1:0] rem_12cyc_st_6_1_0;
  reg [1:0] rem_12cyc_st_6_3_2;
  reg [1:0] rem_12cyc_st_5_1_0;
  reg [1:0] rem_12cyc_st_5_3_2;
  reg [1:0] rem_12cyc_st_4_1_0;
  reg [1:0] rem_12cyc_st_4_3_2;
  reg [1:0] rem_12cyc_st_3_1_0;
  reg [1:0] rem_12cyc_st_3_3_2;
  reg [1:0] rem_12cyc_st_2_1_0;
  reg [1:0] rem_12cyc_st_2_3_2;
  reg [1:0] rem_12cyc_1_0;
  reg [1:0] rem_12cyc_3_2;
  reg [1:0] rem_12cyc_st_12_3_2;
  reg [63:0] result_sva_duc;
  reg [1:0] rem_12cyc_st_12_1_0;
  reg asn_itm_12;
  reg main_stage_0_13;
  reg main_stage_0_3;
  reg asn_itm_1;
  reg main_stage_0_2;
  reg main_stage_0_4;
  reg asn_itm_2;
  reg main_stage_0_5;
  reg asn_itm_3;
  reg main_stage_0_6;
  reg asn_itm_4;
  reg asn_itm_5;
  reg main_stage_0_8;
  reg asn_itm_7;
  reg main_stage_0_9;
  reg asn_itm_8;
  reg main_stage_0_10;
  reg asn_itm_9;
  reg main_stage_0_7;
  reg asn_itm_6;
  reg main_stage_0_11;
  reg asn_itm_10;
  wire and_1173_cse;
  wire and_1175_cse;
  wire and_1177_cse;
  wire and_1179_cse;
  wire and_1181_cse;
  wire and_1183_cse;
  wire and_1185_cse;
  wire and_1187_cse;
  wire and_1189_cse;
  wire and_1191_cse;
  wire and_1193_cse;
  wire and_1195_cse;
  wire and_1197_cse;
  wire or_1_cse;
  wire or_6_cse;
  wire or_10_cse;
  wire or_15_cse;
  wire or_21_cse;
  wire or_28_cse;
  wire or_37_cse;
  wire or_48_cse;
  wire or_83_cse;
  wire nand_276_cse;
  wire or_88_cse;
  wire nand_274_cse;
  wire or_93_cse;
  wire nand_271_cse;
  wire or_100_cse;
  wire nand_267_cse;
  wire or_109_cse;
  wire or_120_cse;
  wire or_133_cse;
  wire or_148_cse;
  wire or_190_cse;
  wire or_195_cse;
  wire or_199_cse;
  wire or_204_cse;
  wire or_210_cse;
  wire or_217_cse;
  wire or_226_cse;
  wire or_237_cse;
  wire or_270_cse;
  wire or_275_cse;
  wire or_280_cse;
  wire or_287_cse;
  wire or_296_cse;
  wire or_307_cse;
  wire or_320_cse;
  wire or_335_cse;
  wire nand_281_cse;
  wire or_377_cse;
  wire or_382_cse;
  wire or_386_cse;
  wire or_391_cse;
  wire or_397_cse;
  wire nand_215_cse;
  wire or_404_cse;
  wire nand_212_cse;
  wire or_413_cse;
  wire nand_208_cse;
  wire or_424_cse;
  wire or_458_cse;
  wire or_463_cse;
  wire nand_198_cse;
  wire or_468_cse;
  wire or_475_cse;
  wire nand_189_cse;
  wire or_484_cse;
  wire or_495_cse;
  wire or_508_cse;
  wire nand_203_cse;
  wire or_523_cse;
  wire nand_250_cse;
  wire or_564_cse;
  wire or_569_cse;
  wire or_573_cse;
  wire or_578_cse;
  wire or_584_cse;
  wire or_591_cse;
  wire or_600_cse;
  wire or_611_cse;
  wire or_643_cse;
  wire or_648_cse;
  wire or_653_cse;
  wire or_660_cse;
  wire or_669_cse;
  wire or_680_cse;
  wire or_693_cse;
  wire or_708_cse;
  wire or_748_cse;
  wire or_753_cse;
  wire or_757_cse;
  wire or_762_cse;
  wire or_768_cse;
  wire or_775_cse;
  wire or_784_cse;
  wire or_795_cse;
  wire or_837_cse;
  wire nand_84_cse;
  wire or_842_cse;
  wire or_847_cse;
  wire nand_79_cse;
  wire or_854_cse;
  wire or_863_cse;
  wire or_874_cse;
  wire or_887_cse;
  wire or_902_cse;
  wire or_952_cse;
  wire or_957_cse;
  wire or_961_cse;
  wire or_966_cse;
  wire or_972_cse;
  wire or_979_cse;
  wire or_988_cse;
  wire or_999_cse;
  wire nand_57_cse;
  wire or_1045_cse;
  wire or_1050_cse;
  wire or_1057_cse;
  wire or_1066_cse;
  wire nand_36_cse;
  wire nand_29_cse;
  wire nand_21_cse;
  wire nand_222_cse;
  wire nand_223_cse;
  reg main_stage_0_12;
  reg [63:0] m_buf_sva_1;
  reg [63:0] m_buf_sva_2;
  reg [63:0] m_buf_sva_3;
  reg [63:0] m_buf_sva_4;
  reg [63:0] m_buf_sva_5;
  reg [63:0] m_buf_sva_6;
  reg [63:0] m_buf_sva_7;
  reg [63:0] m_buf_sva_8;
  reg [63:0] m_buf_sva_9;
  reg [63:0] m_buf_sva_10;
  reg [63:0] m_buf_sva_11;
  reg [63:0] m_buf_sva_12;
  reg asn_itm_11;
  reg [63:0] mut_2_63_0;
  reg [63:0] mut_3_63_0;
  reg [63:0] mut_4_63_0;
  reg [63:0] mut_5_63_0;
  reg [63:0] mut_6_63_0;
  reg [63:0] mut_7_63_0;
  reg [63:0] mut_8_63_0;
  reg [63:0] mut_9_63_0;
  reg [63:0] mut_10_63_0;
  reg [63:0] mut_11_63_0;
  reg [63:0] mut_1_2_63_0;
  reg [63:0] mut_1_3_63_0;
  reg [63:0] mut_1_4_63_0;
  reg [63:0] mut_1_5_63_0;
  reg [63:0] mut_1_6_63_0;
  reg [63:0] mut_1_7_63_0;
  reg [63:0] mut_1_8_63_0;
  reg [63:0] mut_1_9_63_0;
  reg [63:0] mut_1_10_63_0;
  reg [63:0] mut_1_11_63_0;
  reg [63:0] mut_2_2_63_0;
  reg [63:0] mut_2_3_63_0;
  reg [63:0] mut_2_4_63_0;
  reg [63:0] mut_2_5_63_0;
  reg [63:0] mut_2_6_63_0;
  reg [63:0] mut_2_7_63_0;
  reg [63:0] mut_2_8_63_0;
  reg [63:0] mut_2_9_63_0;
  reg [63:0] mut_2_10_63_0;
  reg [63:0] mut_2_11_63_0;
  reg [63:0] mut_3_2_63_0;
  reg [63:0] mut_3_3_63_0;
  reg [63:0] mut_3_4_63_0;
  reg [63:0] mut_3_5_63_0;
  reg [63:0] mut_3_6_63_0;
  reg [63:0] mut_3_7_63_0;
  reg [63:0] mut_3_8_63_0;
  reg [63:0] mut_3_9_63_0;
  reg [63:0] mut_3_10_63_0;
  reg [63:0] mut_3_11_63_0;
  reg [63:0] mut_4_2_63_0;
  reg [63:0] mut_4_3_63_0;
  reg [63:0] mut_4_4_63_0;
  reg [63:0] mut_4_5_63_0;
  reg [63:0] mut_4_6_63_0;
  reg [63:0] mut_4_7_63_0;
  reg [63:0] mut_4_8_63_0;
  reg [63:0] mut_4_9_63_0;
  reg [63:0] mut_4_10_63_0;
  reg [63:0] mut_4_11_63_0;
  reg [63:0] mut_5_2_63_0;
  reg [63:0] mut_5_3_63_0;
  reg [63:0] mut_5_4_63_0;
  reg [63:0] mut_5_5_63_0;
  reg [63:0] mut_5_6_63_0;
  reg [63:0] mut_5_7_63_0;
  reg [63:0] mut_5_8_63_0;
  reg [63:0] mut_5_9_63_0;
  reg [63:0] mut_5_10_63_0;
  reg [63:0] mut_5_11_63_0;
  reg [63:0] mut_6_2_63_0;
  reg [63:0] mut_6_3_63_0;
  reg [63:0] mut_6_4_63_0;
  reg [63:0] mut_6_5_63_0;
  reg [63:0] mut_6_6_63_0;
  reg [63:0] mut_6_7_63_0;
  reg [63:0] mut_6_8_63_0;
  reg [63:0] mut_6_9_63_0;
  reg [63:0] mut_6_10_63_0;
  reg [63:0] mut_6_11_63_0;
  reg [63:0] mut_7_2_63_0;
  reg [63:0] mut_7_3_63_0;
  reg [63:0] mut_7_4_63_0;
  reg [63:0] mut_7_5_63_0;
  reg [63:0] mut_7_6_63_0;
  reg [63:0] mut_7_7_63_0;
  reg [63:0] mut_7_8_63_0;
  reg [63:0] mut_7_9_63_0;
  reg [63:0] mut_7_10_63_0;
  reg [63:0] mut_7_11_63_0;
  reg [63:0] mut_8_2_63_0;
  reg [63:0] mut_8_3_63_0;
  reg [63:0] mut_8_4_63_0;
  reg [63:0] mut_8_5_63_0;
  reg [63:0] mut_8_6_63_0;
  reg [63:0] mut_8_7_63_0;
  reg [63:0] mut_8_8_63_0;
  reg [63:0] mut_8_9_63_0;
  reg [63:0] mut_8_10_63_0;
  reg [63:0] mut_8_11_63_0;
  reg [63:0] mut_9_2_63_0;
  reg [63:0] mut_9_3_63_0;
  reg [63:0] mut_9_4_63_0;
  reg [63:0] mut_9_5_63_0;
  reg [63:0] mut_9_6_63_0;
  reg [63:0] mut_9_7_63_0;
  reg [63:0] mut_9_8_63_0;
  reg [63:0] mut_9_9_63_0;
  reg [63:0] mut_9_10_63_0;
  reg [63:0] mut_9_11_63_0;
  reg [63:0] mut_10_2_63_0;
  reg [63:0] mut_10_3_63_0;
  reg [63:0] mut_10_4_63_0;
  reg [63:0] mut_10_5_63_0;
  reg [63:0] mut_10_6_63_0;
  reg [63:0] mut_10_7_63_0;
  reg [63:0] mut_10_8_63_0;
  reg [63:0] mut_10_9_63_0;
  reg [63:0] mut_10_10_63_0;
  reg [63:0] mut_10_11_63_0;
  reg [63:0] mut_11_2_63_0;
  reg [63:0] mut_11_3_63_0;
  reg [63:0] mut_11_4_63_0;
  reg [63:0] mut_11_5_63_0;
  reg [63:0] mut_11_6_63_0;
  reg [63:0] mut_11_7_63_0;
  reg [63:0] mut_11_8_63_0;
  reg [63:0] mut_11_9_63_0;
  reg [63:0] mut_11_10_63_0;
  reg [63:0] mut_11_11_63_0;
  reg [63:0] mut_12_2_63_0;
  reg [63:0] mut_12_3_63_0;
  reg [63:0] mut_12_4_63_0;
  reg [63:0] mut_12_5_63_0;
  reg [63:0] mut_12_6_63_0;
  reg [63:0] mut_12_7_63_0;
  reg [63:0] mut_12_8_63_0;
  reg [63:0] mut_12_9_63_0;
  reg [63:0] mut_12_10_63_0;
  reg [63:0] mut_12_11_63_0;
  reg [63:0] mut_13_2_63_0;
  reg [63:0] mut_13_3_63_0;
  reg [63:0] mut_13_4_63_0;
  reg [63:0] mut_13_5_63_0;
  reg [63:0] mut_13_6_63_0;
  reg [63:0] mut_13_7_63_0;
  reg [63:0] mut_13_8_63_0;
  reg [63:0] mut_13_9_63_0;
  reg [63:0] mut_13_10_63_0;
  reg [63:0] mut_13_11_63_0;
  reg [63:0] mut_14_2_63_0;
  reg [63:0] mut_14_3_63_0;
  reg [63:0] mut_14_4_63_0;
  reg [63:0] mut_14_5_63_0;
  reg [63:0] mut_14_6_63_0;
  reg [63:0] mut_14_7_63_0;
  reg [63:0] mut_14_8_63_0;
  reg [63:0] mut_14_9_63_0;
  reg [63:0] mut_14_10_63_0;
  reg [63:0] mut_14_11_63_0;
  reg [63:0] mut_15_2_63_0;
  reg [63:0] mut_15_3_63_0;
  reg [63:0] mut_15_4_63_0;
  reg [63:0] mut_15_5_63_0;
  reg [63:0] mut_15_6_63_0;
  reg [63:0] mut_15_7_63_0;
  reg [63:0] mut_15_8_63_0;
  reg [63:0] mut_15_9_63_0;
  reg [63:0] mut_15_10_63_0;
  reg [63:0] mut_15_11_63_0;
  reg [63:0] mut_16_2_63_0;
  reg [63:0] mut_16_3_63_0;
  reg [63:0] mut_16_4_63_0;
  reg [63:0] mut_16_5_63_0;
  reg [63:0] mut_16_6_63_0;
  reg [63:0] mut_16_7_63_0;
  reg [63:0] mut_16_8_63_0;
  reg [63:0] mut_16_9_63_0;
  reg [63:0] mut_16_10_63_0;
  reg [63:0] mut_16_11_63_0;
  reg [63:0] mut_17_2_63_0;
  reg [63:0] mut_17_3_63_0;
  reg [63:0] mut_17_4_63_0;
  reg [63:0] mut_17_5_63_0;
  reg [63:0] mut_17_6_63_0;
  reg [63:0] mut_17_7_63_0;
  reg [63:0] mut_17_8_63_0;
  reg [63:0] mut_17_9_63_0;
  reg [63:0] mut_17_10_63_0;
  reg [63:0] mut_17_11_63_0;
  reg [63:0] mut_18_2_63_0;
  reg [63:0] mut_18_3_63_0;
  reg [63:0] mut_18_4_63_0;
  reg [63:0] mut_18_5_63_0;
  reg [63:0] mut_18_6_63_0;
  reg [63:0] mut_18_7_63_0;
  reg [63:0] mut_18_8_63_0;
  reg [63:0] mut_18_9_63_0;
  reg [63:0] mut_18_10_63_0;
  reg [63:0] mut_18_11_63_0;
  reg [63:0] mut_19_2_63_0;
  reg [63:0] mut_19_3_63_0;
  reg [63:0] mut_19_4_63_0;
  reg [63:0] mut_19_5_63_0;
  reg [63:0] mut_19_6_63_0;
  reg [63:0] mut_19_7_63_0;
  reg [63:0] mut_19_8_63_0;
  reg [63:0] mut_19_9_63_0;
  reg [63:0] mut_19_10_63_0;
  reg [63:0] mut_19_11_63_0;
  reg [63:0] mut_20_2_63_0;
  reg [63:0] mut_20_3_63_0;
  reg [63:0] mut_20_4_63_0;
  reg [63:0] mut_20_5_63_0;
  reg [63:0] mut_20_6_63_0;
  reg [63:0] mut_20_7_63_0;
  reg [63:0] mut_20_8_63_0;
  reg [63:0] mut_20_9_63_0;
  reg [63:0] mut_20_10_63_0;
  reg [63:0] mut_20_11_63_0;
  reg [63:0] mut_21_2_63_0;
  reg [63:0] mut_21_3_63_0;
  reg [63:0] mut_21_4_63_0;
  reg [63:0] mut_21_5_63_0;
  reg [63:0] mut_21_6_63_0;
  reg [63:0] mut_21_7_63_0;
  reg [63:0] mut_21_8_63_0;
  reg [63:0] mut_21_9_63_0;
  reg [63:0] mut_21_10_63_0;
  reg [63:0] mut_21_11_63_0;
  reg [63:0] mut_22_2_63_0;
  reg [63:0] mut_22_3_63_0;
  reg [63:0] mut_22_4_63_0;
  reg [63:0] mut_22_5_63_0;
  reg [63:0] mut_22_6_63_0;
  reg [63:0] mut_22_7_63_0;
  reg [63:0] mut_22_8_63_0;
  reg [63:0] mut_22_9_63_0;
  reg [63:0] mut_22_10_63_0;
  reg [63:0] mut_22_11_63_0;
  reg [63:0] mut_23_2_63_0;
  reg [63:0] mut_23_3_63_0;
  reg [63:0] mut_23_4_63_0;
  reg [63:0] mut_23_5_63_0;
  reg [63:0] mut_23_6_63_0;
  reg [63:0] mut_23_7_63_0;
  reg [63:0] mut_23_8_63_0;
  reg [63:0] mut_23_9_63_0;
  reg [63:0] mut_23_10_63_0;
  reg [63:0] mut_23_11_63_0;
  reg [1:0] rem_12cyc_st_11_3_2;
  reg [1:0] rem_12cyc_st_11_1_0;
  wire [63:0] result_sva_duc_mx0;
  wire and_1203_cse;
  wire and_1205_cse;
  wire and_1207_cse;
  wire and_1209_cse;
  wire and_1211_cse;
  wire and_1213_cse;
  wire and_1215_cse;
  wire and_1217_cse;
  wire and_1219_cse;
  wire and_1221_cse;
  wire and_1223_cse;
  wire and_1225_cse;
  wire and_1227_cse;
  wire and_1229_cse;
  wire and_1231_cse;
  wire and_1233_cse;
  wire and_1235_cse;
  wire and_1237_cse;
  wire and_1239_cse;
  wire and_1241_cse;
  wire and_1243_cse;
  wire and_1245_cse;
  wire and_1247_cse;
  wire and_1249_cse;
  wire and_1251_cse;
  wire and_1253_cse;
  wire and_1255_cse;
  wire and_1257_cse;
  wire and_1259_cse;
  wire and_1261_cse;
  wire and_1263_cse;
  wire and_1265_cse;
  wire and_1267_cse;
  wire and_1269_cse;
  wire and_1271_cse;
  wire and_1273_cse;
  wire and_1275_cse;
  wire and_1277_cse;
  wire and_1279_cse;
  wire and_1281_cse;
  wire and_1283_cse;
  wire and_1285_cse;
  wire and_1287_cse;
  wire and_1289_cse;
  wire and_1291_cse;
  wire and_1293_cse;
  wire and_1295_cse;
  wire and_1297_cse;
  wire and_1299_cse;
  wire and_1301_cse;
  wire and_1303_cse;
  wire and_1305_cse;
  wire and_1307_cse;
  wire and_1309_cse;
  wire and_1311_cse;
  wire and_1313_cse;
  wire and_1315_cse;
  wire and_1317_cse;
  wire and_1319_cse;
  wire and_1321_cse;
  wire and_1323_cse;
  wire and_1325_cse;
  wire and_1327_cse;
  wire and_1329_cse;
  wire and_1331_cse;
  wire and_1333_cse;
  wire and_1335_cse;
  wire and_1337_cse;
  wire and_1339_cse;
  wire and_1341_cse;
  wire and_1343_cse;
  wire and_1345_cse;
  wire and_1347_cse;
  wire and_1349_cse;
  wire and_1351_cse;
  wire and_1353_cse;
  wire and_1355_cse;
  wire and_1357_cse;
  wire and_1359_cse;
  wire and_1361_cse;
  wire and_1363_cse;
  wire and_1365_cse;
  wire and_1367_cse;
  wire and_1369_cse;
  wire and_1371_cse;
  wire and_1373_cse;
  wire and_1375_cse;
  wire and_1377_cse;
  wire and_1379_cse;
  wire and_1381_cse;
  wire and_1383_cse;
  wire and_1385_cse;
  wire and_1387_cse;
  wire and_1389_cse;
  wire and_1391_cse;
  wire and_1393_cse;
  wire and_1395_cse;
  wire and_1397_cse;
  wire and_1399_cse;
  wire and_1401_cse;
  wire and_1403_cse;
  wire and_1405_cse;
  wire and_1407_cse;
  wire and_1409_cse;
  wire and_1411_cse;
  wire and_1413_cse;
  wire and_1415_cse;
  wire and_1417_cse;
  wire and_1419_cse;
  wire and_1421_cse;
  wire and_1423_cse;
  wire and_1425_cse;
  wire and_1427_cse;
  wire and_1429_cse;
  wire and_1431_cse;
  wire and_1433_cse;
  wire and_1435_cse;
  wire and_1437_cse;
  wire and_1439_cse;
  wire and_1441_cse;
  wire and_1443_cse;
  wire and_1445_cse;
  wire and_1447_cse;
  wire and_1449_cse;
  wire and_1451_cse;
  wire and_1453_cse;
  wire and_1455_cse;
  wire and_1457_cse;
  wire and_1459_cse;
  wire and_1461_cse;
  wire and_1463_cse;

  wire[63:0] qelse_acc_nl;
  wire[64:0] nl_qelse_acc_nl;
  wire[0:0] mux_13_nl;
  wire[0:0] mux_12_nl;
  wire[0:0] mux_11_nl;
  wire[0:0] mux_10_nl;
  wire[0:0] mux_9_nl;
  wire[0:0] mux_8_nl;
  wire[0:0] mux_7_nl;
  wire[0:0] mux_6_nl;
  wire[0:0] mux_5_nl;
  wire[0:0] mux_4_nl;
  wire[0:0] mux_3_nl;
  wire[0:0] mux_2_nl;
  wire[0:0] and_273_nl;
  wire[0:0] and_275_nl;
  wire[0:0] and_277_nl;
  wire[0:0] and_279_nl;
  wire[0:0] and_281_nl;
  wire[0:0] and_282_nl;
  wire[0:0] and_283_nl;
  wire[0:0] and_284_nl;
  wire[0:0] and_286_nl;
  wire[0:0] and_287_nl;
  wire[0:0] and_288_nl;
  wire[0:0] and_289_nl;
  wire[0:0] and_290_nl;
  wire[0:0] xor_nl;
  wire[0:0] nor_nl;
  wire[0:0] mux_14_nl;
  wire[0:0] nor_518_nl;
  wire[0:0] mux_15_nl;
  wire[0:0] nor_517_nl;
  wire[0:0] mux_16_nl;
  wire[0:0] nor_516_nl;
  wire[0:0] mux_17_nl;
  wire[0:0] nor_515_nl;
  wire[0:0] mux_18_nl;
  wire[0:0] nor_514_nl;
  wire[0:0] mux_19_nl;
  wire[0:0] nor_512_nl;
  wire[0:0] mux_20_nl;
  wire[0:0] nor_513_nl;
  wire[0:0] nor_509_nl;
  wire[0:0] mux_22_nl;
  wire[0:0] nor_510_nl;
  wire[0:0] mux_23_nl;
  wire[0:0] nor_511_nl;
  wire[0:0] nor_505_nl;
  wire[0:0] nor_506_nl;
  wire[0:0] mux_26_nl;
  wire[0:0] nor_507_nl;
  wire[0:0] mux_27_nl;
  wire[0:0] nor_508_nl;
  wire[0:0] nor_500_nl;
  wire[0:0] or_61_nl;
  wire[0:0] nor_501_nl;
  wire[0:0] nor_502_nl;
  wire[0:0] mux_31_nl;
  wire[0:0] nor_503_nl;
  wire[0:0] mux_32_nl;
  wire[0:0] nor_504_nl;
  wire[0:0] mux_33_nl;
  wire[0:0] nor_499_nl;
  wire[0:0] and_1168_nl;
  wire[0:0] mux_35_nl;
  wire[0:0] nor_498_nl;
  wire[0:0] and_1166_nl;
  wire[0:0] and_1167_nl;
  wire[0:0] mux_38_nl;
  wire[0:0] nor_497_nl;
  wire[0:0] and_1163_nl;
  wire[0:0] and_1164_nl;
  wire[0:0] and_1165_nl;
  wire[0:0] mux_42_nl;
  wire[0:0] nor_496_nl;
  wire[0:0] and_1159_nl;
  wire[0:0] and_1160_nl;
  wire[0:0] and_1161_nl;
  wire[0:0] and_1162_nl;
  wire[0:0] mux_47_nl;
  wire[0:0] nor_495_nl;
  wire[0:0] nor_493_nl;
  wire[0:0] and_1155_nl;
  wire[0:0] and_1156_nl;
  wire[0:0] and_1157_nl;
  wire[0:0] and_1158_nl;
  wire[0:0] mux_53_nl;
  wire[0:0] nor_494_nl;
  wire[0:0] nor_490_nl;
  wire[0:0] nor_491_nl;
  wire[0:0] and_1151_nl;
  wire[0:0] and_1152_nl;
  wire[0:0] and_1153_nl;
  wire[0:0] and_1154_nl;
  wire[0:0] mux_60_nl;
  wire[0:0] nor_492_nl;
  wire[0:0] nor_486_nl;
  wire[0:0] nor_487_nl;
  wire[0:0] nor_488_nl;
  wire[0:0] and_1147_nl;
  wire[0:0] and_1148_nl;
  wire[0:0] and_1149_nl;
  wire[0:0] and_1150_nl;
  wire[0:0] mux_68_nl;
  wire[0:0] nor_489_nl;
  wire[0:0] nor_481_nl;
  wire[0:0] or_165_nl;
  wire[0:0] nor_482_nl;
  wire[0:0] nor_483_nl;
  wire[0:0] nor_484_nl;
  wire[0:0] and_1143_nl;
  wire[0:0] and_1144_nl;
  wire[0:0] and_1145_nl;
  wire[0:0] and_1146_nl;
  wire[0:0] mux_77_nl;
  wire[0:0] nor_485_nl;
  wire[0:0] nor_480_nl;
  wire[0:0] or_175_nl;
  wire[0:0] mux_79_nl;
  wire[0:0] nor_479_nl;
  wire[0:0] mux_80_nl;
  wire[0:0] nor_478_nl;
  wire[0:0] mux_81_nl;
  wire[0:0] nor_477_nl;
  wire[0:0] mux_82_nl;
  wire[0:0] nor_476_nl;
  wire[0:0] mux_83_nl;
  wire[0:0] nor_475_nl;
  wire[0:0] mux_84_nl;
  wire[0:0] nor_473_nl;
  wire[0:0] mux_85_nl;
  wire[0:0] nor_474_nl;
  wire[0:0] nor_470_nl;
  wire[0:0] mux_87_nl;
  wire[0:0] nor_471_nl;
  wire[0:0] mux_88_nl;
  wire[0:0] nor_472_nl;
  wire[0:0] nor_466_nl;
  wire[0:0] nor_467_nl;
  wire[0:0] mux_91_nl;
  wire[0:0] nor_468_nl;
  wire[0:0] mux_92_nl;
  wire[0:0] nor_469_nl;
  wire[0:0] nor_461_nl;
  wire[0:0] or_250_nl;
  wire[0:0] nor_462_nl;
  wire[0:0] nor_463_nl;
  wire[0:0] mux_96_nl;
  wire[0:0] nor_464_nl;
  wire[0:0] mux_97_nl;
  wire[0:0] nor_465_nl;
  wire[0:0] mux_98_nl;
  wire[0:0] nor_460_nl;
  wire[0:0] and_1142_nl;
  wire[0:0] mux_100_nl;
  wire[0:0] nor_459_nl;
  wire[0:0] and_1140_nl;
  wire[0:0] and_1141_nl;
  wire[0:0] mux_103_nl;
  wire[0:0] nor_458_nl;
  wire[0:0] and_1137_nl;
  wire[0:0] and_1138_nl;
  wire[0:0] and_1139_nl;
  wire[0:0] mux_107_nl;
  wire[0:0] nor_457_nl;
  wire[0:0] and_1133_nl;
  wire[0:0] and_1134_nl;
  wire[0:0] and_1135_nl;
  wire[0:0] and_1136_nl;
  wire[0:0] mux_112_nl;
  wire[0:0] nor_456_nl;
  wire[0:0] nor_454_nl;
  wire[0:0] and_1129_nl;
  wire[0:0] and_1130_nl;
  wire[0:0] and_1131_nl;
  wire[0:0] and_1132_nl;
  wire[0:0] mux_118_nl;
  wire[0:0] nor_455_nl;
  wire[0:0] nor_451_nl;
  wire[0:0] nor_452_nl;
  wire[0:0] and_1125_nl;
  wire[0:0] and_1126_nl;
  wire[0:0] and_1127_nl;
  wire[0:0] and_1128_nl;
  wire[0:0] mux_125_nl;
  wire[0:0] nor_453_nl;
  wire[0:0] nor_447_nl;
  wire[0:0] nor_448_nl;
  wire[0:0] nor_449_nl;
  wire[0:0] and_1121_nl;
  wire[0:0] and_1122_nl;
  wire[0:0] and_1123_nl;
  wire[0:0] and_1124_nl;
  wire[0:0] mux_133_nl;
  wire[0:0] nor_450_nl;
  wire[0:0] nor_442_nl;
  wire[0:0] or_352_nl;
  wire[0:0] nor_443_nl;
  wire[0:0] nor_444_nl;
  wire[0:0] nor_445_nl;
  wire[0:0] and_1117_nl;
  wire[0:0] and_1118_nl;
  wire[0:0] and_1119_nl;
  wire[0:0] and_1120_nl;
  wire[0:0] mux_142_nl;
  wire[0:0] nor_446_nl;
  wire[0:0] and_1116_nl;
  wire[0:0] or_362_nl;
  wire[0:0] mux_144_nl;
  wire[0:0] and_1172_nl;
  wire[0:0] mux_145_nl;
  wire[0:0] and_1114_nl;
  wire[0:0] mux_146_nl;
  wire[0:0] and_1113_nl;
  wire[0:0] mux_147_nl;
  wire[0:0] and_1112_nl;
  wire[0:0] mux_148_nl;
  wire[0:0] and_1111_nl;
  wire[0:0] mux_149_nl;
  wire[0:0] and_1109_nl;
  wire[0:0] mux_150_nl;
  wire[0:0] and_1110_nl;
  wire[0:0] and_1106_nl;
  wire[0:0] mux_152_nl;
  wire[0:0] and_1107_nl;
  wire[0:0] mux_153_nl;
  wire[0:0] and_1108_nl;
  wire[0:0] and_1102_nl;
  wire[0:0] and_1103_nl;
  wire[0:0] mux_156_nl;
  wire[0:0] and_1104_nl;
  wire[0:0] mux_157_nl;
  wire[0:0] and_1105_nl;
  wire[0:0] and_1097_nl;
  wire[0:0] or_437_nl;
  wire[0:0] and_1098_nl;
  wire[0:0] and_1099_nl;
  wire[0:0] mux_161_nl;
  wire[0:0] and_1100_nl;
  wire[0:0] mux_162_nl;
  wire[0:0] and_1101_nl;
  wire[0:0] mux_163_nl;
  wire[0:0] and_1171_nl;
  wire[0:0] and_1094_nl;
  wire[0:0] mux_165_nl;
  wire[0:0] and_1095_nl;
  wire[0:0] and_1091_nl;
  wire[0:0] and_1092_nl;
  wire[0:0] mux_168_nl;
  wire[0:0] and_1093_nl;
  wire[0:0] and_1087_nl;
  wire[0:0] and_1088_nl;
  wire[0:0] and_1089_nl;
  wire[0:0] mux_172_nl;
  wire[0:0] and_1090_nl;
  wire[0:0] and_1082_nl;
  wire[0:0] and_1083_nl;
  wire[0:0] and_1084_nl;
  wire[0:0] and_1085_nl;
  wire[0:0] mux_177_nl;
  wire[0:0] and_1086_nl;
  wire[0:0] and_1076_nl;
  wire[0:0] and_1077_nl;
  wire[0:0] and_1078_nl;
  wire[0:0] and_1079_nl;
  wire[0:0] and_1080_nl;
  wire[0:0] mux_183_nl;
  wire[0:0] and_1081_nl;
  wire[0:0] and_1069_nl;
  wire[0:0] and_1070_nl;
  wire[0:0] and_1071_nl;
  wire[0:0] and_1072_nl;
  wire[0:0] and_1073_nl;
  wire[0:0] and_1074_nl;
  wire[0:0] mux_190_nl;
  wire[0:0] and_1075_nl;
  wire[0:0] and_1061_nl;
  wire[0:0] and_1062_nl;
  wire[0:0] and_1063_nl;
  wire[0:0] and_1064_nl;
  wire[0:0] and_1065_nl;
  wire[0:0] and_1066_nl;
  wire[0:0] and_1067_nl;
  wire[0:0] mux_198_nl;
  wire[0:0] and_1068_nl;
  wire[0:0] and_1052_nl;
  wire[0:0] or_540_nl;
  wire[0:0] and_1053_nl;
  wire[0:0] and_1054_nl;
  wire[0:0] and_1055_nl;
  wire[0:0] and_1056_nl;
  wire[0:0] and_1057_nl;
  wire[0:0] and_1058_nl;
  wire[0:0] and_1059_nl;
  wire[0:0] mux_207_nl;
  wire[0:0] and_1060_nl;
  wire[0:0] nor_439_nl;
  wire[0:0] or_550_nl;
  wire[0:0] mux_209_nl;
  wire[0:0] and_1170_nl;
  wire[0:0] mux_210_nl;
  wire[0:0] and_1050_nl;
  wire[0:0] mux_211_nl;
  wire[0:0] and_1049_nl;
  wire[0:0] mux_212_nl;
  wire[0:0] and_1048_nl;
  wire[0:0] mux_213_nl;
  wire[0:0] and_1047_nl;
  wire[0:0] mux_214_nl;
  wire[0:0] and_1045_nl;
  wire[0:0] mux_215_nl;
  wire[0:0] and_1046_nl;
  wire[0:0] and_1042_nl;
  wire[0:0] mux_217_nl;
  wire[0:0] and_1043_nl;
  wire[0:0] mux_218_nl;
  wire[0:0] and_1044_nl;
  wire[0:0] and_1038_nl;
  wire[0:0] and_1039_nl;
  wire[0:0] mux_221_nl;
  wire[0:0] and_1040_nl;
  wire[0:0] mux_222_nl;
  wire[0:0] and_1041_nl;
  wire[0:0] and_1033_nl;
  wire[0:0] or_624_nl;
  wire[0:0] and_1034_nl;
  wire[0:0] and_1035_nl;
  wire[0:0] mux_226_nl;
  wire[0:0] and_1036_nl;
  wire[0:0] mux_227_nl;
  wire[0:0] and_1037_nl;
  wire[0:0] mux_228_nl;
  wire[0:0] and_1169_nl;
  wire[0:0] and_1030_nl;
  wire[0:0] mux_230_nl;
  wire[0:0] and_1031_nl;
  wire[0:0] and_1027_nl;
  wire[0:0] and_1028_nl;
  wire[0:0] mux_233_nl;
  wire[0:0] and_1029_nl;
  wire[0:0] and_1023_nl;
  wire[0:0] and_1024_nl;
  wire[0:0] and_1025_nl;
  wire[0:0] mux_237_nl;
  wire[0:0] and_1026_nl;
  wire[0:0] and_1018_nl;
  wire[0:0] and_1019_nl;
  wire[0:0] and_1020_nl;
  wire[0:0] and_1021_nl;
  wire[0:0] mux_242_nl;
  wire[0:0] and_1022_nl;
  wire[0:0] and_1012_nl;
  wire[0:0] and_1013_nl;
  wire[0:0] and_1014_nl;
  wire[0:0] and_1015_nl;
  wire[0:0] and_1016_nl;
  wire[0:0] mux_248_nl;
  wire[0:0] and_1017_nl;
  wire[0:0] and_1005_nl;
  wire[0:0] and_1006_nl;
  wire[0:0] and_1007_nl;
  wire[0:0] and_1008_nl;
  wire[0:0] and_1009_nl;
  wire[0:0] and_1010_nl;
  wire[0:0] mux_255_nl;
  wire[0:0] and_1011_nl;
  wire[0:0] and_997_nl;
  wire[0:0] and_998_nl;
  wire[0:0] and_999_nl;
  wire[0:0] and_1000_nl;
  wire[0:0] and_1001_nl;
  wire[0:0] and_1002_nl;
  wire[0:0] and_1003_nl;
  wire[0:0] mux_263_nl;
  wire[0:0] and_1004_nl;
  wire[0:0] and_988_nl;
  wire[0:0] or_725_nl;
  wire[0:0] and_989_nl;
  wire[0:0] and_990_nl;
  wire[0:0] and_991_nl;
  wire[0:0] and_992_nl;
  wire[0:0] and_993_nl;
  wire[0:0] and_994_nl;
  wire[0:0] and_995_nl;
  wire[0:0] mux_272_nl;
  wire[0:0] and_996_nl;
  wire[0:0] and_987_nl;
  wire[0:0] or_735_nl;
  wire[0:0] mux_274_nl;
  wire[0:0] nor_436_nl;
  wire[0:0] mux_275_nl;
  wire[0:0] nor_435_nl;
  wire[0:0] mux_276_nl;
  wire[0:0] nor_434_nl;
  wire[0:0] mux_277_nl;
  wire[0:0] nor_433_nl;
  wire[0:0] mux_278_nl;
  wire[0:0] nor_432_nl;
  wire[0:0] mux_279_nl;
  wire[0:0] nor_430_nl;
  wire[0:0] mux_280_nl;
  wire[0:0] nor_431_nl;
  wire[0:0] nor_427_nl;
  wire[0:0] mux_282_nl;
  wire[0:0] nor_428_nl;
  wire[0:0] mux_283_nl;
  wire[0:0] nor_429_nl;
  wire[0:0] nor_423_nl;
  wire[0:0] nor_424_nl;
  wire[0:0] mux_286_nl;
  wire[0:0] nor_425_nl;
  wire[0:0] mux_287_nl;
  wire[0:0] nor_426_nl;
  wire[0:0] nor_418_nl;
  wire[0:0] or_808_nl;
  wire[0:0] nor_419_nl;
  wire[0:0] nor_420_nl;
  wire[0:0] mux_291_nl;
  wire[0:0] nor_421_nl;
  wire[0:0] mux_292_nl;
  wire[0:0] nor_422_nl;
  wire[0:0] nor_409_nl;
  wire[0:0] or_823_nl;
  wire[0:0] nor_410_nl;
  wire[0:0] or_822_nl;
  wire[0:0] nor_411_nl;
  wire[0:0] or_821_nl;
  wire[0:0] nor_412_nl;
  wire[0:0] or_820_nl;
  wire[0:0] nor_413_nl;
  wire[0:0] or_819_nl;
  wire[0:0] nor_414_nl;
  wire[0:0] or_818_nl;
  wire[0:0] nor_415_nl;
  wire[0:0] or_817_nl;
  wire[0:0] nor_416_nl;
  wire[0:0] or_816_nl;
  wire[0:0] mux_301_nl;
  wire[0:0] nor_417_nl;
  wire[0:0] or_815_nl;
  wire[0:0] mux_302_nl;
  wire[0:0] nor_408_nl;
  wire[0:0] and_986_nl;
  wire[0:0] mux_304_nl;
  wire[0:0] nor_407_nl;
  wire[0:0] and_984_nl;
  wire[0:0] and_985_nl;
  wire[0:0] mux_307_nl;
  wire[0:0] nor_406_nl;
  wire[0:0] and_981_nl;
  wire[0:0] and_982_nl;
  wire[0:0] and_983_nl;
  wire[0:0] mux_311_nl;
  wire[0:0] nor_405_nl;
  wire[0:0] and_977_nl;
  wire[0:0] and_978_nl;
  wire[0:0] and_979_nl;
  wire[0:0] and_980_nl;
  wire[0:0] mux_316_nl;
  wire[0:0] nor_404_nl;
  wire[0:0] nor_402_nl;
  wire[0:0] and_973_nl;
  wire[0:0] and_974_nl;
  wire[0:0] and_975_nl;
  wire[0:0] and_976_nl;
  wire[0:0] mux_322_nl;
  wire[0:0] nor_403_nl;
  wire[0:0] nor_399_nl;
  wire[0:0] nor_400_nl;
  wire[0:0] and_969_nl;
  wire[0:0] and_970_nl;
  wire[0:0] and_971_nl;
  wire[0:0] and_972_nl;
  wire[0:0] mux_329_nl;
  wire[0:0] nor_401_nl;
  wire[0:0] nor_395_nl;
  wire[0:0] nor_396_nl;
  wire[0:0] nor_397_nl;
  wire[0:0] and_965_nl;
  wire[0:0] and_966_nl;
  wire[0:0] and_967_nl;
  wire[0:0] and_968_nl;
  wire[0:0] mux_337_nl;
  wire[0:0] nor_398_nl;
  wire[0:0] nor_390_nl;
  wire[0:0] or_919_nl;
  wire[0:0] nor_391_nl;
  wire[0:0] nor_392_nl;
  wire[0:0] nor_393_nl;
  wire[0:0] and_961_nl;
  wire[0:0] and_962_nl;
  wire[0:0] and_963_nl;
  wire[0:0] and_964_nl;
  wire[0:0] mux_346_nl;
  wire[0:0] nor_394_nl;
  wire[0:0] nor_380_nl;
  wire[0:0] or_938_nl;
  wire[0:0] nor_381_nl;
  wire[0:0] or_937_nl;
  wire[0:0] nor_382_nl;
  wire[0:0] or_936_nl;
  wire[0:0] nor_383_nl;
  wire[0:0] or_935_nl;
  wire[0:0] nor_384_nl;
  wire[0:0] or_934_nl;
  wire[0:0] nor_385_nl;
  wire[0:0] or_933_nl;
  wire[0:0] nor_386_nl;
  wire[0:0] or_932_nl;
  wire[0:0] nor_387_nl;
  wire[0:0] or_931_nl;
  wire[0:0] nor_388_nl;
  wire[0:0] or_930_nl;
  wire[0:0] nor_389_nl;
  wire[0:0] or_929_nl;
  wire[0:0] mux_357_nl;
  wire[0:0] nor_379_nl;
  wire[0:0] mux_358_nl;
  wire[0:0] nor_378_nl;
  wire[0:0] mux_359_nl;
  wire[0:0] nor_377_nl;
  wire[0:0] mux_360_nl;
  wire[0:0] nor_376_nl;
  wire[0:0] mux_361_nl;
  wire[0:0] nor_375_nl;
  wire[0:0] mux_362_nl;
  wire[0:0] nor_373_nl;
  wire[0:0] mux_363_nl;
  wire[0:0] nor_374_nl;
  wire[0:0] nor_370_nl;
  wire[0:0] mux_365_nl;
  wire[0:0] nor_371_nl;
  wire[0:0] mux_366_nl;
  wire[0:0] nor_372_nl;
  wire[0:0] nor_366_nl;
  wire[0:0] nor_367_nl;
  wire[0:0] mux_369_nl;
  wire[0:0] nor_368_nl;
  wire[0:0] mux_370_nl;
  wire[0:0] nor_369_nl;
  wire[0:0] nor_361_nl;
  wire[0:0] or_1012_nl;
  wire[0:0] nor_362_nl;
  wire[0:0] nor_363_nl;
  wire[0:0] mux_374_nl;
  wire[0:0] nor_364_nl;
  wire[0:0] mux_375_nl;
  wire[0:0] nor_365_nl;
  wire[0:0] nor_352_nl;
  wire[0:0] or_1027_nl;
  wire[0:0] nor_353_nl;
  wire[0:0] or_1026_nl;
  wire[0:0] nor_354_nl;
  wire[0:0] or_1025_nl;
  wire[0:0] nor_355_nl;
  wire[0:0] or_1024_nl;
  wire[0:0] nor_356_nl;
  wire[0:0] or_1023_nl;
  wire[0:0] nor_357_nl;
  wire[0:0] or_1022_nl;
  wire[0:0] nor_358_nl;
  wire[0:0] or_1021_nl;
  wire[0:0] nor_359_nl;
  wire[0:0] or_1020_nl;
  wire[0:0] mux_384_nl;
  wire[0:0] nor_360_nl;
  wire[0:0] or_1019_nl;
  wire[0:0] mux_385_nl;
  wire[0:0] nor_351_nl;
  wire[0:0] and_960_nl;
  wire[0:0] mux_387_nl;
  wire[0:0] nor_350_nl;
  wire[0:0] and_958_nl;
  wire[0:0] and_959_nl;
  wire[0:0] mux_390_nl;
  wire[0:0] nor_349_nl;
  wire[0:0] and_955_nl;
  wire[0:0] and_956_nl;
  wire[0:0] and_957_nl;
  wire[0:0] mux_394_nl;
  wire[0:0] nor_348_nl;
  wire[0:0] and_951_nl;
  wire[0:0] and_952_nl;
  wire[0:0] and_953_nl;
  wire[0:0] and_954_nl;
  wire[0:0] mux_399_nl;
  wire[0:0] nor_347_nl;
  wire[0:0] nor_345_nl;
  wire[0:0] and_947_nl;
  wire[0:0] and_948_nl;
  wire[0:0] and_949_nl;
  wire[0:0] and_950_nl;
  wire[0:0] mux_405_nl;
  wire[0:0] nor_346_nl;
  wire[0:0] nor_342_nl;
  wire[0:0] nor_343_nl;
  wire[0:0] and_943_nl;
  wire[0:0] and_944_nl;
  wire[0:0] and_945_nl;
  wire[0:0] and_946_nl;
  wire[0:0] mux_412_nl;
  wire[0:0] nor_344_nl;
  wire[0:0] nor_338_nl;
  wire[0:0] nor_339_nl;
  wire[0:0] nor_340_nl;
  wire[0:0] and_939_nl;
  wire[0:0] and_940_nl;
  wire[0:0] and_941_nl;
  wire[0:0] and_942_nl;
  wire[0:0] mux_420_nl;
  wire[0:0] nor_341_nl;
  wire[0:0] nor_333_nl;
  wire[0:0] nand_12_nl;
  wire[0:0] nor_334_nl;
  wire[0:0] nor_335_nl;
  wire[0:0] nor_336_nl;
  wire[0:0] and_935_nl;
  wire[0:0] and_936_nl;
  wire[0:0] and_937_nl;
  wire[0:0] and_938_nl;
  wire[0:0] mux_429_nl;
  wire[0:0] nor_337_nl;
  wire[0:0] nor_324_nl;
  wire[0:0] nand_1_nl;
  wire[0:0] nor_325_nl;
  wire[0:0] nand_2_nl;
  wire[0:0] nor_326_nl;
  wire[0:0] nand_3_nl;
  wire[0:0] nor_327_nl;
  wire[0:0] nand_4_nl;
  wire[0:0] nor_328_nl;
  wire[0:0] nand_5_nl;
  wire[0:0] nor_329_nl;
  wire[0:0] nand_6_nl;
  wire[0:0] nor_330_nl;
  wire[0:0] nand_7_nl;
  wire[0:0] nor_331_nl;
  wire[0:0] nand_8_nl;
  wire[0:0] nor_332_nl;
  wire[0:0] nand_9_nl;
  wire[0:0] and_934_nl;
  wire[0:0] nand_11_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [64:0] nl_rem_13_cmp_a;
  assign nl_rem_13_cmp_a = {{1{rem_13_cmp_a_63_0[63]}}, rem_13_cmp_a_63_0};
  wire [64:0] nl_rem_13_cmp_b;
  assign nl_rem_13_cmp_b = {1'b0 , rem_13_cmp_b_63_0};
  wire [64:0] nl_rem_13_cmp_1_a;
  assign nl_rem_13_cmp_1_a = {{1{rem_13_cmp_1_a_63_0[63]}}, rem_13_cmp_1_a_63_0};
  wire [64:0] nl_rem_13_cmp_1_b;
  assign nl_rem_13_cmp_1_b = {1'b0 , rem_13_cmp_1_b_63_0};
  wire [64:0] nl_rem_13_cmp_2_a;
  assign nl_rem_13_cmp_2_a = {{1{rem_13_cmp_2_a_63_0[63]}}, rem_13_cmp_2_a_63_0};
  wire [64:0] nl_rem_13_cmp_2_b;
  assign nl_rem_13_cmp_2_b = {1'b0 , rem_13_cmp_2_b_63_0};
  wire [64:0] nl_rem_13_cmp_3_a;
  assign nl_rem_13_cmp_3_a = {{1{rem_13_cmp_3_a_63_0[63]}}, rem_13_cmp_3_a_63_0};
  wire [64:0] nl_rem_13_cmp_3_b;
  assign nl_rem_13_cmp_3_b = {1'b0 , rem_13_cmp_3_b_63_0};
  wire [64:0] nl_rem_13_cmp_4_a;
  assign nl_rem_13_cmp_4_a = {{1{rem_13_cmp_4_a_63_0[63]}}, rem_13_cmp_4_a_63_0};
  wire [64:0] nl_rem_13_cmp_4_b;
  assign nl_rem_13_cmp_4_b = {1'b0 , rem_13_cmp_4_b_63_0};
  wire [64:0] nl_rem_13_cmp_5_a;
  assign nl_rem_13_cmp_5_a = {{1{rem_13_cmp_5_a_63_0[63]}}, rem_13_cmp_5_a_63_0};
  wire [64:0] nl_rem_13_cmp_5_b;
  assign nl_rem_13_cmp_5_b = {1'b0 , rem_13_cmp_5_b_63_0};
  wire [64:0] nl_rem_13_cmp_6_a;
  assign nl_rem_13_cmp_6_a = {{1{rem_13_cmp_6_a_63_0[63]}}, rem_13_cmp_6_a_63_0};
  wire [64:0] nl_rem_13_cmp_6_b;
  assign nl_rem_13_cmp_6_b = {1'b0 , rem_13_cmp_6_b_63_0};
  wire [64:0] nl_rem_13_cmp_7_a;
  assign nl_rem_13_cmp_7_a = {{1{rem_13_cmp_7_a_63_0[63]}}, rem_13_cmp_7_a_63_0};
  wire [64:0] nl_rem_13_cmp_7_b;
  assign nl_rem_13_cmp_7_b = {1'b0 , rem_13_cmp_7_b_63_0};
  wire [64:0] nl_rem_13_cmp_8_a;
  assign nl_rem_13_cmp_8_a = {{1{rem_13_cmp_8_a_63_0[63]}}, rem_13_cmp_8_a_63_0};
  wire [64:0] nl_rem_13_cmp_8_b;
  assign nl_rem_13_cmp_8_b = {1'b0 , rem_13_cmp_8_b_63_0};
  wire [64:0] nl_rem_13_cmp_9_a;
  assign nl_rem_13_cmp_9_a = {{1{rem_13_cmp_9_a_63_0[63]}}, rem_13_cmp_9_a_63_0};
  wire [64:0] nl_rem_13_cmp_9_b;
  assign nl_rem_13_cmp_9_b = {1'b0 , rem_13_cmp_9_b_63_0};
  wire [64:0] nl_rem_13_cmp_10_a;
  assign nl_rem_13_cmp_10_a = {{1{rem_13_cmp_10_a_63_0[63]}}, rem_13_cmp_10_a_63_0};
  wire [64:0] nl_rem_13_cmp_10_b;
  assign nl_rem_13_cmp_10_b = {1'b0 , rem_13_cmp_10_b_63_0};
  wire [64:0] nl_rem_13_cmp_11_a;
  assign nl_rem_13_cmp_11_a = {{1{rem_13_cmp_11_a_63_0[63]}}, rem_13_cmp_11_a_63_0};
  wire [64:0] nl_rem_13_cmp_11_b;
  assign nl_rem_13_cmp_11_b = {1'b0 , rem_13_cmp_11_b_63_0};
  ccs_in_v1 #(.rscid(32'sd1),
  .width(32'sd64)) base_rsci (
      .dat(base_rsc_dat),
      .idat(base_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd2),
  .width(32'sd64)) m_rsci (
      .dat(m_rsc_dat),
      .idat(m_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd3),
  .width(32'sd64)) return_rsci (
      .d(return_rsci_d),
      .z(return_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd7),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  mgc_rem #(.width_a(32'sd65),
  .width_b(32'sd65),
  .signd(32'sd1)) rem_13_cmp (
      .a(nl_rem_13_cmp_a[64:0]),
      .b(nl_rem_13_cmp_b[64:0]),
      .z(rem_13_cmp_z)
    );
  mgc_rem #(.width_a(32'sd65),
  .width_b(32'sd65),
  .signd(32'sd1)) rem_13_cmp_1 (
      .a(nl_rem_13_cmp_1_a[64:0]),
      .b(nl_rem_13_cmp_1_b[64:0]),
      .z(rem_13_cmp_1_z)
    );
  mgc_rem #(.width_a(32'sd65),
  .width_b(32'sd65),
  .signd(32'sd1)) rem_13_cmp_2 (
      .a(nl_rem_13_cmp_2_a[64:0]),
      .b(nl_rem_13_cmp_2_b[64:0]),
      .z(rem_13_cmp_2_z)
    );
  mgc_rem #(.width_a(32'sd65),
  .width_b(32'sd65),
  .signd(32'sd1)) rem_13_cmp_3 (
      .a(nl_rem_13_cmp_3_a[64:0]),
      .b(nl_rem_13_cmp_3_b[64:0]),
      .z(rem_13_cmp_3_z)
    );
  mgc_rem #(.width_a(32'sd65),
  .width_b(32'sd65),
  .signd(32'sd1)) rem_13_cmp_4 (
      .a(nl_rem_13_cmp_4_a[64:0]),
      .b(nl_rem_13_cmp_4_b[64:0]),
      .z(rem_13_cmp_4_z)
    );
  mgc_rem #(.width_a(32'sd65),
  .width_b(32'sd65),
  .signd(32'sd1)) rem_13_cmp_5 (
      .a(nl_rem_13_cmp_5_a[64:0]),
      .b(nl_rem_13_cmp_5_b[64:0]),
      .z(rem_13_cmp_5_z)
    );
  mgc_rem #(.width_a(32'sd65),
  .width_b(32'sd65),
  .signd(32'sd1)) rem_13_cmp_6 (
      .a(nl_rem_13_cmp_6_a[64:0]),
      .b(nl_rem_13_cmp_6_b[64:0]),
      .z(rem_13_cmp_6_z)
    );
  mgc_rem #(.width_a(32'sd65),
  .width_b(32'sd65),
  .signd(32'sd1)) rem_13_cmp_7 (
      .a(nl_rem_13_cmp_7_a[64:0]),
      .b(nl_rem_13_cmp_7_b[64:0]),
      .z(rem_13_cmp_7_z)
    );
  mgc_rem #(.width_a(32'sd65),
  .width_b(32'sd65),
  .signd(32'sd1)) rem_13_cmp_8 (
      .a(nl_rem_13_cmp_8_a[64:0]),
      .b(nl_rem_13_cmp_8_b[64:0]),
      .z(rem_13_cmp_8_z)
    );
  mgc_rem #(.width_a(32'sd65),
  .width_b(32'sd65),
  .signd(32'sd1)) rem_13_cmp_9 (
      .a(nl_rem_13_cmp_9_a[64:0]),
      .b(nl_rem_13_cmp_9_b[64:0]),
      .z(rem_13_cmp_9_z)
    );
  mgc_rem #(.width_a(32'sd65),
  .width_b(32'sd65),
  .signd(32'sd1)) rem_13_cmp_10 (
      .a(nl_rem_13_cmp_10_a[64:0]),
      .b(nl_rem_13_cmp_10_b[64:0]),
      .z(rem_13_cmp_10_z)
    );
  mgc_rem #(.width_a(32'sd65),
  .width_b(32'sd65),
  .signd(32'sd1)) rem_13_cmp_11 (
      .a(nl_rem_13_cmp_11_a[64:0]),
      .b(nl_rem_13_cmp_11_b[64:0]),
      .z(rem_13_cmp_11_z)
    );
  assign and_1203_cse = ccs_ccore_en & main_stage_0_12 & asn_itm_11;
  assign and_1173_cse = ccs_ccore_en & (and_dcpl_294 | and_dcpl_300 | and_dcpl_306
      | and_dcpl_312 | and_dcpl_318 | and_dcpl_324 | and_dcpl_330 | and_dcpl_336
      | and_dcpl_342 | and_dcpl_348 | and_tmp_35);
  assign and_1175_cse = ccs_ccore_en & (and_dcpl_356 | and_dcpl_360 | and_dcpl_364
      | and_dcpl_368 | and_dcpl_372 | and_dcpl_376 | and_dcpl_379 | and_dcpl_382
      | and_dcpl_385 | and_dcpl_388 | mux_tmp_76);
  assign and_1177_cse = ccs_ccore_en & (and_dcpl_394 | and_dcpl_397 | and_dcpl_400
      | and_dcpl_403 | and_dcpl_406 | and_dcpl_409 | and_dcpl_413 | and_dcpl_417
      | and_dcpl_421 | and_dcpl_425 | and_tmp_80);
  assign and_1179_cse = ccs_ccore_en & (and_dcpl_431 | and_dcpl_433 | and_dcpl_435
      | and_dcpl_437 | and_dcpl_439 | and_dcpl_442 | and_dcpl_445 | and_dcpl_448
      | and_dcpl_451 | and_dcpl_454 | mux_tmp_141);
  assign and_1181_cse = ccs_ccore_en & (and_dcpl_461 | and_dcpl_465 | and_dcpl_469
      | and_dcpl_473 | and_dcpl_477 | and_dcpl_480 | and_dcpl_483 | and_dcpl_486
      | and_dcpl_489 | and_dcpl_492 | and_tmp_125);
  assign and_1183_cse = ccs_ccore_en & (and_dcpl_498 | and_dcpl_500 | and_dcpl_502
      | and_dcpl_504 | and_dcpl_506 | and_dcpl_508 | and_dcpl_510 | and_dcpl_512
      | and_dcpl_514 | and_dcpl_516 | mux_tmp_206);
  assign and_1185_cse = ccs_ccore_en & (and_dcpl_520 | and_dcpl_523 | and_dcpl_526
      | and_dcpl_529 | and_dcpl_532 | and_dcpl_534 | and_dcpl_536 | and_dcpl_538
      | and_dcpl_540 | and_dcpl_542 | and_tmp_170);
  assign and_1187_cse = ccs_ccore_en & (and_dcpl_546 | and_dcpl_548 | and_dcpl_550
      | and_dcpl_552 | and_dcpl_554 | and_dcpl_556 | and_dcpl_558 | and_dcpl_560
      | and_dcpl_562 | and_dcpl_564 | mux_tmp_271);
  assign and_1189_cse = ccs_ccore_en & (and_dcpl_569 | and_dcpl_573 | and_dcpl_577
      | and_dcpl_581 | and_dcpl_585 | and_dcpl_589 | and_dcpl_593 | and_dcpl_597
      | and_dcpl_601 | and_dcpl_605 | and_tmp_206);
  assign and_1191_cse = ccs_ccore_en & (and_dcpl_610 | and_dcpl_612 | and_dcpl_614
      | and_dcpl_616 | and_dcpl_618 | and_dcpl_622 | and_dcpl_625 | and_dcpl_628
      | and_dcpl_631 | and_dcpl_634 | mux_tmp_354);
  assign and_1193_cse = ccs_ccore_en & (and_dcpl_638 | and_dcpl_641 | and_dcpl_644
      | and_dcpl_647 | and_dcpl_650 | and_dcpl_653 | and_dcpl_657 | and_dcpl_661
      | and_dcpl_665 | and_dcpl_669 | and_tmp_233);
  assign and_1195_cse = ccs_ccore_en & (and_dcpl_673 | and_dcpl_675 | and_dcpl_677
      | and_dcpl_679 | and_dcpl_681 | and_dcpl_684 | and_dcpl_687 | and_dcpl_690
      | and_dcpl_693 | and_dcpl_696 | mux_tmp_437);
  assign and_1205_cse = ccs_ccore_en & and_dcpl_4 & and_dcpl_2;
  assign and_1207_cse = ccs_ccore_en & and_dcpl_4 & and_dcpl_6;
  assign and_1209_cse = ccs_ccore_en & and_dcpl_4 & and_dcpl_9;
  assign and_1211_cse = ccs_ccore_en & and_dcpl_4 & and_dcpl_11;
  assign and_1213_cse = ccs_ccore_en & and_dcpl_13 & and_dcpl_2;
  assign and_1215_cse = ccs_ccore_en & and_dcpl_13 & and_dcpl_6;
  assign and_1217_cse = ccs_ccore_en & and_dcpl_13 & and_dcpl_9;
  assign and_1219_cse = ccs_ccore_en & and_dcpl_13 & and_dcpl_11;
  assign and_1221_cse = ccs_ccore_en & and_dcpl_4 & and_dcpl_18 & (~ (rem_12cyc_st_10_1_0[0]));
  assign and_1223_cse = ccs_ccore_en & and_dcpl_4 & and_dcpl_18 & (rem_12cyc_st_10_1_0[0]);
  assign and_1225_cse = ccs_ccore_en & and_dcpl_4 & and_dcpl_23 & (~ (rem_12cyc_st_10_1_0[0]));
  assign and_1227_cse = ccs_ccore_en & and_dcpl_4 & and_dcpl_23 & (rem_12cyc_st_10_1_0[0]);
  assign and_1229_cse = ccs_ccore_en & and_dcpl_3;
  assign and_1231_cse = ccs_ccore_en & and_dcpl_31 & and_dcpl_29;
  assign and_1233_cse = ccs_ccore_en & and_dcpl_31 & and_dcpl_33;
  assign and_1235_cse = ccs_ccore_en & and_dcpl_31 & and_dcpl_36;
  assign and_1237_cse = ccs_ccore_en & and_dcpl_31 & and_dcpl_38;
  assign and_1239_cse = ccs_ccore_en & and_dcpl_40 & and_dcpl_29;
  assign and_1241_cse = ccs_ccore_en & and_dcpl_40 & and_dcpl_33;
  assign and_1243_cse = ccs_ccore_en & and_dcpl_40 & and_dcpl_36;
  assign and_1245_cse = ccs_ccore_en & and_dcpl_40 & and_dcpl_38;
  assign and_1247_cse = ccs_ccore_en & and_dcpl_31 & and_dcpl_45 & (~ (rem_12cyc_st_9_1_0[0]));
  assign and_1249_cse = ccs_ccore_en & and_dcpl_31 & and_dcpl_45 & (rem_12cyc_st_9_1_0[0]);
  assign and_1251_cse = ccs_ccore_en & and_dcpl_31 & and_dcpl_50 & (~ (rem_12cyc_st_9_1_0[0]));
  assign and_1253_cse = ccs_ccore_en & and_dcpl_31 & and_dcpl_50 & (rem_12cyc_st_9_1_0[0]);
  assign and_1255_cse = ccs_ccore_en & and_dcpl_30;
  assign and_1257_cse = ccs_ccore_en & and_dcpl_58 & and_dcpl_56;
  assign and_1259_cse = ccs_ccore_en & and_dcpl_58 & and_dcpl_60;
  assign and_1261_cse = ccs_ccore_en & and_dcpl_58 & and_dcpl_63;
  assign and_1263_cse = ccs_ccore_en & and_dcpl_58 & and_dcpl_65;
  assign and_1265_cse = ccs_ccore_en & and_dcpl_67 & and_dcpl_56;
  assign and_1267_cse = ccs_ccore_en & and_dcpl_67 & and_dcpl_60;
  assign and_1269_cse = ccs_ccore_en & and_dcpl_67 & and_dcpl_63;
  assign and_1271_cse = ccs_ccore_en & and_dcpl_67 & and_dcpl_65;
  assign and_1273_cse = ccs_ccore_en & and_dcpl_58 & and_dcpl_72 & (~ (rem_12cyc_st_8_1_0[0]));
  assign and_1275_cse = ccs_ccore_en & and_dcpl_58 & and_dcpl_72 & (rem_12cyc_st_8_1_0[0]);
  assign and_1277_cse = ccs_ccore_en & and_dcpl_58 & and_dcpl_77 & (~ (rem_12cyc_st_8_1_0[0]));
  assign and_1279_cse = ccs_ccore_en & and_dcpl_58 & and_dcpl_77 & (rem_12cyc_st_8_1_0[0]);
  assign and_1281_cse = ccs_ccore_en & and_dcpl_57;
  assign and_1283_cse = ccs_ccore_en & and_dcpl_85 & and_dcpl_83;
  assign and_1285_cse = ccs_ccore_en & and_dcpl_85 & and_dcpl_87;
  assign and_1287_cse = ccs_ccore_en & and_dcpl_85 & and_dcpl_90;
  assign and_1289_cse = ccs_ccore_en & and_dcpl_85 & and_dcpl_92;
  assign and_1291_cse = ccs_ccore_en & and_dcpl_94 & and_dcpl_83;
  assign and_1293_cse = ccs_ccore_en & and_dcpl_94 & and_dcpl_87;
  assign and_1295_cse = ccs_ccore_en & and_dcpl_94 & and_dcpl_90;
  assign and_1297_cse = ccs_ccore_en & and_dcpl_94 & and_dcpl_92;
  assign and_1299_cse = ccs_ccore_en & and_dcpl_85 & and_dcpl_99 & (~ (rem_12cyc_st_7_1_0[0]));
  assign and_1301_cse = ccs_ccore_en & and_dcpl_85 & and_dcpl_99 & (rem_12cyc_st_7_1_0[0]);
  assign and_1303_cse = ccs_ccore_en & and_dcpl_85 & and_dcpl_104 & (~ (rem_12cyc_st_7_1_0[0]));
  assign and_1305_cse = ccs_ccore_en & and_dcpl_85 & and_dcpl_104 & (rem_12cyc_st_7_1_0[0]);
  assign and_1307_cse = ccs_ccore_en & and_dcpl_84;
  assign and_1309_cse = ccs_ccore_en & and_dcpl_112 & and_dcpl_110;
  assign and_1311_cse = ccs_ccore_en & and_dcpl_112 & and_dcpl_115;
  assign and_1313_cse = ccs_ccore_en & and_dcpl_112 & and_dcpl_117;
  assign and_1315_cse = ccs_ccore_en & and_dcpl_112 & and_dcpl_119;
  assign and_1317_cse = ccs_ccore_en & and_dcpl_121 & and_dcpl_110;
  assign and_1319_cse = ccs_ccore_en & and_dcpl_121 & and_dcpl_115;
  assign and_1321_cse = ccs_ccore_en & and_dcpl_121 & and_dcpl_117;
  assign and_1323_cse = ccs_ccore_en & and_dcpl_121 & and_dcpl_119;
  assign and_1325_cse = ccs_ccore_en & and_dcpl_112 & and_dcpl_126 & (~ (rem_12cyc_st_6_1_0[1]));
  assign and_1327_cse = ccs_ccore_en & and_dcpl_112 & and_dcpl_129 & (~ (rem_12cyc_st_6_1_0[1]));
  assign and_1329_cse = ccs_ccore_en & and_dcpl_112 & and_dcpl_126 & (rem_12cyc_st_6_1_0[1]);
  assign and_1331_cse = ccs_ccore_en & and_dcpl_112 & and_dcpl_129 & (rem_12cyc_st_6_1_0[1]);
  assign and_1333_cse = ccs_ccore_en & and_dcpl_111;
  assign and_1335_cse = ccs_ccore_en & and_dcpl_139 & and_dcpl_137;
  assign and_1337_cse = ccs_ccore_en & and_dcpl_139 & and_dcpl_141;
  assign and_1339_cse = ccs_ccore_en & and_dcpl_139 & and_dcpl_144;
  assign and_1341_cse = ccs_ccore_en & and_dcpl_139 & and_dcpl_146;
  assign and_1343_cse = ccs_ccore_en & and_dcpl_148 & and_dcpl_137;
  assign and_1345_cse = ccs_ccore_en & and_dcpl_148 & and_dcpl_141;
  assign and_1347_cse = ccs_ccore_en & and_dcpl_148 & and_dcpl_144;
  assign and_1349_cse = ccs_ccore_en & and_dcpl_148 & and_dcpl_146;
  assign and_1351_cse = ccs_ccore_en & and_dcpl_139 & and_dcpl_153 & (~ (rem_12cyc_st_5_1_0[0]));
  assign and_1353_cse = ccs_ccore_en & and_dcpl_139 & and_dcpl_153 & (rem_12cyc_st_5_1_0[0]);
  assign and_1355_cse = ccs_ccore_en & and_dcpl_139 & and_dcpl_158 & (~ (rem_12cyc_st_5_1_0[0]));
  assign and_1357_cse = ccs_ccore_en & and_dcpl_139 & and_dcpl_158 & (rem_12cyc_st_5_1_0[0]);
  assign and_1359_cse = ccs_ccore_en & and_dcpl_138;
  assign and_1361_cse = ccs_ccore_en & and_dcpl_166 & and_dcpl_164;
  assign and_1363_cse = ccs_ccore_en & and_dcpl_166 & and_dcpl_168;
  assign and_1365_cse = ccs_ccore_en & and_dcpl_166 & and_dcpl_171;
  assign and_1367_cse = ccs_ccore_en & and_dcpl_166 & and_dcpl_173;
  assign and_1369_cse = ccs_ccore_en & and_dcpl_166 & and_dcpl_175 & (~ (rem_12cyc_st_4_1_0[0]));
  assign and_1371_cse = ccs_ccore_en & and_dcpl_166 & and_dcpl_175 & (rem_12cyc_st_4_1_0[0]);
  assign and_1373_cse = ccs_ccore_en & and_dcpl_166 & and_dcpl_180 & (~ (rem_12cyc_st_4_1_0[0]));
  assign and_1375_cse = ccs_ccore_en & and_dcpl_166 & and_dcpl_180 & (rem_12cyc_st_4_1_0[0]);
  assign and_1377_cse = ccs_ccore_en & and_dcpl_185 & and_dcpl_164;
  assign and_1379_cse = ccs_ccore_en & and_dcpl_185 & and_dcpl_168;
  assign and_1381_cse = ccs_ccore_en & and_dcpl_185 & and_dcpl_171;
  assign and_1383_cse = ccs_ccore_en & and_dcpl_185 & and_dcpl_173;
  assign and_1385_cse = ccs_ccore_en & and_dcpl_165;
  assign and_1387_cse = ccs_ccore_en & and_dcpl_193 & and_dcpl_191;
  assign and_1389_cse = ccs_ccore_en & and_dcpl_193 & and_dcpl_195;
  assign and_1391_cse = ccs_ccore_en & and_dcpl_193 & and_dcpl_198;
  assign and_1393_cse = ccs_ccore_en & and_dcpl_193 & and_dcpl_200;
  assign and_1395_cse = ccs_ccore_en & and_dcpl_202 & and_dcpl_191;
  assign and_1397_cse = ccs_ccore_en & and_dcpl_202 & and_dcpl_195;
  assign and_1399_cse = ccs_ccore_en & and_dcpl_202 & and_dcpl_198;
  assign and_1401_cse = ccs_ccore_en & and_dcpl_202 & and_dcpl_200;
  assign and_1403_cse = ccs_ccore_en & and_dcpl_193 & and_dcpl_207 & (~ (rem_12cyc_st_3_1_0[0]));
  assign and_1405_cse = ccs_ccore_en & and_dcpl_193 & and_dcpl_207 & (rem_12cyc_st_3_1_0[0]);
  assign and_1407_cse = ccs_ccore_en & and_dcpl_193 & and_dcpl_212 & (~ (rem_12cyc_st_3_1_0[0]));
  assign and_1409_cse = ccs_ccore_en & and_dcpl_193 & and_dcpl_212 & (rem_12cyc_st_3_1_0[0]);
  assign and_1411_cse = ccs_ccore_en & and_dcpl_192;
  assign and_1413_cse = ccs_ccore_en & and_dcpl_220 & and_dcpl_218;
  assign and_1415_cse = ccs_ccore_en & and_dcpl_220 & and_dcpl_222;
  assign and_1417_cse = ccs_ccore_en & and_dcpl_220 & and_dcpl_225;
  assign and_1419_cse = ccs_ccore_en & and_dcpl_220 & and_dcpl_227;
  assign and_1421_cse = ccs_ccore_en & and_dcpl_220 & and_dcpl_229 & (~ (rem_12cyc_st_2_1_0[0]));
  assign and_1423_cse = ccs_ccore_en & and_dcpl_220 & and_dcpl_229 & (rem_12cyc_st_2_1_0[0]);
  assign and_1425_cse = ccs_ccore_en & and_dcpl_220 & and_dcpl_234 & (~ (rem_12cyc_st_2_1_0[0]));
  assign and_1427_cse = ccs_ccore_en & and_dcpl_220 & and_dcpl_234 & (rem_12cyc_st_2_1_0[0]);
  assign and_1429_cse = ccs_ccore_en & and_dcpl_239 & and_dcpl_218;
  assign and_1431_cse = ccs_ccore_en & and_dcpl_239 & and_dcpl_222;
  assign and_1433_cse = ccs_ccore_en & and_dcpl_239 & and_dcpl_225;
  assign and_1435_cse = ccs_ccore_en & and_dcpl_239 & and_dcpl_227;
  assign and_1437_cse = ccs_ccore_en & and_dcpl_219;
  assign and_1439_cse = ccs_ccore_en & and_dcpl_247 & and_dcpl_245;
  assign and_1441_cse = ccs_ccore_en & and_dcpl_247 & and_dcpl_249;
  assign and_1443_cse = ccs_ccore_en & and_dcpl_247 & and_dcpl_252;
  assign and_1445_cse = ccs_ccore_en & and_dcpl_247 & and_dcpl_254;
  assign and_1447_cse = ccs_ccore_en & and_dcpl_256 & and_dcpl_245;
  assign and_1449_cse = ccs_ccore_en & and_dcpl_256 & and_dcpl_249;
  assign and_1451_cse = ccs_ccore_en & and_dcpl_256 & and_dcpl_252;
  assign and_1453_cse = ccs_ccore_en & and_dcpl_256 & and_dcpl_254;
  assign and_1455_cse = ccs_ccore_en & and_dcpl_247 & and_dcpl_261 & (~ (rem_12cyc_1_0[0]));
  assign and_1457_cse = ccs_ccore_en & and_dcpl_247 & and_dcpl_261 & (rem_12cyc_1_0[0]);
  assign and_1459_cse = ccs_ccore_en & and_dcpl_247 & and_dcpl_266 & (~ (rem_12cyc_1_0[0]));
  assign and_1461_cse = ccs_ccore_en & and_dcpl_247 & and_dcpl_266 & (rem_12cyc_1_0[0]);
  assign and_1463_cse = ccs_ccore_en & and_dcpl_246;
  assign and_1197_cse = ccs_ccore_en & ccs_ccore_start_rsci_idat;
  assign and_273_nl = and_dcpl_272 & and_dcpl_271;
  assign and_275_nl = and_dcpl_272 & and_dcpl_274;
  assign and_277_nl = and_dcpl_272 & and_dcpl_276;
  assign and_279_nl = and_dcpl_272 & and_dcpl_278;
  assign and_281_nl = and_dcpl_280 & and_dcpl_271;
  assign and_282_nl = and_dcpl_280 & and_dcpl_274;
  assign and_283_nl = and_dcpl_280 & and_dcpl_276;
  assign and_284_nl = and_dcpl_280 & and_dcpl_278;
  assign and_286_nl = and_dcpl_285 & and_dcpl_271;
  assign and_287_nl = and_dcpl_285 & and_dcpl_274;
  assign and_288_nl = and_dcpl_285 & and_dcpl_276;
  assign and_289_nl = and_dcpl_285 & and_dcpl_278;
  assign and_290_nl = (rem_12cyc_st_12_3_2==2'b11);
  assign result_sva_duc_mx0 = MUX1HOT_v_64_13_2((rem_13_cmp_1_z[63:0]), (rem_13_cmp_2_z[63:0]),
      (rem_13_cmp_3_z[63:0]), (rem_13_cmp_4_z[63:0]), (rem_13_cmp_5_z[63:0]), (rem_13_cmp_6_z[63:0]),
      (rem_13_cmp_7_z[63:0]), (rem_13_cmp_8_z[63:0]), (rem_13_cmp_9_z[63:0]), (rem_13_cmp_10_z[63:0]),
      (rem_13_cmp_11_z[63:0]), (rem_13_cmp_z[63:0]), result_sva_duc, {and_273_nl
      , and_275_nl , and_277_nl , and_279_nl , and_281_nl , and_282_nl , and_283_nl
      , and_284_nl , and_286_nl , and_287_nl , and_288_nl , and_289_nl , and_290_nl});
  assign nl_acc_1_tmp = ({rem_12cyc_3_2 , rem_12cyc_1_0}) + 4'b0001;
  assign acc_1_tmp = nl_acc_1_tmp[3:0];
  assign xor_nl = (acc_1_tmp[2]) ^ (acc_1_tmp[3]);
  assign nor_nl = ~((acc_1_tmp[3:2]!=2'b10));
  assign nl_acc_tmp = conv_u2u_1_2(xor_nl) + conv_u2u_1_2(nor_nl);
  assign acc_tmp = nl_acc_tmp[1:0];
  assign and_dcpl_1 = ~((rem_12cyc_st_10_3_2[1]) | (rem_12cyc_st_10_1_0[1]));
  assign and_dcpl_2 = and_dcpl_1 & (~ (rem_12cyc_st_10_1_0[0]));
  assign and_dcpl_3 = main_stage_0_11 & asn_itm_10;
  assign and_dcpl_4 = and_dcpl_3 & (~ (rem_12cyc_st_10_3_2[0]));
  assign and_dcpl_6 = and_dcpl_1 & (rem_12cyc_st_10_1_0[0]);
  assign and_dcpl_8 = (~ (rem_12cyc_st_10_3_2[1])) & (rem_12cyc_st_10_1_0[1]);
  assign and_dcpl_9 = and_dcpl_8 & (~ (rem_12cyc_st_10_1_0[0]));
  assign and_dcpl_11 = and_dcpl_8 & (rem_12cyc_st_10_1_0[0]);
  assign and_dcpl_13 = and_dcpl_3 & (rem_12cyc_st_10_3_2[0]);
  assign and_dcpl_18 = (rem_12cyc_st_10_3_2[1]) & (~ (rem_12cyc_st_10_1_0[1]));
  assign and_dcpl_23 = (rem_12cyc_st_10_3_2[1]) & (rem_12cyc_st_10_1_0[1]);
  assign and_dcpl_28 = ~((rem_12cyc_st_9_3_2[1]) | (rem_12cyc_st_9_1_0[1]));
  assign and_dcpl_29 = and_dcpl_28 & (~ (rem_12cyc_st_9_1_0[0]));
  assign and_dcpl_30 = main_stage_0_10 & asn_itm_9;
  assign and_dcpl_31 = and_dcpl_30 & (~ (rem_12cyc_st_9_3_2[0]));
  assign and_dcpl_33 = and_dcpl_28 & (rem_12cyc_st_9_1_0[0]);
  assign and_dcpl_35 = (~ (rem_12cyc_st_9_3_2[1])) & (rem_12cyc_st_9_1_0[1]);
  assign and_dcpl_36 = and_dcpl_35 & (~ (rem_12cyc_st_9_1_0[0]));
  assign and_dcpl_38 = and_dcpl_35 & (rem_12cyc_st_9_1_0[0]);
  assign and_dcpl_40 = and_dcpl_30 & (rem_12cyc_st_9_3_2[0]);
  assign and_dcpl_45 = (rem_12cyc_st_9_3_2[1]) & (~ (rem_12cyc_st_9_1_0[1]));
  assign and_dcpl_50 = (rem_12cyc_st_9_3_2[1]) & (rem_12cyc_st_9_1_0[1]);
  assign and_dcpl_55 = ~((rem_12cyc_st_8_3_2[1]) | (rem_12cyc_st_8_1_0[1]));
  assign and_dcpl_56 = and_dcpl_55 & (~ (rem_12cyc_st_8_1_0[0]));
  assign and_dcpl_57 = main_stage_0_9 & asn_itm_8;
  assign and_dcpl_58 = and_dcpl_57 & (~ (rem_12cyc_st_8_3_2[0]));
  assign and_dcpl_60 = and_dcpl_55 & (rem_12cyc_st_8_1_0[0]);
  assign and_dcpl_62 = (~ (rem_12cyc_st_8_3_2[1])) & (rem_12cyc_st_8_1_0[1]);
  assign and_dcpl_63 = and_dcpl_62 & (~ (rem_12cyc_st_8_1_0[0]));
  assign and_dcpl_65 = and_dcpl_62 & (rem_12cyc_st_8_1_0[0]);
  assign and_dcpl_67 = and_dcpl_57 & (rem_12cyc_st_8_3_2[0]);
  assign and_dcpl_72 = (rem_12cyc_st_8_3_2[1]) & (~ (rem_12cyc_st_8_1_0[1]));
  assign and_dcpl_77 = (rem_12cyc_st_8_3_2[1]) & (rem_12cyc_st_8_1_0[1]);
  assign and_dcpl_82 = ~((rem_12cyc_st_7_3_2[1]) | (rem_12cyc_st_7_1_0[1]));
  assign and_dcpl_83 = and_dcpl_82 & (~ (rem_12cyc_st_7_1_0[0]));
  assign and_dcpl_84 = main_stage_0_8 & asn_itm_7;
  assign and_dcpl_85 = and_dcpl_84 & (~ (rem_12cyc_st_7_3_2[0]));
  assign and_dcpl_87 = and_dcpl_82 & (rem_12cyc_st_7_1_0[0]);
  assign and_dcpl_89 = (~ (rem_12cyc_st_7_3_2[1])) & (rem_12cyc_st_7_1_0[1]);
  assign and_dcpl_90 = and_dcpl_89 & (~ (rem_12cyc_st_7_1_0[0]));
  assign and_dcpl_92 = and_dcpl_89 & (rem_12cyc_st_7_1_0[0]);
  assign and_dcpl_94 = and_dcpl_84 & (rem_12cyc_st_7_3_2[0]);
  assign and_dcpl_99 = (rem_12cyc_st_7_3_2[1]) & (~ (rem_12cyc_st_7_1_0[1]));
  assign and_dcpl_104 = (rem_12cyc_st_7_3_2[1]) & (rem_12cyc_st_7_1_0[1]);
  assign and_dcpl_109 = ~((rem_12cyc_st_6_3_2[1]) | (rem_12cyc_st_6_1_0[0]));
  assign and_dcpl_110 = and_dcpl_109 & (~ (rem_12cyc_st_6_1_0[1]));
  assign and_dcpl_111 = main_stage_0_7 & asn_itm_6;
  assign and_dcpl_112 = and_dcpl_111 & (~ (rem_12cyc_st_6_3_2[0]));
  assign and_dcpl_114 = (~ (rem_12cyc_st_6_3_2[1])) & (rem_12cyc_st_6_1_0[0]);
  assign and_dcpl_115 = and_dcpl_114 & (~ (rem_12cyc_st_6_1_0[1]));
  assign and_dcpl_117 = and_dcpl_109 & (rem_12cyc_st_6_1_0[1]);
  assign and_dcpl_119 = and_dcpl_114 & (rem_12cyc_st_6_1_0[1]);
  assign and_dcpl_121 = and_dcpl_111 & (rem_12cyc_st_6_3_2[0]);
  assign and_dcpl_126 = (rem_12cyc_st_6_3_2[1]) & (~ (rem_12cyc_st_6_1_0[0]));
  assign and_dcpl_129 = (rem_12cyc_st_6_3_2[1]) & (rem_12cyc_st_6_1_0[0]);
  assign and_dcpl_136 = ~((rem_12cyc_st_5_3_2[1]) | (rem_12cyc_st_5_1_0[1]));
  assign and_dcpl_137 = and_dcpl_136 & (~ (rem_12cyc_st_5_1_0[0]));
  assign and_dcpl_138 = main_stage_0_6 & asn_itm_5;
  assign and_dcpl_139 = and_dcpl_138 & (~ (rem_12cyc_st_5_3_2[0]));
  assign and_dcpl_141 = and_dcpl_136 & (rem_12cyc_st_5_1_0[0]);
  assign and_dcpl_143 = (~ (rem_12cyc_st_5_3_2[1])) & (rem_12cyc_st_5_1_0[1]);
  assign and_dcpl_144 = and_dcpl_143 & (~ (rem_12cyc_st_5_1_0[0]));
  assign and_dcpl_146 = and_dcpl_143 & (rem_12cyc_st_5_1_0[0]);
  assign and_dcpl_148 = and_dcpl_138 & (rem_12cyc_st_5_3_2[0]);
  assign and_dcpl_153 = (rem_12cyc_st_5_3_2[1]) & (~ (rem_12cyc_st_5_1_0[1]));
  assign and_dcpl_158 = (rem_12cyc_st_5_3_2[1]) & (rem_12cyc_st_5_1_0[1]);
  assign and_dcpl_163 = ~((rem_12cyc_st_4_3_2[0]) | (rem_12cyc_st_4_1_0[1]));
  assign and_dcpl_164 = and_dcpl_163 & (~ (rem_12cyc_st_4_1_0[0]));
  assign and_dcpl_165 = main_stage_0_5 & asn_itm_4;
  assign and_dcpl_166 = and_dcpl_165 & (~ (rem_12cyc_st_4_3_2[1]));
  assign and_dcpl_168 = and_dcpl_163 & (rem_12cyc_st_4_1_0[0]);
  assign and_dcpl_170 = (~ (rem_12cyc_st_4_3_2[0])) & (rem_12cyc_st_4_1_0[1]);
  assign and_dcpl_171 = and_dcpl_170 & (~ (rem_12cyc_st_4_1_0[0]));
  assign and_dcpl_173 = and_dcpl_170 & (rem_12cyc_st_4_1_0[0]);
  assign and_dcpl_175 = (rem_12cyc_st_4_3_2[0]) & (~ (rem_12cyc_st_4_1_0[1]));
  assign and_dcpl_180 = (rem_12cyc_st_4_3_2[0]) & (rem_12cyc_st_4_1_0[1]);
  assign and_dcpl_185 = and_dcpl_165 & (rem_12cyc_st_4_3_2[1]);
  assign and_dcpl_190 = ~((rem_12cyc_st_3_3_2[1]) | (rem_12cyc_st_3_1_0[1]));
  assign and_dcpl_191 = and_dcpl_190 & (~ (rem_12cyc_st_3_1_0[0]));
  assign and_dcpl_192 = main_stage_0_4 & asn_itm_3;
  assign and_dcpl_193 = and_dcpl_192 & (~ (rem_12cyc_st_3_3_2[0]));
  assign and_dcpl_195 = and_dcpl_190 & (rem_12cyc_st_3_1_0[0]);
  assign and_dcpl_197 = (~ (rem_12cyc_st_3_3_2[1])) & (rem_12cyc_st_3_1_0[1]);
  assign and_dcpl_198 = and_dcpl_197 & (~ (rem_12cyc_st_3_1_0[0]));
  assign and_dcpl_200 = and_dcpl_197 & (rem_12cyc_st_3_1_0[0]);
  assign and_dcpl_202 = and_dcpl_192 & (rem_12cyc_st_3_3_2[0]);
  assign and_dcpl_207 = (rem_12cyc_st_3_3_2[1]) & (~ (rem_12cyc_st_3_1_0[1]));
  assign and_dcpl_212 = (rem_12cyc_st_3_3_2[1]) & (rem_12cyc_st_3_1_0[1]);
  assign and_dcpl_217 = ~((rem_12cyc_st_2_3_2[0]) | (rem_12cyc_st_2_1_0[1]));
  assign and_dcpl_218 = and_dcpl_217 & (~ (rem_12cyc_st_2_1_0[0]));
  assign and_dcpl_219 = main_stage_0_3 & asn_itm_2;
  assign and_dcpl_220 = and_dcpl_219 & (~ (rem_12cyc_st_2_3_2[1]));
  assign and_dcpl_222 = and_dcpl_217 & (rem_12cyc_st_2_1_0[0]);
  assign and_dcpl_224 = (~ (rem_12cyc_st_2_3_2[0])) & (rem_12cyc_st_2_1_0[1]);
  assign and_dcpl_225 = and_dcpl_224 & (~ (rem_12cyc_st_2_1_0[0]));
  assign and_dcpl_227 = and_dcpl_224 & (rem_12cyc_st_2_1_0[0]);
  assign and_dcpl_229 = (rem_12cyc_st_2_3_2[0]) & (~ (rem_12cyc_st_2_1_0[1]));
  assign and_dcpl_234 = (rem_12cyc_st_2_3_2[0]) & (rem_12cyc_st_2_1_0[1]);
  assign and_dcpl_239 = and_dcpl_219 & (rem_12cyc_st_2_3_2[1]);
  assign and_dcpl_244 = ~((rem_12cyc_3_2[1]) | (rem_12cyc_1_0[1]));
  assign and_dcpl_245 = and_dcpl_244 & (~ (rem_12cyc_1_0[0]));
  assign and_dcpl_246 = main_stage_0_2 & asn_itm_1;
  assign and_dcpl_247 = and_dcpl_246 & (~ (rem_12cyc_3_2[0]));
  assign and_dcpl_249 = and_dcpl_244 & (rem_12cyc_1_0[0]);
  assign and_dcpl_251 = (~ (rem_12cyc_3_2[1])) & (rem_12cyc_1_0[1]);
  assign and_dcpl_252 = and_dcpl_251 & (~ (rem_12cyc_1_0[0]));
  assign and_dcpl_254 = and_dcpl_251 & (rem_12cyc_1_0[0]);
  assign and_dcpl_256 = and_dcpl_246 & (rem_12cyc_3_2[0]);
  assign and_dcpl_261 = (rem_12cyc_3_2[1]) & (~ (rem_12cyc_1_0[1]));
  assign and_dcpl_266 = (rem_12cyc_3_2[1]) & (rem_12cyc_1_0[1]);
  assign and_dcpl_271 = ~((rem_12cyc_st_12_1_0!=2'b00));
  assign and_dcpl_272 = ~((rem_12cyc_st_12_3_2!=2'b00));
  assign and_dcpl_274 = (rem_12cyc_st_12_1_0==2'b01);
  assign and_dcpl_276 = (rem_12cyc_st_12_1_0==2'b10);
  assign and_dcpl_278 = (rem_12cyc_st_12_1_0==2'b11);
  assign and_dcpl_280 = (rem_12cyc_st_12_3_2==2'b01);
  assign and_dcpl_285 = (rem_12cyc_st_12_3_2==2'b10);
  assign and_dcpl_291 = ~((acc_1_tmp[1:0]!=2'b00));
  assign and_dcpl_292 = ccs_ccore_start_rsci_idat & (~ (acc_tmp[0]));
  assign and_dcpl_293 = and_dcpl_292 & (~ (acc_tmp[1]));
  assign and_dcpl_294 = and_dcpl_293 & and_dcpl_291;
  assign and_dcpl_295 = ~((rem_12cyc_st_2_3_2!=2'b00));
  assign and_dcpl_296 = and_dcpl_295 & (~ (rem_12cyc_st_2_1_0[1]));
  assign and_dcpl_298 = (~ (rem_12cyc_st_2_1_0[0])) & main_stage_0_3 & asn_itm_2;
  assign not_tmp_54 = ~(asn_itm_1 & main_stage_0_2);
  assign or_tmp_2 = (rem_12cyc_1_0!=2'b00) | (rem_12cyc_3_2!=2'b00) | not_tmp_54;
  assign or_1_cse = (acc_1_tmp[1:0]!=2'b00) | (acc_tmp!=2'b00);
  assign nor_518_nl = ~(ccs_ccore_start_rsci_idat | (~ or_tmp_2));
  assign mux_14_nl = MUX_s_1_2_2(nor_518_nl, or_tmp_2, or_1_cse);
  assign and_dcpl_300 = mux_14_nl & and_dcpl_298 & and_dcpl_296;
  assign and_dcpl_301 = ~((rem_12cyc_st_3_3_2!=2'b00));
  assign and_dcpl_302 = and_dcpl_301 & (~ (rem_12cyc_st_3_1_0[1]));
  assign and_dcpl_304 = (~ (rem_12cyc_st_3_1_0[0])) & main_stage_0_4 & asn_itm_3;
  assign or_6_cse = (rem_12cyc_st_2_1_0[1]) | (rem_12cyc_st_2_3_2!=2'b00) | (~ asn_itm_2)
      | (~ main_stage_0_3) | (rem_12cyc_st_2_1_0[0]);
  assign and_tmp = or_6_cse & or_tmp_2;
  assign nor_517_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp));
  assign mux_15_nl = MUX_s_1_2_2(nor_517_nl, and_tmp, or_1_cse);
  assign and_dcpl_306 = mux_15_nl & and_dcpl_304 & and_dcpl_302;
  assign and_dcpl_307 = ~((rem_12cyc_st_4_3_2!=2'b00));
  assign and_dcpl_308 = and_dcpl_307 & (~ (rem_12cyc_st_4_1_0[1]));
  assign and_dcpl_310 = (~ (rem_12cyc_st_4_1_0[0])) & main_stage_0_5 & asn_itm_4;
  assign or_10_cse = (rem_12cyc_st_3_1_0[1]) | (rem_12cyc_st_3_3_2!=2'b00) | (~ asn_itm_3)
      | (~ main_stage_0_4) | (rem_12cyc_st_3_1_0[0]);
  assign and_tmp_2 = or_6_cse & or_10_cse & or_tmp_2;
  assign nor_516_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_2));
  assign mux_16_nl = MUX_s_1_2_2(nor_516_nl, and_tmp_2, or_1_cse);
  assign and_dcpl_312 = mux_16_nl & and_dcpl_310 & and_dcpl_308;
  assign and_dcpl_313 = ~((rem_12cyc_st_5_3_2!=2'b00));
  assign and_dcpl_314 = and_dcpl_313 & (~ (rem_12cyc_st_5_1_0[1]));
  assign and_dcpl_316 = (~ (rem_12cyc_st_5_1_0[0])) & main_stage_0_6 & asn_itm_5;
  assign or_15_cse = (rem_12cyc_st_4_1_0[1]) | (rem_12cyc_st_4_3_2!=2'b00) | (~ asn_itm_4)
      | (~ main_stage_0_5) | (rem_12cyc_st_4_1_0[0]);
  assign and_tmp_5 = or_6_cse & or_10_cse & or_15_cse & or_tmp_2;
  assign nor_515_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_5));
  assign mux_17_nl = MUX_s_1_2_2(nor_515_nl, and_tmp_5, or_1_cse);
  assign and_dcpl_318 = mux_17_nl & and_dcpl_316 & and_dcpl_314;
  assign or_21_cse = (rem_12cyc_st_5_1_0[1]) | (rem_12cyc_st_5_3_2!=2'b00) | (~ asn_itm_5)
      | (~ main_stage_0_6) | (rem_12cyc_st_5_1_0[0]);
  assign and_tmp_9 = or_6_cse & or_10_cse & or_15_cse & or_21_cse & or_tmp_2;
  assign nor_514_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_9));
  assign mux_18_nl = MUX_s_1_2_2(nor_514_nl, and_tmp_9, or_1_cse);
  assign and_dcpl_324 = mux_18_nl & and_dcpl_112 & and_dcpl_110;
  assign or_28_cse = (rem_12cyc_st_6_1_0!=2'b00) | (rem_12cyc_st_6_3_2!=2'b00);
  assign nor_512_nl = ~(and_dcpl_111 | (~ or_tmp_2));
  assign mux_19_nl = MUX_s_1_2_2(nor_512_nl, or_tmp_2, or_28_cse);
  assign and_tmp_13 = or_6_cse & or_10_cse & or_15_cse & or_21_cse & mux_19_nl;
  assign nor_513_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_13));
  assign mux_20_nl = MUX_s_1_2_2(nor_513_nl, and_tmp_13, or_1_cse);
  assign and_dcpl_330 = mux_20_nl & and_dcpl_85 & and_dcpl_83;
  assign or_37_cse = (rem_12cyc_st_7_1_0!=2'b00) | (rem_12cyc_st_7_3_2!=2'b00);
  assign nor_509_nl = ~(and_dcpl_84 | (~ or_tmp_2));
  assign mux_tmp_19 = MUX_s_1_2_2(nor_509_nl, or_tmp_2, or_37_cse);
  assign nor_510_nl = ~(and_dcpl_111 | (~ mux_tmp_19));
  assign mux_22_nl = MUX_s_1_2_2(nor_510_nl, mux_tmp_19, or_28_cse);
  assign and_tmp_17 = or_6_cse & or_10_cse & or_15_cse & or_21_cse & mux_22_nl;
  assign nor_511_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_17));
  assign mux_23_nl = MUX_s_1_2_2(nor_511_nl, and_tmp_17, or_1_cse);
  assign and_dcpl_336 = mux_23_nl & and_dcpl_58 & and_dcpl_56;
  assign or_48_cse = (rem_12cyc_st_8_1_0!=2'b00) | (rem_12cyc_st_8_3_2!=2'b00);
  assign nor_505_nl = ~(and_dcpl_57 | (~ or_tmp_2));
  assign mux_tmp_22 = MUX_s_1_2_2(nor_505_nl, or_tmp_2, or_48_cse);
  assign nor_506_nl = ~(and_dcpl_84 | (~ mux_tmp_22));
  assign mux_tmp_23 = MUX_s_1_2_2(nor_506_nl, mux_tmp_22, or_37_cse);
  assign nor_507_nl = ~(and_dcpl_111 | (~ mux_tmp_23));
  assign mux_26_nl = MUX_s_1_2_2(nor_507_nl, mux_tmp_23, or_28_cse);
  assign and_tmp_21 = or_6_cse & or_10_cse & or_15_cse & or_21_cse & mux_26_nl;
  assign nor_508_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_21));
  assign mux_27_nl = MUX_s_1_2_2(nor_508_nl, and_tmp_21, or_1_cse);
  assign and_dcpl_342 = mux_27_nl & and_dcpl_31 & and_dcpl_29;
  assign nor_500_nl = ~(and_dcpl_30 | (~ or_tmp_2));
  assign or_61_nl = (rem_12cyc_st_9_1_0!=2'b00) | (rem_12cyc_st_9_3_2!=2'b00);
  assign mux_tmp_26 = MUX_s_1_2_2(nor_500_nl, or_tmp_2, or_61_nl);
  assign nor_501_nl = ~(and_dcpl_57 | (~ mux_tmp_26));
  assign mux_tmp_27 = MUX_s_1_2_2(nor_501_nl, mux_tmp_26, or_48_cse);
  assign nor_502_nl = ~(and_dcpl_84 | (~ mux_tmp_27));
  assign mux_tmp_28 = MUX_s_1_2_2(nor_502_nl, mux_tmp_27, or_37_cse);
  assign nor_503_nl = ~(and_dcpl_111 | (~ mux_tmp_28));
  assign mux_31_nl = MUX_s_1_2_2(nor_503_nl, mux_tmp_28, or_28_cse);
  assign and_tmp_25 = or_6_cse & or_10_cse & or_15_cse & or_21_cse & mux_31_nl;
  assign nor_504_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_25));
  assign mux_32_nl = MUX_s_1_2_2(nor_504_nl, and_tmp_25, or_1_cse);
  assign and_dcpl_348 = mux_32_nl & and_dcpl_4 & and_dcpl_2;
  assign and_tmp_35 = ((~ main_stage_0_2) | (~ asn_itm_1) | (rem_12cyc_3_2!=2'b00)
      | (rem_12cyc_1_0!=2'b00)) & ((~ main_stage_0_8) | (~ asn_itm_7) | (rem_12cyc_st_7_1_0!=2'b00)
      | (rem_12cyc_st_7_3_2!=2'b00)) & ((~ main_stage_0_9) | (~ asn_itm_8) | (rem_12cyc_st_8_1_0!=2'b00)
      | (rem_12cyc_st_8_3_2!=2'b00)) & ((~ main_stage_0_10) | (~ asn_itm_9) | (rem_12cyc_st_9_1_0!=2'b00)
      | (rem_12cyc_st_9_3_2!=2'b00)) & or_6_cse & or_10_cse & or_15_cse & or_21_cse
      & ((~ main_stage_0_7) | (~ asn_itm_6) | (rem_12cyc_st_6_1_0!=2'b00) | (rem_12cyc_st_6_3_2!=2'b00))
      & ((~ main_stage_0_11) | (~ asn_itm_10) | (rem_12cyc_st_10_1_0!=2'b00) | (rem_12cyc_st_10_3_2!=2'b00))
      & ((acc_tmp!=2'b00) | (acc_1_tmp[1:0]!=2'b00) | (~ ccs_ccore_start_rsci_idat));
  assign and_dcpl_355 = (acc_1_tmp[1:0]==2'b01);
  assign and_dcpl_356 = and_dcpl_293 & and_dcpl_355;
  assign and_dcpl_358 = (rem_12cyc_st_2_1_0[0]) & main_stage_0_3 & asn_itm_2;
  assign or_tmp_80 = (rem_12cyc_1_0!=2'b01) | (rem_12cyc_3_2!=2'b00) | not_tmp_54;
  assign or_83_cse = (acc_1_tmp[1:0]!=2'b01) | (acc_tmp!=2'b00);
  assign nor_499_nl = ~(ccs_ccore_start_rsci_idat | (~ or_tmp_80));
  assign mux_33_nl = MUX_s_1_2_2(nor_499_nl, or_tmp_80, or_83_cse);
  assign and_dcpl_360 = mux_33_nl & and_dcpl_358 & and_dcpl_296;
  assign and_dcpl_362 = (rem_12cyc_st_3_1_0[0]) & main_stage_0_4 & asn_itm_3;
  assign nand_276_cse = ~(asn_itm_2 & main_stage_0_3 & (rem_12cyc_st_2_1_0[0]));
  assign or_88_cse = (rem_12cyc_st_2_1_0[1]) | (rem_12cyc_st_2_3_2!=2'b00);
  assign and_1168_nl = nand_276_cse & or_tmp_80;
  assign mux_tmp_32 = MUX_s_1_2_2(and_1168_nl, or_tmp_80, or_88_cse);
  assign nor_498_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_32));
  assign mux_35_nl = MUX_s_1_2_2(nor_498_nl, mux_tmp_32, or_83_cse);
  assign and_dcpl_364 = mux_35_nl & and_dcpl_362 & and_dcpl_302;
  assign and_dcpl_366 = (rem_12cyc_st_4_1_0[0]) & main_stage_0_5 & asn_itm_4;
  assign nand_274_cse = ~(asn_itm_3 & main_stage_0_4 & (rem_12cyc_st_3_1_0[0]));
  assign or_93_cse = (rem_12cyc_st_3_1_0[1]) | (rem_12cyc_st_3_3_2!=2'b00);
  assign and_1166_nl = nand_274_cse & or_tmp_80;
  assign mux_tmp_34 = MUX_s_1_2_2(and_1166_nl, or_tmp_80, or_93_cse);
  assign and_1167_nl = nand_276_cse & mux_tmp_34;
  assign mux_tmp_35 = MUX_s_1_2_2(and_1167_nl, mux_tmp_34, or_88_cse);
  assign nor_497_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_35));
  assign mux_38_nl = MUX_s_1_2_2(nor_497_nl, mux_tmp_35, or_83_cse);
  assign and_dcpl_368 = mux_38_nl & and_dcpl_366 & and_dcpl_308;
  assign and_dcpl_370 = (rem_12cyc_st_5_1_0[0]) & main_stage_0_6 & asn_itm_5;
  assign nand_271_cse = ~(asn_itm_4 & main_stage_0_5 & (rem_12cyc_st_4_1_0[0]));
  assign or_100_cse = (rem_12cyc_st_4_1_0[1]) | (rem_12cyc_st_4_3_2!=2'b00);
  assign and_1163_nl = nand_271_cse & or_tmp_80;
  assign mux_tmp_37 = MUX_s_1_2_2(and_1163_nl, or_tmp_80, or_100_cse);
  assign and_1164_nl = nand_274_cse & mux_tmp_37;
  assign mux_tmp_38 = MUX_s_1_2_2(and_1164_nl, mux_tmp_37, or_93_cse);
  assign and_1165_nl = nand_276_cse & mux_tmp_38;
  assign mux_tmp_39 = MUX_s_1_2_2(and_1165_nl, mux_tmp_38, or_88_cse);
  assign nor_496_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_39));
  assign mux_42_nl = MUX_s_1_2_2(nor_496_nl, mux_tmp_39, or_83_cse);
  assign and_dcpl_372 = mux_42_nl & and_dcpl_370 & and_dcpl_314;
  assign nand_267_cse = ~(asn_itm_5 & main_stage_0_6 & (rem_12cyc_st_5_1_0[0]));
  assign or_109_cse = (rem_12cyc_st_5_1_0[1]) | (rem_12cyc_st_5_3_2!=2'b00);
  assign and_1159_nl = nand_267_cse & or_tmp_80;
  assign mux_tmp_41 = MUX_s_1_2_2(and_1159_nl, or_tmp_80, or_109_cse);
  assign and_1160_nl = nand_271_cse & mux_tmp_41;
  assign mux_tmp_42 = MUX_s_1_2_2(and_1160_nl, mux_tmp_41, or_100_cse);
  assign and_1161_nl = nand_274_cse & mux_tmp_42;
  assign mux_tmp_43 = MUX_s_1_2_2(and_1161_nl, mux_tmp_42, or_93_cse);
  assign and_1162_nl = nand_276_cse & mux_tmp_43;
  assign mux_tmp_44 = MUX_s_1_2_2(and_1162_nl, mux_tmp_43, or_88_cse);
  assign nor_495_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_44));
  assign mux_47_nl = MUX_s_1_2_2(nor_495_nl, mux_tmp_44, or_83_cse);
  assign and_dcpl_376 = mux_47_nl & and_dcpl_112 & and_dcpl_115;
  assign or_120_cse = (rem_12cyc_st_6_1_0!=2'b01) | (rem_12cyc_st_6_3_2!=2'b00);
  assign nor_493_nl = ~(and_dcpl_111 | (~ or_tmp_80));
  assign mux_tmp_46 = MUX_s_1_2_2(nor_493_nl, or_tmp_80, or_120_cse);
  assign and_1155_nl = nand_267_cse & mux_tmp_46;
  assign mux_tmp_47 = MUX_s_1_2_2(and_1155_nl, mux_tmp_46, or_109_cse);
  assign and_1156_nl = nand_271_cse & mux_tmp_47;
  assign mux_tmp_48 = MUX_s_1_2_2(and_1156_nl, mux_tmp_47, or_100_cse);
  assign and_1157_nl = nand_274_cse & mux_tmp_48;
  assign mux_tmp_49 = MUX_s_1_2_2(and_1157_nl, mux_tmp_48, or_93_cse);
  assign and_1158_nl = nand_276_cse & mux_tmp_49;
  assign mux_tmp_50 = MUX_s_1_2_2(and_1158_nl, mux_tmp_49, or_88_cse);
  assign nor_494_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_50));
  assign mux_53_nl = MUX_s_1_2_2(nor_494_nl, mux_tmp_50, or_83_cse);
  assign and_dcpl_379 = mux_53_nl & and_dcpl_85 & and_dcpl_87;
  assign or_133_cse = (rem_12cyc_st_7_1_0!=2'b01) | (rem_12cyc_st_7_3_2!=2'b00);
  assign nor_490_nl = ~(and_dcpl_84 | (~ or_tmp_80));
  assign mux_tmp_52 = MUX_s_1_2_2(nor_490_nl, or_tmp_80, or_133_cse);
  assign nor_491_nl = ~(and_dcpl_111 | (~ mux_tmp_52));
  assign mux_tmp_53 = MUX_s_1_2_2(nor_491_nl, mux_tmp_52, or_120_cse);
  assign and_1151_nl = nand_267_cse & mux_tmp_53;
  assign mux_tmp_54 = MUX_s_1_2_2(and_1151_nl, mux_tmp_53, or_109_cse);
  assign and_1152_nl = nand_271_cse & mux_tmp_54;
  assign mux_tmp_55 = MUX_s_1_2_2(and_1152_nl, mux_tmp_54, or_100_cse);
  assign and_1153_nl = nand_274_cse & mux_tmp_55;
  assign mux_tmp_56 = MUX_s_1_2_2(and_1153_nl, mux_tmp_55, or_93_cse);
  assign and_1154_nl = nand_276_cse & mux_tmp_56;
  assign mux_tmp_57 = MUX_s_1_2_2(and_1154_nl, mux_tmp_56, or_88_cse);
  assign nor_492_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_57));
  assign mux_60_nl = MUX_s_1_2_2(nor_492_nl, mux_tmp_57, or_83_cse);
  assign and_dcpl_382 = mux_60_nl & and_dcpl_58 & and_dcpl_60;
  assign or_148_cse = (rem_12cyc_st_8_1_0!=2'b01) | (rem_12cyc_st_8_3_2!=2'b00);
  assign nor_486_nl = ~(and_dcpl_57 | (~ or_tmp_80));
  assign mux_tmp_59 = MUX_s_1_2_2(nor_486_nl, or_tmp_80, or_148_cse);
  assign nor_487_nl = ~(and_dcpl_84 | (~ mux_tmp_59));
  assign mux_tmp_60 = MUX_s_1_2_2(nor_487_nl, mux_tmp_59, or_133_cse);
  assign nor_488_nl = ~(and_dcpl_111 | (~ mux_tmp_60));
  assign mux_tmp_61 = MUX_s_1_2_2(nor_488_nl, mux_tmp_60, or_120_cse);
  assign and_1147_nl = nand_267_cse & mux_tmp_61;
  assign mux_tmp_62 = MUX_s_1_2_2(and_1147_nl, mux_tmp_61, or_109_cse);
  assign and_1148_nl = nand_271_cse & mux_tmp_62;
  assign mux_tmp_63 = MUX_s_1_2_2(and_1148_nl, mux_tmp_62, or_100_cse);
  assign and_1149_nl = nand_274_cse & mux_tmp_63;
  assign mux_tmp_64 = MUX_s_1_2_2(and_1149_nl, mux_tmp_63, or_93_cse);
  assign and_1150_nl = nand_276_cse & mux_tmp_64;
  assign mux_tmp_65 = MUX_s_1_2_2(and_1150_nl, mux_tmp_64, or_88_cse);
  assign nor_489_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_65));
  assign mux_68_nl = MUX_s_1_2_2(nor_489_nl, mux_tmp_65, or_83_cse);
  assign and_dcpl_385 = mux_68_nl & and_dcpl_31 & and_dcpl_33;
  assign nor_481_nl = ~(and_dcpl_30 | (~ or_tmp_80));
  assign or_165_nl = (rem_12cyc_st_9_1_0!=2'b01) | (rem_12cyc_st_9_3_2!=2'b00);
  assign mux_tmp_67 = MUX_s_1_2_2(nor_481_nl, or_tmp_80, or_165_nl);
  assign nor_482_nl = ~(and_dcpl_57 | (~ mux_tmp_67));
  assign mux_tmp_68 = MUX_s_1_2_2(nor_482_nl, mux_tmp_67, or_148_cse);
  assign nor_483_nl = ~(and_dcpl_84 | (~ mux_tmp_68));
  assign mux_tmp_69 = MUX_s_1_2_2(nor_483_nl, mux_tmp_68, or_133_cse);
  assign nor_484_nl = ~(and_dcpl_111 | (~ mux_tmp_69));
  assign mux_tmp_70 = MUX_s_1_2_2(nor_484_nl, mux_tmp_69, or_120_cse);
  assign and_1143_nl = nand_267_cse & mux_tmp_70;
  assign mux_tmp_71 = MUX_s_1_2_2(and_1143_nl, mux_tmp_70, or_109_cse);
  assign and_1144_nl = nand_271_cse & mux_tmp_71;
  assign mux_tmp_72 = MUX_s_1_2_2(and_1144_nl, mux_tmp_71, or_100_cse);
  assign and_1145_nl = nand_274_cse & mux_tmp_72;
  assign mux_tmp_73 = MUX_s_1_2_2(and_1145_nl, mux_tmp_72, or_93_cse);
  assign and_1146_nl = nand_276_cse & mux_tmp_73;
  assign mux_tmp_74 = MUX_s_1_2_2(and_1146_nl, mux_tmp_73, or_88_cse);
  assign nor_485_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_74));
  assign mux_77_nl = MUX_s_1_2_2(nor_485_nl, mux_tmp_74, or_83_cse);
  assign and_dcpl_388 = mux_77_nl & and_dcpl_4 & and_dcpl_6;
  assign nand_250_cse = ~((acc_1_tmp[0]) & ccs_ccore_start_rsci_idat);
  assign and_tmp_44 = ((~ main_stage_0_8) | (~ asn_itm_7) | (rem_12cyc_st_7_1_0!=2'b01)
      | (rem_12cyc_st_7_3_2!=2'b00)) & ((~ main_stage_0_9) | (~ asn_itm_8) | (rem_12cyc_st_8_1_0!=2'b01)
      | (rem_12cyc_st_8_3_2!=2'b00)) & ((~ main_stage_0_10) | (~ asn_itm_9) | (rem_12cyc_st_9_1_0!=2'b01)
      | (rem_12cyc_st_9_3_2!=2'b00)) & ((~ main_stage_0_3) | (~ asn_itm_2) | (rem_12cyc_st_2_1_0!=2'b01)
      | (rem_12cyc_st_2_3_2!=2'b00)) & ((~ main_stage_0_4) | (~ asn_itm_3) | (rem_12cyc_st_3_1_0!=2'b01)
      | (rem_12cyc_st_3_3_2!=2'b00)) & ((~ main_stage_0_5) | (~ asn_itm_4) | (rem_12cyc_st_4_1_0!=2'b01)
      | (rem_12cyc_st_4_3_2!=2'b00)) & ((~ main_stage_0_6) | (~ asn_itm_5) | (rem_12cyc_st_5_1_0!=2'b01)
      | (rem_12cyc_st_5_3_2!=2'b00)) & ((~ main_stage_0_7) | (~ asn_itm_6) | (rem_12cyc_st_6_1_0!=2'b01)
      | (rem_12cyc_st_6_3_2!=2'b00)) & ((~ main_stage_0_11) | (~ asn_itm_10) | (rem_12cyc_st_10_1_0!=2'b01)
      | (rem_12cyc_st_10_3_2!=2'b00)) & ((acc_tmp!=2'b00) | (acc_1_tmp[1]) | nand_250_cse);
  assign nor_480_nl = ~((rem_12cyc_1_0[0]) | (~ and_tmp_44));
  assign or_175_nl = (~ main_stage_0_2) | (~ asn_itm_1) | (rem_12cyc_3_2!=2'b00)
      | (rem_12cyc_1_0[1]);
  assign mux_tmp_76 = MUX_s_1_2_2(nor_480_nl, and_tmp_44, or_175_nl);
  assign and_dcpl_393 = (acc_1_tmp[1:0]==2'b10);
  assign and_dcpl_394 = and_dcpl_293 & and_dcpl_393;
  assign and_dcpl_395 = and_dcpl_295 & (rem_12cyc_st_2_1_0[1]);
  assign or_tmp_185 = (rem_12cyc_1_0!=2'b10) | (rem_12cyc_3_2!=2'b00) | not_tmp_54;
  assign or_190_cse = (acc_1_tmp[1:0]!=2'b10) | (acc_tmp!=2'b00);
  assign nor_479_nl = ~(ccs_ccore_start_rsci_idat | (~ or_tmp_185));
  assign mux_79_nl = MUX_s_1_2_2(nor_479_nl, or_tmp_185, or_190_cse);
  assign and_dcpl_397 = mux_79_nl & and_dcpl_298 & and_dcpl_395;
  assign and_dcpl_398 = and_dcpl_301 & (rem_12cyc_st_3_1_0[1]);
  assign or_195_cse = (~ (rem_12cyc_st_2_1_0[1])) | (rem_12cyc_st_2_3_2!=2'b00) |
      (~ asn_itm_2) | (~ main_stage_0_3) | (rem_12cyc_st_2_1_0[0]);
  assign and_tmp_45 = or_195_cse & or_tmp_185;
  assign nor_478_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_45));
  assign mux_80_nl = MUX_s_1_2_2(nor_478_nl, and_tmp_45, or_190_cse);
  assign and_dcpl_400 = mux_80_nl & and_dcpl_304 & and_dcpl_398;
  assign and_dcpl_401 = and_dcpl_307 & (rem_12cyc_st_4_1_0[1]);
  assign or_199_cse = (~ (rem_12cyc_st_3_1_0[1])) | (rem_12cyc_st_3_3_2!=2'b00) |
      (~ asn_itm_3) | (~ main_stage_0_4) | (rem_12cyc_st_3_1_0[0]);
  assign and_tmp_47 = or_195_cse & or_199_cse & or_tmp_185;
  assign nor_477_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_47));
  assign mux_81_nl = MUX_s_1_2_2(nor_477_nl, and_tmp_47, or_190_cse);
  assign and_dcpl_403 = mux_81_nl & and_dcpl_310 & and_dcpl_401;
  assign and_dcpl_404 = and_dcpl_313 & (rem_12cyc_st_5_1_0[1]);
  assign or_204_cse = (~ (rem_12cyc_st_4_1_0[1])) | (rem_12cyc_st_4_3_2!=2'b00) |
      (~ asn_itm_4) | (~ main_stage_0_5) | (rem_12cyc_st_4_1_0[0]);
  assign and_tmp_50 = or_195_cse & or_199_cse & or_204_cse & or_tmp_185;
  assign nor_476_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_50));
  assign mux_82_nl = MUX_s_1_2_2(nor_476_nl, and_tmp_50, or_190_cse);
  assign and_dcpl_406 = mux_82_nl & and_dcpl_316 & and_dcpl_404;
  assign or_210_cse = (~ (rem_12cyc_st_5_1_0[1])) | (rem_12cyc_st_5_3_2!=2'b00) |
      (~ asn_itm_5) | (~ main_stage_0_6) | (rem_12cyc_st_5_1_0[0]);
  assign and_tmp_54 = or_195_cse & or_199_cse & or_204_cse & or_210_cse & or_tmp_185;
  assign nor_475_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_54));
  assign mux_83_nl = MUX_s_1_2_2(nor_475_nl, and_tmp_54, or_190_cse);
  assign and_dcpl_409 = mux_83_nl & and_dcpl_112 & and_dcpl_117;
  assign or_217_cse = (rem_12cyc_st_6_1_0!=2'b10) | (rem_12cyc_st_6_3_2!=2'b00);
  assign nor_473_nl = ~(and_dcpl_111 | (~ or_tmp_185));
  assign mux_84_nl = MUX_s_1_2_2(nor_473_nl, or_tmp_185, or_217_cse);
  assign and_tmp_58 = or_195_cse & or_199_cse & or_204_cse & or_210_cse & mux_84_nl;
  assign nor_474_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_58));
  assign mux_85_nl = MUX_s_1_2_2(nor_474_nl, and_tmp_58, or_190_cse);
  assign and_dcpl_413 = mux_85_nl & and_dcpl_85 & and_dcpl_90;
  assign or_226_cse = (rem_12cyc_st_7_1_0!=2'b10) | (rem_12cyc_st_7_3_2!=2'b00);
  assign nor_470_nl = ~(and_dcpl_84 | (~ or_tmp_185));
  assign mux_tmp_84 = MUX_s_1_2_2(nor_470_nl, or_tmp_185, or_226_cse);
  assign nor_471_nl = ~(and_dcpl_111 | (~ mux_tmp_84));
  assign mux_87_nl = MUX_s_1_2_2(nor_471_nl, mux_tmp_84, or_217_cse);
  assign and_tmp_62 = or_195_cse & or_199_cse & or_204_cse & or_210_cse & mux_87_nl;
  assign nor_472_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_62));
  assign mux_88_nl = MUX_s_1_2_2(nor_472_nl, and_tmp_62, or_190_cse);
  assign and_dcpl_417 = mux_88_nl & and_dcpl_58 & and_dcpl_63;
  assign or_237_cse = (rem_12cyc_st_8_1_0!=2'b10) | (rem_12cyc_st_8_3_2!=2'b00);
  assign nor_466_nl = ~(and_dcpl_57 | (~ or_tmp_185));
  assign mux_tmp_87 = MUX_s_1_2_2(nor_466_nl, or_tmp_185, or_237_cse);
  assign nor_467_nl = ~(and_dcpl_84 | (~ mux_tmp_87));
  assign mux_tmp_88 = MUX_s_1_2_2(nor_467_nl, mux_tmp_87, or_226_cse);
  assign nor_468_nl = ~(and_dcpl_111 | (~ mux_tmp_88));
  assign mux_91_nl = MUX_s_1_2_2(nor_468_nl, mux_tmp_88, or_217_cse);
  assign and_tmp_66 = or_195_cse & or_199_cse & or_204_cse & or_210_cse & mux_91_nl;
  assign nor_469_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_66));
  assign mux_92_nl = MUX_s_1_2_2(nor_469_nl, and_tmp_66, or_190_cse);
  assign and_dcpl_421 = mux_92_nl & and_dcpl_31 & and_dcpl_36;
  assign nor_461_nl = ~(and_dcpl_30 | (~ or_tmp_185));
  assign or_250_nl = (rem_12cyc_st_9_1_0!=2'b10) | (rem_12cyc_st_9_3_2!=2'b00);
  assign mux_tmp_91 = MUX_s_1_2_2(nor_461_nl, or_tmp_185, or_250_nl);
  assign nor_462_nl = ~(and_dcpl_57 | (~ mux_tmp_91));
  assign mux_tmp_92 = MUX_s_1_2_2(nor_462_nl, mux_tmp_91, or_237_cse);
  assign nor_463_nl = ~(and_dcpl_84 | (~ mux_tmp_92));
  assign mux_tmp_93 = MUX_s_1_2_2(nor_463_nl, mux_tmp_92, or_226_cse);
  assign nor_464_nl = ~(and_dcpl_111 | (~ mux_tmp_93));
  assign mux_96_nl = MUX_s_1_2_2(nor_464_nl, mux_tmp_93, or_217_cse);
  assign and_tmp_70 = or_195_cse & or_199_cse & or_204_cse & or_210_cse & mux_96_nl;
  assign nor_465_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_70));
  assign mux_97_nl = MUX_s_1_2_2(nor_465_nl, and_tmp_70, or_190_cse);
  assign and_dcpl_425 = mux_97_nl & and_dcpl_4 & and_dcpl_9;
  assign and_tmp_80 = ((~ main_stage_0_2) | (~ asn_itm_1) | (rem_12cyc_3_2!=2'b00)
      | (rem_12cyc_1_0!=2'b10)) & ((~ main_stage_0_8) | (~ asn_itm_7) | (rem_12cyc_st_7_1_0!=2'b10)
      | (rem_12cyc_st_7_3_2!=2'b00)) & ((~ main_stage_0_9) | (~ asn_itm_8) | (rem_12cyc_st_8_1_0!=2'b10)
      | (rem_12cyc_st_8_3_2!=2'b00)) & ((~ main_stage_0_10) | (~ asn_itm_9) | (rem_12cyc_st_9_1_0!=2'b10)
      | (rem_12cyc_st_9_3_2!=2'b00)) & or_195_cse & or_199_cse & or_204_cse & or_210_cse
      & ((~ main_stage_0_7) | (~ asn_itm_6) | (rem_12cyc_st_6_1_0!=2'b10) | (rem_12cyc_st_6_3_2!=2'b00))
      & ((~ main_stage_0_11) | (~ asn_itm_10) | (rem_12cyc_st_10_1_0!=2'b10) | (rem_12cyc_st_10_3_2!=2'b00))
      & ((acc_tmp!=2'b00) | (acc_1_tmp[1:0]!=2'b10) | (~ ccs_ccore_start_rsci_idat));
  assign and_dcpl_430 = (acc_1_tmp[1:0]==2'b11);
  assign and_dcpl_431 = and_dcpl_293 & and_dcpl_430;
  assign or_tmp_263 = (rem_12cyc_1_0!=2'b11) | (rem_12cyc_3_2!=2'b00) | not_tmp_54;
  assign or_270_cse = (acc_1_tmp[1:0]!=2'b11) | (acc_tmp!=2'b00);
  assign nor_460_nl = ~(ccs_ccore_start_rsci_idat | (~ or_tmp_263));
  assign mux_98_nl = MUX_s_1_2_2(nor_460_nl, or_tmp_263, or_270_cse);
  assign and_dcpl_433 = mux_98_nl & and_dcpl_358 & and_dcpl_395;
  assign or_275_cse = (~ (rem_12cyc_st_2_1_0[1])) | (rem_12cyc_st_2_3_2!=2'b00);
  assign and_1142_nl = nand_276_cse & or_tmp_263;
  assign mux_tmp_97 = MUX_s_1_2_2(and_1142_nl, or_tmp_263, or_275_cse);
  assign nor_459_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_97));
  assign mux_100_nl = MUX_s_1_2_2(nor_459_nl, mux_tmp_97, or_270_cse);
  assign and_dcpl_435 = mux_100_nl & and_dcpl_362 & and_dcpl_398;
  assign or_280_cse = (~ (rem_12cyc_st_3_1_0[1])) | (rem_12cyc_st_3_3_2!=2'b00);
  assign and_1140_nl = nand_274_cse & or_tmp_263;
  assign mux_tmp_99 = MUX_s_1_2_2(and_1140_nl, or_tmp_263, or_280_cse);
  assign and_1141_nl = nand_276_cse & mux_tmp_99;
  assign mux_tmp_100 = MUX_s_1_2_2(and_1141_nl, mux_tmp_99, or_275_cse);
  assign nor_458_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_100));
  assign mux_103_nl = MUX_s_1_2_2(nor_458_nl, mux_tmp_100, or_270_cse);
  assign and_dcpl_437 = mux_103_nl & and_dcpl_366 & and_dcpl_401;
  assign or_287_cse = (~ (rem_12cyc_st_4_1_0[1])) | (rem_12cyc_st_4_3_2!=2'b00);
  assign and_1137_nl = nand_271_cse & or_tmp_263;
  assign mux_tmp_102 = MUX_s_1_2_2(and_1137_nl, or_tmp_263, or_287_cse);
  assign and_1138_nl = nand_274_cse & mux_tmp_102;
  assign mux_tmp_103 = MUX_s_1_2_2(and_1138_nl, mux_tmp_102, or_280_cse);
  assign and_1139_nl = nand_276_cse & mux_tmp_103;
  assign mux_tmp_104 = MUX_s_1_2_2(and_1139_nl, mux_tmp_103, or_275_cse);
  assign nor_457_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_104));
  assign mux_107_nl = MUX_s_1_2_2(nor_457_nl, mux_tmp_104, or_270_cse);
  assign and_dcpl_439 = mux_107_nl & and_dcpl_370 & and_dcpl_404;
  assign or_296_cse = (~ (rem_12cyc_st_5_1_0[1])) | (rem_12cyc_st_5_3_2!=2'b00);
  assign and_1133_nl = nand_267_cse & or_tmp_263;
  assign mux_tmp_106 = MUX_s_1_2_2(and_1133_nl, or_tmp_263, or_296_cse);
  assign and_1134_nl = nand_271_cse & mux_tmp_106;
  assign mux_tmp_107 = MUX_s_1_2_2(and_1134_nl, mux_tmp_106, or_287_cse);
  assign and_1135_nl = nand_274_cse & mux_tmp_107;
  assign mux_tmp_108 = MUX_s_1_2_2(and_1135_nl, mux_tmp_107, or_280_cse);
  assign and_1136_nl = nand_276_cse & mux_tmp_108;
  assign mux_tmp_109 = MUX_s_1_2_2(and_1136_nl, mux_tmp_108, or_275_cse);
  assign nor_456_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_109));
  assign mux_112_nl = MUX_s_1_2_2(nor_456_nl, mux_tmp_109, or_270_cse);
  assign and_dcpl_442 = mux_112_nl & and_dcpl_112 & and_dcpl_119;
  assign or_307_cse = (rem_12cyc_st_6_1_0!=2'b11) | (rem_12cyc_st_6_3_2!=2'b00);
  assign nor_454_nl = ~(and_dcpl_111 | (~ or_tmp_263));
  assign mux_tmp_111 = MUX_s_1_2_2(nor_454_nl, or_tmp_263, or_307_cse);
  assign and_1129_nl = nand_267_cse & mux_tmp_111;
  assign mux_tmp_112 = MUX_s_1_2_2(and_1129_nl, mux_tmp_111, or_296_cse);
  assign and_1130_nl = nand_271_cse & mux_tmp_112;
  assign mux_tmp_113 = MUX_s_1_2_2(and_1130_nl, mux_tmp_112, or_287_cse);
  assign and_1131_nl = nand_274_cse & mux_tmp_113;
  assign mux_tmp_114 = MUX_s_1_2_2(and_1131_nl, mux_tmp_113, or_280_cse);
  assign and_1132_nl = nand_276_cse & mux_tmp_114;
  assign mux_tmp_115 = MUX_s_1_2_2(and_1132_nl, mux_tmp_114, or_275_cse);
  assign nor_455_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_115));
  assign mux_118_nl = MUX_s_1_2_2(nor_455_nl, mux_tmp_115, or_270_cse);
  assign and_dcpl_445 = mux_118_nl & and_dcpl_85 & and_dcpl_92;
  assign or_320_cse = (rem_12cyc_st_7_1_0!=2'b11) | (rem_12cyc_st_7_3_2!=2'b00);
  assign nor_451_nl = ~(and_dcpl_84 | (~ or_tmp_263));
  assign mux_tmp_117 = MUX_s_1_2_2(nor_451_nl, or_tmp_263, or_320_cse);
  assign nor_452_nl = ~(and_dcpl_111 | (~ mux_tmp_117));
  assign mux_tmp_118 = MUX_s_1_2_2(nor_452_nl, mux_tmp_117, or_307_cse);
  assign and_1125_nl = nand_267_cse & mux_tmp_118;
  assign mux_tmp_119 = MUX_s_1_2_2(and_1125_nl, mux_tmp_118, or_296_cse);
  assign and_1126_nl = nand_271_cse & mux_tmp_119;
  assign mux_tmp_120 = MUX_s_1_2_2(and_1126_nl, mux_tmp_119, or_287_cse);
  assign and_1127_nl = nand_274_cse & mux_tmp_120;
  assign mux_tmp_121 = MUX_s_1_2_2(and_1127_nl, mux_tmp_120, or_280_cse);
  assign and_1128_nl = nand_276_cse & mux_tmp_121;
  assign mux_tmp_122 = MUX_s_1_2_2(and_1128_nl, mux_tmp_121, or_275_cse);
  assign nor_453_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_122));
  assign mux_125_nl = MUX_s_1_2_2(nor_453_nl, mux_tmp_122, or_270_cse);
  assign and_dcpl_448 = mux_125_nl & and_dcpl_58 & and_dcpl_65;
  assign or_335_cse = (rem_12cyc_st_8_1_0!=2'b11) | (rem_12cyc_st_8_3_2!=2'b00);
  assign nor_447_nl = ~(and_dcpl_57 | (~ or_tmp_263));
  assign mux_tmp_124 = MUX_s_1_2_2(nor_447_nl, or_tmp_263, or_335_cse);
  assign nor_448_nl = ~(and_dcpl_84 | (~ mux_tmp_124));
  assign mux_tmp_125 = MUX_s_1_2_2(nor_448_nl, mux_tmp_124, or_320_cse);
  assign nor_449_nl = ~(and_dcpl_111 | (~ mux_tmp_125));
  assign mux_tmp_126 = MUX_s_1_2_2(nor_449_nl, mux_tmp_125, or_307_cse);
  assign and_1121_nl = nand_267_cse & mux_tmp_126;
  assign mux_tmp_127 = MUX_s_1_2_2(and_1121_nl, mux_tmp_126, or_296_cse);
  assign and_1122_nl = nand_271_cse & mux_tmp_127;
  assign mux_tmp_128 = MUX_s_1_2_2(and_1122_nl, mux_tmp_127, or_287_cse);
  assign and_1123_nl = nand_274_cse & mux_tmp_128;
  assign mux_tmp_129 = MUX_s_1_2_2(and_1123_nl, mux_tmp_128, or_280_cse);
  assign and_1124_nl = nand_276_cse & mux_tmp_129;
  assign mux_tmp_130 = MUX_s_1_2_2(and_1124_nl, mux_tmp_129, or_275_cse);
  assign nor_450_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_130));
  assign mux_133_nl = MUX_s_1_2_2(nor_450_nl, mux_tmp_130, or_270_cse);
  assign and_dcpl_451 = mux_133_nl & and_dcpl_31 & and_dcpl_38;
  assign nor_442_nl = ~(and_dcpl_30 | (~ or_tmp_263));
  assign or_352_nl = (rem_12cyc_st_9_1_0!=2'b11) | (rem_12cyc_st_9_3_2!=2'b00);
  assign mux_tmp_132 = MUX_s_1_2_2(nor_442_nl, or_tmp_263, or_352_nl);
  assign nor_443_nl = ~(and_dcpl_57 | (~ mux_tmp_132));
  assign mux_tmp_133 = MUX_s_1_2_2(nor_443_nl, mux_tmp_132, or_335_cse);
  assign nor_444_nl = ~(and_dcpl_84 | (~ mux_tmp_133));
  assign mux_tmp_134 = MUX_s_1_2_2(nor_444_nl, mux_tmp_133, or_320_cse);
  assign nor_445_nl = ~(and_dcpl_111 | (~ mux_tmp_134));
  assign mux_tmp_135 = MUX_s_1_2_2(nor_445_nl, mux_tmp_134, or_307_cse);
  assign and_1117_nl = nand_267_cse & mux_tmp_135;
  assign mux_tmp_136 = MUX_s_1_2_2(and_1117_nl, mux_tmp_135, or_296_cse);
  assign and_1118_nl = nand_271_cse & mux_tmp_136;
  assign mux_tmp_137 = MUX_s_1_2_2(and_1118_nl, mux_tmp_136, or_287_cse);
  assign and_1119_nl = nand_274_cse & mux_tmp_137;
  assign mux_tmp_138 = MUX_s_1_2_2(and_1119_nl, mux_tmp_137, or_280_cse);
  assign and_1120_nl = nand_276_cse & mux_tmp_138;
  assign mux_tmp_139 = MUX_s_1_2_2(and_1120_nl, mux_tmp_138, or_275_cse);
  assign nor_446_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_139));
  assign mux_142_nl = MUX_s_1_2_2(nor_446_nl, mux_tmp_139, or_270_cse);
  assign and_dcpl_454 = mux_142_nl & and_dcpl_4 & and_dcpl_11;
  assign nand_222_cse = ~((acc_1_tmp[1:0]==2'b11) & ccs_ccore_start_rsci_idat);
  assign and_tmp_89 = ((~ main_stage_0_8) | (~ asn_itm_7) | (rem_12cyc_st_7_1_0!=2'b11)
      | (rem_12cyc_st_7_3_2!=2'b00)) & ((~ main_stage_0_9) | (~ asn_itm_8) | (rem_12cyc_st_8_1_0!=2'b11)
      | (rem_12cyc_st_8_3_2!=2'b00)) & ((~ main_stage_0_10) | (~ asn_itm_9) | (rem_12cyc_st_9_1_0!=2'b11)
      | (rem_12cyc_st_9_3_2!=2'b00)) & ((~ main_stage_0_3) | (~ asn_itm_2) | (rem_12cyc_st_2_1_0!=2'b11)
      | (rem_12cyc_st_2_3_2!=2'b00)) & ((~ main_stage_0_4) | (~ asn_itm_3) | (rem_12cyc_st_3_1_0!=2'b11)
      | (rem_12cyc_st_3_3_2!=2'b00)) & ((~ main_stage_0_5) | (~ asn_itm_4) | (rem_12cyc_st_4_1_0!=2'b11)
      | (rem_12cyc_st_4_3_2!=2'b00)) & ((~ main_stage_0_6) | (~ asn_itm_5) | (rem_12cyc_st_5_1_0!=2'b11)
      | (rem_12cyc_st_5_3_2!=2'b00)) & ((~ main_stage_0_7) | (~ asn_itm_6) | (rem_12cyc_st_6_1_0!=2'b11)
      | (rem_12cyc_st_6_3_2!=2'b00)) & ((~ main_stage_0_11) | (~ asn_itm_10) | (rem_12cyc_st_10_1_0!=2'b11)
      | (rem_12cyc_st_10_3_2!=2'b00)) & ((acc_tmp!=2'b00) | nand_222_cse);
  assign nand_223_cse = ~((rem_12cyc_1_0==2'b11));
  assign and_1116_nl = nand_223_cse & and_tmp_89;
  assign or_362_nl = (~ main_stage_0_2) | (~ asn_itm_1) | (rem_12cyc_3_2!=2'b00);
  assign mux_tmp_141 = MUX_s_1_2_2(and_1116_nl, and_tmp_89, or_362_nl);
  assign and_dcpl_460 = ccs_ccore_start_rsci_idat & (acc_tmp==2'b01);
  assign and_dcpl_461 = and_dcpl_460 & and_dcpl_291;
  assign and_dcpl_462 = (rem_12cyc_st_2_3_2==2'b01);
  assign and_dcpl_463 = and_dcpl_462 & (~ (rem_12cyc_st_2_1_0[1]));
  assign not_tmp_332 = ~((rem_12cyc_3_2[0]) & asn_itm_1 & main_stage_0_2);
  assign or_tmp_368 = (rem_12cyc_1_0!=2'b00) | (rem_12cyc_3_2[1]) | not_tmp_332;
  assign nand_281_cse = ~((acc_tmp[0]) & ccs_ccore_start_rsci_idat);
  assign or_377_cse = (acc_1_tmp[1:0]!=2'b00) | (acc_tmp[1]);
  assign and_1172_nl = nand_281_cse & or_tmp_368;
  assign mux_144_nl = MUX_s_1_2_2(and_1172_nl, or_tmp_368, or_377_cse);
  assign and_dcpl_465 = mux_144_nl & and_dcpl_298 & and_dcpl_463;
  assign and_dcpl_466 = (rem_12cyc_st_3_3_2==2'b01);
  assign and_dcpl_467 = and_dcpl_466 & (~ (rem_12cyc_st_3_1_0[1]));
  assign or_382_cse = (rem_12cyc_st_2_1_0[1]) | (rem_12cyc_st_2_3_2!=2'b01) | (~
      asn_itm_2) | (~ main_stage_0_3) | (rem_12cyc_st_2_1_0[0]);
  assign and_tmp_90 = or_382_cse & or_tmp_368;
  assign and_1114_nl = nand_281_cse & and_tmp_90;
  assign mux_145_nl = MUX_s_1_2_2(and_1114_nl, and_tmp_90, or_377_cse);
  assign and_dcpl_469 = mux_145_nl & and_dcpl_304 & and_dcpl_467;
  assign and_dcpl_470 = (rem_12cyc_st_4_3_2==2'b01);
  assign and_dcpl_471 = and_dcpl_470 & (~ (rem_12cyc_st_4_1_0[1]));
  assign or_386_cse = (rem_12cyc_st_3_1_0[1]) | (rem_12cyc_st_3_3_2!=2'b01) | (~
      asn_itm_3) | (~ main_stage_0_4) | (rem_12cyc_st_3_1_0[0]);
  assign and_tmp_92 = or_382_cse & or_386_cse & or_tmp_368;
  assign and_1113_nl = nand_281_cse & and_tmp_92;
  assign mux_146_nl = MUX_s_1_2_2(and_1113_nl, and_tmp_92, or_377_cse);
  assign and_dcpl_473 = mux_146_nl & and_dcpl_310 & and_dcpl_471;
  assign and_dcpl_474 = (rem_12cyc_st_5_3_2==2'b01);
  assign and_dcpl_475 = and_dcpl_474 & (~ (rem_12cyc_st_5_1_0[1]));
  assign or_391_cse = (rem_12cyc_st_4_1_0[1]) | (rem_12cyc_st_4_3_2!=2'b01) | (~
      asn_itm_4) | (~ main_stage_0_5) | (rem_12cyc_st_4_1_0[0]);
  assign and_tmp_95 = or_382_cse & or_386_cse & or_391_cse & or_tmp_368;
  assign and_1112_nl = nand_281_cse & and_tmp_95;
  assign mux_147_nl = MUX_s_1_2_2(and_1112_nl, and_tmp_95, or_377_cse);
  assign and_dcpl_477 = mux_147_nl & and_dcpl_316 & and_dcpl_475;
  assign or_397_cse = (rem_12cyc_st_5_1_0[1]) | (rem_12cyc_st_5_3_2!=2'b01) | (~
      asn_itm_5) | (~ main_stage_0_6) | (rem_12cyc_st_5_1_0[0]);
  assign and_tmp_99 = or_382_cse & or_386_cse & or_391_cse & or_397_cse & or_tmp_368;
  assign and_1111_nl = nand_281_cse & and_tmp_99;
  assign mux_148_nl = MUX_s_1_2_2(and_1111_nl, and_tmp_99, or_377_cse);
  assign and_dcpl_480 = mux_148_nl & and_dcpl_121 & and_dcpl_110;
  assign nand_215_cse = ~((rem_12cyc_st_6_3_2[0]) & asn_itm_6 & main_stage_0_7);
  assign or_404_cse = (rem_12cyc_st_6_1_0!=2'b00) | (rem_12cyc_st_6_3_2[1]);
  assign and_1109_nl = nand_215_cse & or_tmp_368;
  assign mux_149_nl = MUX_s_1_2_2(and_1109_nl, or_tmp_368, or_404_cse);
  assign and_tmp_103 = or_382_cse & or_386_cse & or_391_cse & or_397_cse & mux_149_nl;
  assign and_1110_nl = nand_281_cse & and_tmp_103;
  assign mux_150_nl = MUX_s_1_2_2(and_1110_nl, and_tmp_103, or_377_cse);
  assign and_dcpl_483 = mux_150_nl & and_dcpl_94 & and_dcpl_83;
  assign nand_212_cse = ~((rem_12cyc_st_7_3_2[0]) & asn_itm_7 & main_stage_0_8);
  assign or_413_cse = (rem_12cyc_st_7_1_0!=2'b00) | (rem_12cyc_st_7_3_2[1]);
  assign and_1106_nl = nand_212_cse & or_tmp_368;
  assign mux_tmp_149 = MUX_s_1_2_2(and_1106_nl, or_tmp_368, or_413_cse);
  assign and_1107_nl = nand_215_cse & mux_tmp_149;
  assign mux_152_nl = MUX_s_1_2_2(and_1107_nl, mux_tmp_149, or_404_cse);
  assign and_tmp_107 = or_382_cse & or_386_cse & or_391_cse & or_397_cse & mux_152_nl;
  assign and_1108_nl = nand_281_cse & and_tmp_107;
  assign mux_153_nl = MUX_s_1_2_2(and_1108_nl, and_tmp_107, or_377_cse);
  assign and_dcpl_486 = mux_153_nl & and_dcpl_67 & and_dcpl_56;
  assign nand_208_cse = ~((rem_12cyc_st_8_3_2[0]) & asn_itm_8 & main_stage_0_9);
  assign or_424_cse = (rem_12cyc_st_8_1_0!=2'b00) | (rem_12cyc_st_8_3_2[1]);
  assign and_1102_nl = nand_208_cse & or_tmp_368;
  assign mux_tmp_152 = MUX_s_1_2_2(and_1102_nl, or_tmp_368, or_424_cse);
  assign and_1103_nl = nand_212_cse & mux_tmp_152;
  assign mux_tmp_153 = MUX_s_1_2_2(and_1103_nl, mux_tmp_152, or_413_cse);
  assign and_1104_nl = nand_215_cse & mux_tmp_153;
  assign mux_156_nl = MUX_s_1_2_2(and_1104_nl, mux_tmp_153, or_404_cse);
  assign and_tmp_111 = or_382_cse & or_386_cse & or_391_cse & or_397_cse & mux_156_nl;
  assign and_1105_nl = nand_281_cse & and_tmp_111;
  assign mux_157_nl = MUX_s_1_2_2(and_1105_nl, and_tmp_111, or_377_cse);
  assign and_dcpl_489 = mux_157_nl & and_dcpl_40 & and_dcpl_29;
  assign nand_203_cse = ~((rem_12cyc_st_9_3_2[0]) & asn_itm_9 & main_stage_0_10);
  assign and_1097_nl = nand_203_cse & or_tmp_368;
  assign or_437_nl = (rem_12cyc_st_9_1_0!=2'b00) | (rem_12cyc_st_9_3_2[1]);
  assign mux_tmp_156 = MUX_s_1_2_2(and_1097_nl, or_tmp_368, or_437_nl);
  assign and_1098_nl = nand_208_cse & mux_tmp_156;
  assign mux_tmp_157 = MUX_s_1_2_2(and_1098_nl, mux_tmp_156, or_424_cse);
  assign and_1099_nl = nand_212_cse & mux_tmp_157;
  assign mux_tmp_158 = MUX_s_1_2_2(and_1099_nl, mux_tmp_157, or_413_cse);
  assign and_1100_nl = nand_215_cse & mux_tmp_158;
  assign mux_161_nl = MUX_s_1_2_2(and_1100_nl, mux_tmp_158, or_404_cse);
  assign and_tmp_115 = or_382_cse & or_386_cse & or_391_cse & or_397_cse & mux_161_nl;
  assign and_1101_nl = nand_281_cse & and_tmp_115;
  assign mux_162_nl = MUX_s_1_2_2(and_1101_nl, and_tmp_115, or_377_cse);
  assign and_dcpl_492 = mux_162_nl & and_dcpl_13 & and_dcpl_2;
  assign and_tmp_125 = ((~ main_stage_0_2) | (~ asn_itm_1) | (rem_12cyc_3_2!=2'b01)
      | (rem_12cyc_1_0!=2'b00)) & ((~ main_stage_0_8) | (~ asn_itm_7) | (rem_12cyc_st_7_1_0!=2'b00)
      | (rem_12cyc_st_7_3_2!=2'b01)) & ((~ main_stage_0_9) | (~ asn_itm_8) | (rem_12cyc_st_8_1_0!=2'b00)
      | (rem_12cyc_st_8_3_2!=2'b01)) & ((~ main_stage_0_10) | (~ asn_itm_9) | (rem_12cyc_st_9_1_0!=2'b00)
      | (rem_12cyc_st_9_3_2!=2'b01)) & or_382_cse & or_386_cse & or_391_cse & or_397_cse
      & ((~ main_stage_0_7) | (~ asn_itm_6) | (rem_12cyc_st_6_1_0!=2'b00) | (rem_12cyc_st_6_3_2!=2'b01))
      & ((~ main_stage_0_11) | (~ asn_itm_10) | (rem_12cyc_st_10_1_0!=2'b00) | (rem_12cyc_st_10_3_2!=2'b01))
      & ((acc_tmp!=2'b01) | (acc_1_tmp[1:0]!=2'b00) | (~ ccs_ccore_start_rsci_idat));
  assign and_dcpl_498 = and_dcpl_460 & and_dcpl_355;
  assign or_tmp_446 = (rem_12cyc_1_0!=2'b01) | (rem_12cyc_3_2[1]) | not_tmp_332;
  assign or_458_cse = (acc_1_tmp[1:0]!=2'b01) | (acc_tmp[1]);
  assign and_1171_nl = nand_281_cse & or_tmp_446;
  assign mux_163_nl = MUX_s_1_2_2(and_1171_nl, or_tmp_446, or_458_cse);
  assign and_dcpl_500 = mux_163_nl & and_dcpl_358 & and_dcpl_463;
  assign or_463_cse = (rem_12cyc_st_2_1_0[1]) | (rem_12cyc_st_2_3_2!=2'b01);
  assign and_1094_nl = nand_276_cse & or_tmp_446;
  assign mux_tmp_162 = MUX_s_1_2_2(and_1094_nl, or_tmp_446, or_463_cse);
  assign and_1095_nl = nand_281_cse & mux_tmp_162;
  assign mux_165_nl = MUX_s_1_2_2(and_1095_nl, mux_tmp_162, or_458_cse);
  assign and_dcpl_502 = mux_165_nl & and_dcpl_362 & and_dcpl_467;
  assign nand_198_cse = ~((rem_12cyc_st_3_3_2[0]) & asn_itm_3 & main_stage_0_4 &
      (rem_12cyc_st_3_1_0[0]));
  assign or_468_cse = (rem_12cyc_st_3_1_0[1]) | (rem_12cyc_st_3_3_2[1]);
  assign and_1091_nl = nand_198_cse & or_tmp_446;
  assign mux_tmp_164 = MUX_s_1_2_2(and_1091_nl, or_tmp_446, or_468_cse);
  assign and_1092_nl = nand_276_cse & mux_tmp_164;
  assign mux_tmp_165 = MUX_s_1_2_2(and_1092_nl, mux_tmp_164, or_463_cse);
  assign and_1093_nl = nand_281_cse & mux_tmp_165;
  assign mux_168_nl = MUX_s_1_2_2(and_1093_nl, mux_tmp_165, or_458_cse);
  assign and_dcpl_504 = mux_168_nl & and_dcpl_366 & and_dcpl_471;
  assign or_475_cse = (rem_12cyc_st_4_1_0[1]) | (rem_12cyc_st_4_3_2!=2'b01);
  assign and_1087_nl = nand_271_cse & or_tmp_446;
  assign mux_tmp_167 = MUX_s_1_2_2(and_1087_nl, or_tmp_446, or_475_cse);
  assign and_1088_nl = nand_198_cse & mux_tmp_167;
  assign mux_tmp_168 = MUX_s_1_2_2(and_1088_nl, mux_tmp_167, or_468_cse);
  assign and_1089_nl = nand_276_cse & mux_tmp_168;
  assign mux_tmp_169 = MUX_s_1_2_2(and_1089_nl, mux_tmp_168, or_463_cse);
  assign and_1090_nl = nand_281_cse & mux_tmp_169;
  assign mux_172_nl = MUX_s_1_2_2(and_1090_nl, mux_tmp_169, or_458_cse);
  assign and_dcpl_506 = mux_172_nl & and_dcpl_370 & and_dcpl_475;
  assign nand_189_cse = ~((rem_12cyc_st_5_3_2[0]) & asn_itm_5 & main_stage_0_6 &
      (rem_12cyc_st_5_1_0[0]));
  assign or_484_cse = (rem_12cyc_st_5_1_0[1]) | (rem_12cyc_st_5_3_2[1]);
  assign and_1082_nl = nand_189_cse & or_tmp_446;
  assign mux_tmp_171 = MUX_s_1_2_2(and_1082_nl, or_tmp_446, or_484_cse);
  assign and_1083_nl = nand_271_cse & mux_tmp_171;
  assign mux_tmp_172 = MUX_s_1_2_2(and_1083_nl, mux_tmp_171, or_475_cse);
  assign and_1084_nl = nand_198_cse & mux_tmp_172;
  assign mux_tmp_173 = MUX_s_1_2_2(and_1084_nl, mux_tmp_172, or_468_cse);
  assign and_1085_nl = nand_276_cse & mux_tmp_173;
  assign mux_tmp_174 = MUX_s_1_2_2(and_1085_nl, mux_tmp_173, or_463_cse);
  assign and_1086_nl = nand_281_cse & mux_tmp_174;
  assign mux_177_nl = MUX_s_1_2_2(and_1086_nl, mux_tmp_174, or_458_cse);
  assign and_dcpl_508 = mux_177_nl & and_dcpl_121 & and_dcpl_115;
  assign or_495_cse = (rem_12cyc_st_6_1_0!=2'b01) | (rem_12cyc_st_6_3_2[1]);
  assign and_1076_nl = nand_215_cse & or_tmp_446;
  assign mux_tmp_176 = MUX_s_1_2_2(and_1076_nl, or_tmp_446, or_495_cse);
  assign and_1077_nl = nand_189_cse & mux_tmp_176;
  assign mux_tmp_177 = MUX_s_1_2_2(and_1077_nl, mux_tmp_176, or_484_cse);
  assign and_1078_nl = nand_271_cse & mux_tmp_177;
  assign mux_tmp_178 = MUX_s_1_2_2(and_1078_nl, mux_tmp_177, or_475_cse);
  assign and_1079_nl = nand_198_cse & mux_tmp_178;
  assign mux_tmp_179 = MUX_s_1_2_2(and_1079_nl, mux_tmp_178, or_468_cse);
  assign and_1080_nl = nand_276_cse & mux_tmp_179;
  assign mux_tmp_180 = MUX_s_1_2_2(and_1080_nl, mux_tmp_179, or_463_cse);
  assign and_1081_nl = nand_281_cse & mux_tmp_180;
  assign mux_183_nl = MUX_s_1_2_2(and_1081_nl, mux_tmp_180, or_458_cse);
  assign and_dcpl_510 = mux_183_nl & and_dcpl_94 & and_dcpl_87;
  assign or_508_cse = (rem_12cyc_st_7_1_0!=2'b01) | (rem_12cyc_st_7_3_2[1]);
  assign and_1069_nl = nand_212_cse & or_tmp_446;
  assign mux_tmp_182 = MUX_s_1_2_2(and_1069_nl, or_tmp_446, or_508_cse);
  assign and_1070_nl = nand_215_cse & mux_tmp_182;
  assign mux_tmp_183 = MUX_s_1_2_2(and_1070_nl, mux_tmp_182, or_495_cse);
  assign and_1071_nl = nand_189_cse & mux_tmp_183;
  assign mux_tmp_184 = MUX_s_1_2_2(and_1071_nl, mux_tmp_183, or_484_cse);
  assign and_1072_nl = nand_271_cse & mux_tmp_184;
  assign mux_tmp_185 = MUX_s_1_2_2(and_1072_nl, mux_tmp_184, or_475_cse);
  assign and_1073_nl = nand_198_cse & mux_tmp_185;
  assign mux_tmp_186 = MUX_s_1_2_2(and_1073_nl, mux_tmp_185, or_468_cse);
  assign and_1074_nl = nand_276_cse & mux_tmp_186;
  assign mux_tmp_187 = MUX_s_1_2_2(and_1074_nl, mux_tmp_186, or_463_cse);
  assign and_1075_nl = nand_281_cse & mux_tmp_187;
  assign mux_190_nl = MUX_s_1_2_2(and_1075_nl, mux_tmp_187, or_458_cse);
  assign and_dcpl_512 = mux_190_nl & and_dcpl_67 & and_dcpl_60;
  assign or_523_cse = (rem_12cyc_st_8_1_0!=2'b01) | (rem_12cyc_st_8_3_2[1]);
  assign and_1061_nl = nand_208_cse & or_tmp_446;
  assign mux_tmp_189 = MUX_s_1_2_2(and_1061_nl, or_tmp_446, or_523_cse);
  assign and_1062_nl = nand_212_cse & mux_tmp_189;
  assign mux_tmp_190 = MUX_s_1_2_2(and_1062_nl, mux_tmp_189, or_508_cse);
  assign and_1063_nl = nand_215_cse & mux_tmp_190;
  assign mux_tmp_191 = MUX_s_1_2_2(and_1063_nl, mux_tmp_190, or_495_cse);
  assign and_1064_nl = nand_189_cse & mux_tmp_191;
  assign mux_tmp_192 = MUX_s_1_2_2(and_1064_nl, mux_tmp_191, or_484_cse);
  assign and_1065_nl = nand_271_cse & mux_tmp_192;
  assign mux_tmp_193 = MUX_s_1_2_2(and_1065_nl, mux_tmp_192, or_475_cse);
  assign and_1066_nl = nand_198_cse & mux_tmp_193;
  assign mux_tmp_194 = MUX_s_1_2_2(and_1066_nl, mux_tmp_193, or_468_cse);
  assign and_1067_nl = nand_276_cse & mux_tmp_194;
  assign mux_tmp_195 = MUX_s_1_2_2(and_1067_nl, mux_tmp_194, or_463_cse);
  assign and_1068_nl = nand_281_cse & mux_tmp_195;
  assign mux_198_nl = MUX_s_1_2_2(and_1068_nl, mux_tmp_195, or_458_cse);
  assign and_dcpl_514 = mux_198_nl & and_dcpl_40 & and_dcpl_33;
  assign and_1052_nl = nand_203_cse & or_tmp_446;
  assign or_540_nl = (rem_12cyc_st_9_1_0!=2'b01) | (rem_12cyc_st_9_3_2[1]);
  assign mux_tmp_197 = MUX_s_1_2_2(and_1052_nl, or_tmp_446, or_540_nl);
  assign and_1053_nl = nand_208_cse & mux_tmp_197;
  assign mux_tmp_198 = MUX_s_1_2_2(and_1053_nl, mux_tmp_197, or_523_cse);
  assign and_1054_nl = nand_212_cse & mux_tmp_198;
  assign mux_tmp_199 = MUX_s_1_2_2(and_1054_nl, mux_tmp_198, or_508_cse);
  assign and_1055_nl = nand_215_cse & mux_tmp_199;
  assign mux_tmp_200 = MUX_s_1_2_2(and_1055_nl, mux_tmp_199, or_495_cse);
  assign and_1056_nl = nand_189_cse & mux_tmp_200;
  assign mux_tmp_201 = MUX_s_1_2_2(and_1056_nl, mux_tmp_200, or_484_cse);
  assign and_1057_nl = nand_271_cse & mux_tmp_201;
  assign mux_tmp_202 = MUX_s_1_2_2(and_1057_nl, mux_tmp_201, or_475_cse);
  assign and_1058_nl = nand_198_cse & mux_tmp_202;
  assign mux_tmp_203 = MUX_s_1_2_2(and_1058_nl, mux_tmp_202, or_468_cse);
  assign and_1059_nl = nand_276_cse & mux_tmp_203;
  assign mux_tmp_204 = MUX_s_1_2_2(and_1059_nl, mux_tmp_203, or_463_cse);
  assign and_1060_nl = nand_281_cse & mux_tmp_204;
  assign mux_207_nl = MUX_s_1_2_2(and_1060_nl, mux_tmp_204, or_458_cse);
  assign and_dcpl_516 = mux_207_nl & and_dcpl_13 & and_dcpl_6;
  assign and_tmp_134 = ((~ main_stage_0_8) | (~ asn_itm_7) | (rem_12cyc_st_7_1_0!=2'b01)
      | (rem_12cyc_st_7_3_2!=2'b01)) & ((~ main_stage_0_9) | (~ asn_itm_8) | (rem_12cyc_st_8_1_0!=2'b01)
      | (rem_12cyc_st_8_3_2!=2'b01)) & ((~ main_stage_0_10) | (~ asn_itm_9) | (rem_12cyc_st_9_1_0!=2'b01)
      | (rem_12cyc_st_9_3_2!=2'b01)) & ((~ main_stage_0_3) | (~ asn_itm_2) | (rem_12cyc_st_2_1_0!=2'b01)
      | (rem_12cyc_st_2_3_2!=2'b01)) & ((~ main_stage_0_4) | (~ asn_itm_3) | (rem_12cyc_st_3_1_0!=2'b01)
      | (rem_12cyc_st_3_3_2!=2'b01)) & ((~ main_stage_0_5) | (~ asn_itm_4) | (rem_12cyc_st_4_1_0!=2'b01)
      | (rem_12cyc_st_4_3_2!=2'b01)) & ((~ main_stage_0_6) | (~ asn_itm_5) | (rem_12cyc_st_5_1_0!=2'b01)
      | (rem_12cyc_st_5_3_2!=2'b01)) & ((~ main_stage_0_7) | (~ asn_itm_6) | (rem_12cyc_st_6_1_0!=2'b01)
      | (rem_12cyc_st_6_3_2!=2'b01)) & ((~ main_stage_0_11) | (~ asn_itm_10) | (rem_12cyc_st_10_1_0!=2'b01)
      | (rem_12cyc_st_10_3_2!=2'b01)) & ((acc_tmp!=2'b01) | (acc_1_tmp[1]) | nand_250_cse);
  assign nor_439_nl = ~((rem_12cyc_1_0[0]) | (~ and_tmp_134));
  assign or_550_nl = (~ main_stage_0_2) | (~ asn_itm_1) | (rem_12cyc_3_2!=2'b01)
      | (rem_12cyc_1_0[1]);
  assign mux_tmp_206 = MUX_s_1_2_2(nor_439_nl, and_tmp_134, or_550_nl);
  assign and_dcpl_520 = and_dcpl_460 & and_dcpl_393;
  assign and_dcpl_521 = and_dcpl_462 & (rem_12cyc_st_2_1_0[1]);
  assign or_tmp_551 = (rem_12cyc_1_0!=2'b10) | (rem_12cyc_3_2[1]) | not_tmp_332;
  assign or_564_cse = (acc_1_tmp[1:0]!=2'b10) | (acc_tmp[1]);
  assign and_1170_nl = nand_281_cse & or_tmp_551;
  assign mux_209_nl = MUX_s_1_2_2(and_1170_nl, or_tmp_551, or_564_cse);
  assign and_dcpl_523 = mux_209_nl & and_dcpl_298 & and_dcpl_521;
  assign and_dcpl_524 = and_dcpl_466 & (rem_12cyc_st_3_1_0[1]);
  assign or_569_cse = (~ (rem_12cyc_st_2_1_0[1])) | (rem_12cyc_st_2_3_2!=2'b01) |
      (~ asn_itm_2) | (~ main_stage_0_3) | (rem_12cyc_st_2_1_0[0]);
  assign and_tmp_135 = or_569_cse & or_tmp_551;
  assign and_1050_nl = nand_281_cse & and_tmp_135;
  assign mux_210_nl = MUX_s_1_2_2(and_1050_nl, and_tmp_135, or_564_cse);
  assign and_dcpl_526 = mux_210_nl & and_dcpl_304 & and_dcpl_524;
  assign and_dcpl_527 = and_dcpl_470 & (rem_12cyc_st_4_1_0[1]);
  assign or_573_cse = (~ (rem_12cyc_st_3_1_0[1])) | (rem_12cyc_st_3_3_2!=2'b01) |
      (~ asn_itm_3) | (~ main_stage_0_4) | (rem_12cyc_st_3_1_0[0]);
  assign and_tmp_137 = or_569_cse & or_573_cse & or_tmp_551;
  assign and_1049_nl = nand_281_cse & and_tmp_137;
  assign mux_211_nl = MUX_s_1_2_2(and_1049_nl, and_tmp_137, or_564_cse);
  assign and_dcpl_529 = mux_211_nl & and_dcpl_310 & and_dcpl_527;
  assign and_dcpl_530 = and_dcpl_474 & (rem_12cyc_st_5_1_0[1]);
  assign or_578_cse = (~ (rem_12cyc_st_4_1_0[1])) | (rem_12cyc_st_4_3_2!=2'b01) |
      (~ asn_itm_4) | (~ main_stage_0_5) | (rem_12cyc_st_4_1_0[0]);
  assign and_tmp_140 = or_569_cse & or_573_cse & or_578_cse & or_tmp_551;
  assign and_1048_nl = nand_281_cse & and_tmp_140;
  assign mux_212_nl = MUX_s_1_2_2(and_1048_nl, and_tmp_140, or_564_cse);
  assign and_dcpl_532 = mux_212_nl & and_dcpl_316 & and_dcpl_530;
  assign or_584_cse = (~ (rem_12cyc_st_5_1_0[1])) | (rem_12cyc_st_5_3_2!=2'b01) |
      (~ asn_itm_5) | (~ main_stage_0_6) | (rem_12cyc_st_5_1_0[0]);
  assign and_tmp_144 = or_569_cse & or_573_cse & or_578_cse & or_584_cse & or_tmp_551;
  assign and_1047_nl = nand_281_cse & and_tmp_144;
  assign mux_213_nl = MUX_s_1_2_2(and_1047_nl, and_tmp_144, or_564_cse);
  assign and_dcpl_534 = mux_213_nl & and_dcpl_121 & and_dcpl_117;
  assign or_591_cse = (rem_12cyc_st_6_1_0!=2'b10) | (rem_12cyc_st_6_3_2[1]);
  assign and_1045_nl = nand_215_cse & or_tmp_551;
  assign mux_214_nl = MUX_s_1_2_2(and_1045_nl, or_tmp_551, or_591_cse);
  assign and_tmp_148 = or_569_cse & or_573_cse & or_578_cse & or_584_cse & mux_214_nl;
  assign and_1046_nl = nand_281_cse & and_tmp_148;
  assign mux_215_nl = MUX_s_1_2_2(and_1046_nl, and_tmp_148, or_564_cse);
  assign and_dcpl_536 = mux_215_nl & and_dcpl_94 & and_dcpl_90;
  assign or_600_cse = (rem_12cyc_st_7_1_0!=2'b10) | (rem_12cyc_st_7_3_2[1]);
  assign and_1042_nl = nand_212_cse & or_tmp_551;
  assign mux_tmp_214 = MUX_s_1_2_2(and_1042_nl, or_tmp_551, or_600_cse);
  assign and_1043_nl = nand_215_cse & mux_tmp_214;
  assign mux_217_nl = MUX_s_1_2_2(and_1043_nl, mux_tmp_214, or_591_cse);
  assign and_tmp_152 = or_569_cse & or_573_cse & or_578_cse & or_584_cse & mux_217_nl;
  assign and_1044_nl = nand_281_cse & and_tmp_152;
  assign mux_218_nl = MUX_s_1_2_2(and_1044_nl, and_tmp_152, or_564_cse);
  assign and_dcpl_538 = mux_218_nl & and_dcpl_67 & and_dcpl_63;
  assign or_611_cse = (rem_12cyc_st_8_1_0!=2'b10) | (rem_12cyc_st_8_3_2[1]);
  assign and_1038_nl = nand_208_cse & or_tmp_551;
  assign mux_tmp_217 = MUX_s_1_2_2(and_1038_nl, or_tmp_551, or_611_cse);
  assign and_1039_nl = nand_212_cse & mux_tmp_217;
  assign mux_tmp_218 = MUX_s_1_2_2(and_1039_nl, mux_tmp_217, or_600_cse);
  assign and_1040_nl = nand_215_cse & mux_tmp_218;
  assign mux_221_nl = MUX_s_1_2_2(and_1040_nl, mux_tmp_218, or_591_cse);
  assign and_tmp_156 = or_569_cse & or_573_cse & or_578_cse & or_584_cse & mux_221_nl;
  assign and_1041_nl = nand_281_cse & and_tmp_156;
  assign mux_222_nl = MUX_s_1_2_2(and_1041_nl, and_tmp_156, or_564_cse);
  assign and_dcpl_540 = mux_222_nl & and_dcpl_40 & and_dcpl_36;
  assign and_1033_nl = nand_203_cse & or_tmp_551;
  assign or_624_nl = (rem_12cyc_st_9_1_0!=2'b10) | (rem_12cyc_st_9_3_2[1]);
  assign mux_tmp_221 = MUX_s_1_2_2(and_1033_nl, or_tmp_551, or_624_nl);
  assign and_1034_nl = nand_208_cse & mux_tmp_221;
  assign mux_tmp_222 = MUX_s_1_2_2(and_1034_nl, mux_tmp_221, or_611_cse);
  assign and_1035_nl = nand_212_cse & mux_tmp_222;
  assign mux_tmp_223 = MUX_s_1_2_2(and_1035_nl, mux_tmp_222, or_600_cse);
  assign and_1036_nl = nand_215_cse & mux_tmp_223;
  assign mux_226_nl = MUX_s_1_2_2(and_1036_nl, mux_tmp_223, or_591_cse);
  assign and_tmp_160 = or_569_cse & or_573_cse & or_578_cse & or_584_cse & mux_226_nl;
  assign and_1037_nl = nand_281_cse & and_tmp_160;
  assign mux_227_nl = MUX_s_1_2_2(and_1037_nl, and_tmp_160, or_564_cse);
  assign and_dcpl_542 = mux_227_nl & and_dcpl_13 & and_dcpl_9;
  assign and_tmp_170 = ((~ main_stage_0_2) | (~ asn_itm_1) | (rem_12cyc_3_2!=2'b01)
      | (rem_12cyc_1_0!=2'b10)) & ((~ main_stage_0_8) | (~ asn_itm_7) | (rem_12cyc_st_7_1_0!=2'b10)
      | (rem_12cyc_st_7_3_2!=2'b01)) & ((~ main_stage_0_9) | (~ asn_itm_8) | (rem_12cyc_st_8_1_0!=2'b10)
      | (rem_12cyc_st_8_3_2!=2'b01)) & ((~ main_stage_0_10) | (~ asn_itm_9) | (rem_12cyc_st_9_1_0!=2'b10)
      | (rem_12cyc_st_9_3_2!=2'b01)) & or_569_cse & or_573_cse & or_578_cse & or_584_cse
      & ((~ main_stage_0_7) | (~ asn_itm_6) | (rem_12cyc_st_6_1_0!=2'b10) | (rem_12cyc_st_6_3_2!=2'b01))
      & ((~ main_stage_0_11) | (~ asn_itm_10) | (rem_12cyc_st_10_1_0!=2'b10) | (rem_12cyc_st_10_3_2!=2'b01))
      & ((acc_tmp!=2'b01) | (acc_1_tmp[1:0]!=2'b10) | (~ ccs_ccore_start_rsci_idat));
  assign and_dcpl_546 = and_dcpl_460 & and_dcpl_430;
  assign or_tmp_629 = (rem_12cyc_1_0!=2'b11) | (rem_12cyc_3_2[1]) | not_tmp_332;
  assign or_643_cse = (acc_1_tmp[1:0]!=2'b11) | (acc_tmp[1]);
  assign and_1169_nl = nand_281_cse & or_tmp_629;
  assign mux_228_nl = MUX_s_1_2_2(and_1169_nl, or_tmp_629, or_643_cse);
  assign and_dcpl_548 = mux_228_nl & and_dcpl_358 & and_dcpl_521;
  assign or_648_cse = (~ (rem_12cyc_st_2_1_0[1])) | (rem_12cyc_st_2_3_2!=2'b01);
  assign and_1030_nl = nand_276_cse & or_tmp_629;
  assign mux_tmp_227 = MUX_s_1_2_2(and_1030_nl, or_tmp_629, or_648_cse);
  assign and_1031_nl = nand_281_cse & mux_tmp_227;
  assign mux_230_nl = MUX_s_1_2_2(and_1031_nl, mux_tmp_227, or_643_cse);
  assign and_dcpl_550 = mux_230_nl & and_dcpl_362 & and_dcpl_524;
  assign or_653_cse = (~ (rem_12cyc_st_3_1_0[1])) | (rem_12cyc_st_3_3_2[1]);
  assign and_1027_nl = nand_198_cse & or_tmp_629;
  assign mux_tmp_229 = MUX_s_1_2_2(and_1027_nl, or_tmp_629, or_653_cse);
  assign and_1028_nl = nand_276_cse & mux_tmp_229;
  assign mux_tmp_230 = MUX_s_1_2_2(and_1028_nl, mux_tmp_229, or_648_cse);
  assign and_1029_nl = nand_281_cse & mux_tmp_230;
  assign mux_233_nl = MUX_s_1_2_2(and_1029_nl, mux_tmp_230, or_643_cse);
  assign and_dcpl_552 = mux_233_nl & and_dcpl_366 & and_dcpl_527;
  assign or_660_cse = (~ (rem_12cyc_st_4_1_0[1])) | (rem_12cyc_st_4_3_2!=2'b01);
  assign and_1023_nl = nand_271_cse & or_tmp_629;
  assign mux_tmp_232 = MUX_s_1_2_2(and_1023_nl, or_tmp_629, or_660_cse);
  assign and_1024_nl = nand_198_cse & mux_tmp_232;
  assign mux_tmp_233 = MUX_s_1_2_2(and_1024_nl, mux_tmp_232, or_653_cse);
  assign and_1025_nl = nand_276_cse & mux_tmp_233;
  assign mux_tmp_234 = MUX_s_1_2_2(and_1025_nl, mux_tmp_233, or_648_cse);
  assign and_1026_nl = nand_281_cse & mux_tmp_234;
  assign mux_237_nl = MUX_s_1_2_2(and_1026_nl, mux_tmp_234, or_643_cse);
  assign and_dcpl_554 = mux_237_nl & and_dcpl_370 & and_dcpl_530;
  assign or_669_cse = (~ (rem_12cyc_st_5_1_0[1])) | (rem_12cyc_st_5_3_2[1]);
  assign and_1018_nl = nand_189_cse & or_tmp_629;
  assign mux_tmp_236 = MUX_s_1_2_2(and_1018_nl, or_tmp_629, or_669_cse);
  assign and_1019_nl = nand_271_cse & mux_tmp_236;
  assign mux_tmp_237 = MUX_s_1_2_2(and_1019_nl, mux_tmp_236, or_660_cse);
  assign and_1020_nl = nand_198_cse & mux_tmp_237;
  assign mux_tmp_238 = MUX_s_1_2_2(and_1020_nl, mux_tmp_237, or_653_cse);
  assign and_1021_nl = nand_276_cse & mux_tmp_238;
  assign mux_tmp_239 = MUX_s_1_2_2(and_1021_nl, mux_tmp_238, or_648_cse);
  assign and_1022_nl = nand_281_cse & mux_tmp_239;
  assign mux_242_nl = MUX_s_1_2_2(and_1022_nl, mux_tmp_239, or_643_cse);
  assign and_dcpl_556 = mux_242_nl & and_dcpl_121 & and_dcpl_119;
  assign or_680_cse = (rem_12cyc_st_6_1_0!=2'b11) | (rem_12cyc_st_6_3_2[1]);
  assign and_1012_nl = nand_215_cse & or_tmp_629;
  assign mux_tmp_241 = MUX_s_1_2_2(and_1012_nl, or_tmp_629, or_680_cse);
  assign and_1013_nl = nand_189_cse & mux_tmp_241;
  assign mux_tmp_242 = MUX_s_1_2_2(and_1013_nl, mux_tmp_241, or_669_cse);
  assign and_1014_nl = nand_271_cse & mux_tmp_242;
  assign mux_tmp_243 = MUX_s_1_2_2(and_1014_nl, mux_tmp_242, or_660_cse);
  assign and_1015_nl = nand_198_cse & mux_tmp_243;
  assign mux_tmp_244 = MUX_s_1_2_2(and_1015_nl, mux_tmp_243, or_653_cse);
  assign and_1016_nl = nand_276_cse & mux_tmp_244;
  assign mux_tmp_245 = MUX_s_1_2_2(and_1016_nl, mux_tmp_244, or_648_cse);
  assign and_1017_nl = nand_281_cse & mux_tmp_245;
  assign mux_248_nl = MUX_s_1_2_2(and_1017_nl, mux_tmp_245, or_643_cse);
  assign and_dcpl_558 = mux_248_nl & and_dcpl_94 & and_dcpl_92;
  assign or_693_cse = (rem_12cyc_st_7_1_0!=2'b11) | (rem_12cyc_st_7_3_2[1]);
  assign and_1005_nl = nand_212_cse & or_tmp_629;
  assign mux_tmp_247 = MUX_s_1_2_2(and_1005_nl, or_tmp_629, or_693_cse);
  assign and_1006_nl = nand_215_cse & mux_tmp_247;
  assign mux_tmp_248 = MUX_s_1_2_2(and_1006_nl, mux_tmp_247, or_680_cse);
  assign and_1007_nl = nand_189_cse & mux_tmp_248;
  assign mux_tmp_249 = MUX_s_1_2_2(and_1007_nl, mux_tmp_248, or_669_cse);
  assign and_1008_nl = nand_271_cse & mux_tmp_249;
  assign mux_tmp_250 = MUX_s_1_2_2(and_1008_nl, mux_tmp_249, or_660_cse);
  assign and_1009_nl = nand_198_cse & mux_tmp_250;
  assign mux_tmp_251 = MUX_s_1_2_2(and_1009_nl, mux_tmp_250, or_653_cse);
  assign and_1010_nl = nand_276_cse & mux_tmp_251;
  assign mux_tmp_252 = MUX_s_1_2_2(and_1010_nl, mux_tmp_251, or_648_cse);
  assign and_1011_nl = nand_281_cse & mux_tmp_252;
  assign mux_255_nl = MUX_s_1_2_2(and_1011_nl, mux_tmp_252, or_643_cse);
  assign and_dcpl_560 = mux_255_nl & and_dcpl_67 & and_dcpl_65;
  assign or_708_cse = (rem_12cyc_st_8_1_0!=2'b11) | (rem_12cyc_st_8_3_2[1]);
  assign and_997_nl = nand_208_cse & or_tmp_629;
  assign mux_tmp_254 = MUX_s_1_2_2(and_997_nl, or_tmp_629, or_708_cse);
  assign and_998_nl = nand_212_cse & mux_tmp_254;
  assign mux_tmp_255 = MUX_s_1_2_2(and_998_nl, mux_tmp_254, or_693_cse);
  assign and_999_nl = nand_215_cse & mux_tmp_255;
  assign mux_tmp_256 = MUX_s_1_2_2(and_999_nl, mux_tmp_255, or_680_cse);
  assign and_1000_nl = nand_189_cse & mux_tmp_256;
  assign mux_tmp_257 = MUX_s_1_2_2(and_1000_nl, mux_tmp_256, or_669_cse);
  assign and_1001_nl = nand_271_cse & mux_tmp_257;
  assign mux_tmp_258 = MUX_s_1_2_2(and_1001_nl, mux_tmp_257, or_660_cse);
  assign and_1002_nl = nand_198_cse & mux_tmp_258;
  assign mux_tmp_259 = MUX_s_1_2_2(and_1002_nl, mux_tmp_258, or_653_cse);
  assign and_1003_nl = nand_276_cse & mux_tmp_259;
  assign mux_tmp_260 = MUX_s_1_2_2(and_1003_nl, mux_tmp_259, or_648_cse);
  assign and_1004_nl = nand_281_cse & mux_tmp_260;
  assign mux_263_nl = MUX_s_1_2_2(and_1004_nl, mux_tmp_260, or_643_cse);
  assign and_dcpl_562 = mux_263_nl & and_dcpl_40 & and_dcpl_38;
  assign and_988_nl = nand_203_cse & or_tmp_629;
  assign or_725_nl = (rem_12cyc_st_9_1_0!=2'b11) | (rem_12cyc_st_9_3_2[1]);
  assign mux_tmp_262 = MUX_s_1_2_2(and_988_nl, or_tmp_629, or_725_nl);
  assign and_989_nl = nand_208_cse & mux_tmp_262;
  assign mux_tmp_263 = MUX_s_1_2_2(and_989_nl, mux_tmp_262, or_708_cse);
  assign and_990_nl = nand_212_cse & mux_tmp_263;
  assign mux_tmp_264 = MUX_s_1_2_2(and_990_nl, mux_tmp_263, or_693_cse);
  assign and_991_nl = nand_215_cse & mux_tmp_264;
  assign mux_tmp_265 = MUX_s_1_2_2(and_991_nl, mux_tmp_264, or_680_cse);
  assign and_992_nl = nand_189_cse & mux_tmp_265;
  assign mux_tmp_266 = MUX_s_1_2_2(and_992_nl, mux_tmp_265, or_669_cse);
  assign and_993_nl = nand_271_cse & mux_tmp_266;
  assign mux_tmp_267 = MUX_s_1_2_2(and_993_nl, mux_tmp_266, or_660_cse);
  assign and_994_nl = nand_198_cse & mux_tmp_267;
  assign mux_tmp_268 = MUX_s_1_2_2(and_994_nl, mux_tmp_267, or_653_cse);
  assign and_995_nl = nand_276_cse & mux_tmp_268;
  assign mux_tmp_269 = MUX_s_1_2_2(and_995_nl, mux_tmp_268, or_648_cse);
  assign and_996_nl = nand_281_cse & mux_tmp_269;
  assign mux_272_nl = MUX_s_1_2_2(and_996_nl, mux_tmp_269, or_643_cse);
  assign and_dcpl_564 = mux_272_nl & and_dcpl_13 & and_dcpl_11;
  assign and_tmp_179 = (~(main_stage_0_8 & asn_itm_7 & (rem_12cyc_st_7_1_0==2'b11)
      & (rem_12cyc_st_7_3_2==2'b01))) & (~(main_stage_0_9 & asn_itm_8 & (rem_12cyc_st_8_1_0==2'b11)
      & (rem_12cyc_st_8_3_2==2'b01))) & (~(main_stage_0_10 & asn_itm_9 & (rem_12cyc_st_9_1_0==2'b11)
      & (rem_12cyc_st_9_3_2==2'b01))) & (~(main_stage_0_3 & asn_itm_2 & (rem_12cyc_st_2_1_0==2'b11)
      & (rem_12cyc_st_2_3_2==2'b01))) & (~(main_stage_0_4 & asn_itm_3 & (rem_12cyc_st_3_1_0==2'b11)
      & (rem_12cyc_st_3_3_2==2'b01))) & (~(main_stage_0_5 & asn_itm_4 & (rem_12cyc_st_4_1_0==2'b11)
      & (rem_12cyc_st_4_3_2==2'b01))) & (~(main_stage_0_6 & asn_itm_5 & (rem_12cyc_st_5_1_0==2'b11)
      & (rem_12cyc_st_5_3_2==2'b01))) & (~(main_stage_0_7 & asn_itm_6 & (rem_12cyc_st_6_1_0==2'b11)
      & (rem_12cyc_st_6_3_2==2'b01))) & (~(main_stage_0_11 & asn_itm_10 & (rem_12cyc_st_10_1_0==2'b11)
      & (rem_12cyc_st_10_3_2==2'b01))) & ((acc_tmp[1]) | (~((acc_tmp[0]) & (acc_1_tmp[1:0]==2'b11)
      & ccs_ccore_start_rsci_idat)));
  assign and_987_nl = (~((rem_12cyc_3_2[0]) & (rem_12cyc_1_0==2'b11))) & and_tmp_179;
  assign or_735_nl = (~ main_stage_0_2) | (~ asn_itm_1) | (rem_12cyc_3_2[1]);
  assign mux_tmp_271 = MUX_s_1_2_2(and_987_nl, and_tmp_179, or_735_nl);
  assign and_dcpl_568 = and_dcpl_292 & (acc_tmp[1]);
  assign and_dcpl_569 = and_dcpl_568 & and_dcpl_291;
  assign and_dcpl_570 = (rem_12cyc_st_2_3_2==2'b10);
  assign and_dcpl_571 = and_dcpl_570 & (~ (rem_12cyc_st_2_1_0[1]));
  assign or_tmp_733 = (rem_12cyc_1_0!=2'b00) | (rem_12cyc_3_2!=2'b10) | not_tmp_54;
  assign or_748_cse = (acc_1_tmp[1:0]!=2'b00) | (acc_tmp!=2'b10);
  assign nor_436_nl = ~(ccs_ccore_start_rsci_idat | (~ or_tmp_733));
  assign mux_274_nl = MUX_s_1_2_2(nor_436_nl, or_tmp_733, or_748_cse);
  assign and_dcpl_573 = mux_274_nl & and_dcpl_298 & and_dcpl_571;
  assign and_dcpl_574 = (rem_12cyc_st_3_3_2==2'b10);
  assign and_dcpl_575 = and_dcpl_574 & (~ (rem_12cyc_st_3_1_0[1]));
  assign or_753_cse = (rem_12cyc_st_2_1_0[1]) | (rem_12cyc_st_2_3_2!=2'b10) | (~
      asn_itm_2) | (~ main_stage_0_3) | (rem_12cyc_st_2_1_0[0]);
  assign and_tmp_180 = or_753_cse & or_tmp_733;
  assign nor_435_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_180));
  assign mux_275_nl = MUX_s_1_2_2(nor_435_nl, and_tmp_180, or_748_cse);
  assign and_dcpl_577 = mux_275_nl & and_dcpl_304 & and_dcpl_575;
  assign and_dcpl_578 = (rem_12cyc_st_4_3_2==2'b10);
  assign and_dcpl_579 = and_dcpl_578 & (~ (rem_12cyc_st_4_1_0[1]));
  assign or_757_cse = (rem_12cyc_st_3_1_0[1]) | (rem_12cyc_st_3_3_2!=2'b10) | (~
      asn_itm_3) | (~ main_stage_0_4) | (rem_12cyc_st_3_1_0[0]);
  assign and_tmp_182 = or_753_cse & or_757_cse & or_tmp_733;
  assign nor_434_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_182));
  assign mux_276_nl = MUX_s_1_2_2(nor_434_nl, and_tmp_182, or_748_cse);
  assign and_dcpl_581 = mux_276_nl & and_dcpl_310 & and_dcpl_579;
  assign and_dcpl_582 = (rem_12cyc_st_5_3_2==2'b10);
  assign and_dcpl_583 = and_dcpl_582 & (~ (rem_12cyc_st_5_1_0[1]));
  assign or_762_cse = (rem_12cyc_st_4_1_0[1]) | (rem_12cyc_st_4_3_2!=2'b10) | (~
      asn_itm_4) | (~ main_stage_0_5) | (rem_12cyc_st_4_1_0[0]);
  assign and_tmp_185 = or_753_cse & or_757_cse & or_762_cse & or_tmp_733;
  assign nor_433_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_185));
  assign mux_277_nl = MUX_s_1_2_2(nor_433_nl, and_tmp_185, or_748_cse);
  assign and_dcpl_585 = mux_277_nl & and_dcpl_316 & and_dcpl_583;
  assign or_768_cse = (rem_12cyc_st_5_1_0[1]) | (rem_12cyc_st_5_3_2!=2'b10) | (~
      asn_itm_5) | (~ main_stage_0_6) | (rem_12cyc_st_5_1_0[0]);
  assign and_tmp_189 = or_753_cse & or_757_cse & or_762_cse & or_768_cse & or_tmp_733;
  assign nor_432_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_189));
  assign mux_278_nl = MUX_s_1_2_2(nor_432_nl, and_tmp_189, or_748_cse);
  assign and_dcpl_589 = mux_278_nl & and_dcpl_112 & and_dcpl_126 & (~ (rem_12cyc_st_6_1_0[1]));
  assign or_775_cse = (rem_12cyc_st_6_1_0!=2'b00) | (rem_12cyc_st_6_3_2!=2'b10);
  assign nor_430_nl = ~(and_dcpl_111 | (~ or_tmp_733));
  assign mux_279_nl = MUX_s_1_2_2(nor_430_nl, or_tmp_733, or_775_cse);
  assign and_tmp_193 = or_753_cse & or_757_cse & or_762_cse & or_768_cse & mux_279_nl;
  assign nor_431_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_193));
  assign mux_280_nl = MUX_s_1_2_2(nor_431_nl, and_tmp_193, or_748_cse);
  assign and_dcpl_593 = mux_280_nl & and_dcpl_85 & and_dcpl_99 & (~ (rem_12cyc_st_7_1_0[0]));
  assign or_784_cse = (rem_12cyc_st_7_1_0!=2'b00) | (rem_12cyc_st_7_3_2!=2'b10);
  assign nor_427_nl = ~(and_dcpl_84 | (~ or_tmp_733));
  assign mux_tmp_279 = MUX_s_1_2_2(nor_427_nl, or_tmp_733, or_784_cse);
  assign nor_428_nl = ~(and_dcpl_111 | (~ mux_tmp_279));
  assign mux_282_nl = MUX_s_1_2_2(nor_428_nl, mux_tmp_279, or_775_cse);
  assign and_tmp_197 = or_753_cse & or_757_cse & or_762_cse & or_768_cse & mux_282_nl;
  assign nor_429_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_197));
  assign mux_283_nl = MUX_s_1_2_2(nor_429_nl, and_tmp_197, or_748_cse);
  assign and_dcpl_597 = mux_283_nl & and_dcpl_58 & and_dcpl_72 & (~ (rem_12cyc_st_8_1_0[0]));
  assign or_795_cse = (rem_12cyc_st_8_1_0!=2'b00) | (rem_12cyc_st_8_3_2!=2'b10);
  assign nor_423_nl = ~(and_dcpl_57 | (~ or_tmp_733));
  assign mux_tmp_282 = MUX_s_1_2_2(nor_423_nl, or_tmp_733, or_795_cse);
  assign nor_424_nl = ~(and_dcpl_84 | (~ mux_tmp_282));
  assign mux_tmp_283 = MUX_s_1_2_2(nor_424_nl, mux_tmp_282, or_784_cse);
  assign nor_425_nl = ~(and_dcpl_111 | (~ mux_tmp_283));
  assign mux_286_nl = MUX_s_1_2_2(nor_425_nl, mux_tmp_283, or_775_cse);
  assign and_tmp_201 = or_753_cse & or_757_cse & or_762_cse & or_768_cse & mux_286_nl;
  assign nor_426_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_201));
  assign mux_287_nl = MUX_s_1_2_2(nor_426_nl, and_tmp_201, or_748_cse);
  assign and_dcpl_601 = mux_287_nl & and_dcpl_31 & and_dcpl_45 & (~ (rem_12cyc_st_9_1_0[0]));
  assign nor_418_nl = ~(and_dcpl_30 | (~ or_tmp_733));
  assign or_808_nl = (rem_12cyc_st_9_1_0!=2'b00) | (rem_12cyc_st_9_3_2!=2'b10);
  assign mux_tmp_286 = MUX_s_1_2_2(nor_418_nl, or_tmp_733, or_808_nl);
  assign nor_419_nl = ~(and_dcpl_57 | (~ mux_tmp_286));
  assign mux_tmp_287 = MUX_s_1_2_2(nor_419_nl, mux_tmp_286, or_795_cse);
  assign nor_420_nl = ~(and_dcpl_84 | (~ mux_tmp_287));
  assign mux_tmp_288 = MUX_s_1_2_2(nor_420_nl, mux_tmp_287, or_784_cse);
  assign nor_421_nl = ~(and_dcpl_111 | (~ mux_tmp_288));
  assign mux_291_nl = MUX_s_1_2_2(nor_421_nl, mux_tmp_288, or_775_cse);
  assign and_tmp_205 = or_753_cse & or_757_cse & or_762_cse & or_768_cse & mux_291_nl;
  assign nor_422_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_205));
  assign mux_292_nl = MUX_s_1_2_2(nor_422_nl, and_tmp_205, or_748_cse);
  assign and_dcpl_605 = mux_292_nl & and_dcpl_4 & and_dcpl_18 & (~ (rem_12cyc_st_10_1_0[0]));
  assign or_tmp_808 = (acc_tmp!=2'b10) | (acc_1_tmp[1:0]!=2'b00) | (~ ccs_ccore_start_rsci_idat);
  assign nor_409_nl = ~((rem_12cyc_st_10_3_2[1]) | (~ or_tmp_808));
  assign or_823_nl = (~ main_stage_0_11) | (~ asn_itm_10) | (rem_12cyc_st_10_1_0!=2'b00)
      | (rem_12cyc_st_10_3_2[0]);
  assign mux_tmp_291 = MUX_s_1_2_2(nor_409_nl, or_tmp_808, or_823_nl);
  assign nor_410_nl = ~((rem_12cyc_st_6_3_2[1]) | (~ mux_tmp_291));
  assign or_822_nl = (~ main_stage_0_7) | (~ asn_itm_6) | (rem_12cyc_st_6_1_0!=2'b00)
      | (rem_12cyc_st_6_3_2[0]);
  assign mux_tmp_292 = MUX_s_1_2_2(nor_410_nl, mux_tmp_291, or_822_nl);
  assign nor_411_nl = ~((rem_12cyc_st_5_3_2[1]) | (~ mux_tmp_292));
  assign or_821_nl = (~ main_stage_0_6) | (~ asn_itm_5) | (rem_12cyc_st_5_1_0!=2'b00)
      | (rem_12cyc_st_5_3_2[0]);
  assign mux_tmp_293 = MUX_s_1_2_2(nor_411_nl, mux_tmp_292, or_821_nl);
  assign nor_412_nl = ~((rem_12cyc_st_4_3_2[1]) | (~ mux_tmp_293));
  assign or_820_nl = (~ main_stage_0_5) | (~ asn_itm_4) | (rem_12cyc_st_4_1_0!=2'b00)
      | (rem_12cyc_st_4_3_2[0]);
  assign mux_tmp_294 = MUX_s_1_2_2(nor_412_nl, mux_tmp_293, or_820_nl);
  assign nor_413_nl = ~((rem_12cyc_st_3_3_2[1]) | (~ mux_tmp_294));
  assign or_819_nl = (~ main_stage_0_4) | (~ asn_itm_3) | (rem_12cyc_st_3_1_0!=2'b00)
      | (rem_12cyc_st_3_3_2[0]);
  assign mux_tmp_295 = MUX_s_1_2_2(nor_413_nl, mux_tmp_294, or_819_nl);
  assign nor_414_nl = ~((rem_12cyc_st_2_3_2[1]) | (~ mux_tmp_295));
  assign or_818_nl = (~ main_stage_0_3) | (~ asn_itm_2) | (rem_12cyc_st_2_1_0!=2'b00)
      | (rem_12cyc_st_2_3_2[0]);
  assign mux_tmp_296 = MUX_s_1_2_2(nor_414_nl, mux_tmp_295, or_818_nl);
  assign nor_415_nl = ~((rem_12cyc_st_9_3_2[1]) | (~ mux_tmp_296));
  assign or_817_nl = (~ main_stage_0_10) | (~ asn_itm_9) | (rem_12cyc_st_9_1_0!=2'b00)
      | (rem_12cyc_st_9_3_2[0]);
  assign mux_tmp_297 = MUX_s_1_2_2(nor_415_nl, mux_tmp_296, or_817_nl);
  assign nor_416_nl = ~((rem_12cyc_st_8_3_2[1]) | (~ mux_tmp_297));
  assign or_816_nl = (~ main_stage_0_9) | (~ asn_itm_8) | (rem_12cyc_st_8_1_0!=2'b00)
      | (rem_12cyc_st_8_3_2[0]);
  assign mux_tmp_298 = MUX_s_1_2_2(nor_416_nl, mux_tmp_297, or_816_nl);
  assign nor_417_nl = ~((rem_12cyc_st_7_3_2[1]) | (~ mux_tmp_298));
  assign or_815_nl = (~ main_stage_0_8) | (~ asn_itm_7) | (rem_12cyc_st_7_1_0!=2'b00)
      | (rem_12cyc_st_7_3_2[0]);
  assign mux_301_nl = MUX_s_1_2_2(nor_417_nl, mux_tmp_298, or_815_nl);
  assign and_tmp_206 = ((~ main_stage_0_2) | (~ asn_itm_1) | (rem_12cyc_3_2!=2'b10)
      | (rem_12cyc_1_0!=2'b00)) & mux_301_nl;
  assign and_dcpl_610 = and_dcpl_568 & and_dcpl_355;
  assign or_tmp_820 = (rem_12cyc_1_0!=2'b01) | (rem_12cyc_3_2!=2'b10) | not_tmp_54;
  assign or_837_cse = (acc_1_tmp[1:0]!=2'b01) | (acc_tmp!=2'b10);
  assign nor_408_nl = ~(ccs_ccore_start_rsci_idat | (~ or_tmp_820));
  assign mux_302_nl = MUX_s_1_2_2(nor_408_nl, or_tmp_820, or_837_cse);
  assign and_dcpl_612 = mux_302_nl & and_dcpl_358 & and_dcpl_571;
  assign nand_84_cse = ~((rem_12cyc_st_2_3_2[1]) & asn_itm_2 & main_stage_0_3 & (rem_12cyc_st_2_1_0[0]));
  assign or_842_cse = (rem_12cyc_st_2_1_0[1]) | (rem_12cyc_st_2_3_2[0]);
  assign and_986_nl = nand_84_cse & or_tmp_820;
  assign mux_tmp_301 = MUX_s_1_2_2(and_986_nl, or_tmp_820, or_842_cse);
  assign nor_407_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_301));
  assign mux_304_nl = MUX_s_1_2_2(nor_407_nl, mux_tmp_301, or_837_cse);
  assign and_dcpl_614 = mux_304_nl & and_dcpl_362 & and_dcpl_575;
  assign or_847_cse = (rem_12cyc_st_3_1_0[1]) | (rem_12cyc_st_3_3_2!=2'b10);
  assign and_984_nl = nand_274_cse & or_tmp_820;
  assign mux_tmp_303 = MUX_s_1_2_2(and_984_nl, or_tmp_820, or_847_cse);
  assign and_985_nl = nand_84_cse & mux_tmp_303;
  assign mux_tmp_304 = MUX_s_1_2_2(and_985_nl, mux_tmp_303, or_842_cse);
  assign nor_406_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_304));
  assign mux_307_nl = MUX_s_1_2_2(nor_406_nl, mux_tmp_304, or_837_cse);
  assign and_dcpl_616 = mux_307_nl & and_dcpl_366 & and_dcpl_579;
  assign nand_79_cse = ~((rem_12cyc_st_4_3_2[1]) & asn_itm_4 & main_stage_0_5 & (rem_12cyc_st_4_1_0[0]));
  assign or_854_cse = (rem_12cyc_st_4_1_0[1]) | (rem_12cyc_st_4_3_2[0]);
  assign and_981_nl = nand_79_cse & or_tmp_820;
  assign mux_tmp_306 = MUX_s_1_2_2(and_981_nl, or_tmp_820, or_854_cse);
  assign and_982_nl = nand_274_cse & mux_tmp_306;
  assign mux_tmp_307 = MUX_s_1_2_2(and_982_nl, mux_tmp_306, or_847_cse);
  assign and_983_nl = nand_84_cse & mux_tmp_307;
  assign mux_tmp_308 = MUX_s_1_2_2(and_983_nl, mux_tmp_307, or_842_cse);
  assign nor_405_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_308));
  assign mux_311_nl = MUX_s_1_2_2(nor_405_nl, mux_tmp_308, or_837_cse);
  assign and_dcpl_618 = mux_311_nl & and_dcpl_370 & and_dcpl_583;
  assign or_863_cse = (rem_12cyc_st_5_1_0[1]) | (rem_12cyc_st_5_3_2!=2'b10);
  assign and_977_nl = nand_267_cse & or_tmp_820;
  assign mux_tmp_310 = MUX_s_1_2_2(and_977_nl, or_tmp_820, or_863_cse);
  assign and_978_nl = nand_79_cse & mux_tmp_310;
  assign mux_tmp_311 = MUX_s_1_2_2(and_978_nl, mux_tmp_310, or_854_cse);
  assign and_979_nl = nand_274_cse & mux_tmp_311;
  assign mux_tmp_312 = MUX_s_1_2_2(and_979_nl, mux_tmp_311, or_847_cse);
  assign and_980_nl = nand_84_cse & mux_tmp_312;
  assign mux_tmp_313 = MUX_s_1_2_2(and_980_nl, mux_tmp_312, or_842_cse);
  assign nor_404_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_313));
  assign mux_316_nl = MUX_s_1_2_2(nor_404_nl, mux_tmp_313, or_837_cse);
  assign and_dcpl_622 = mux_316_nl & and_dcpl_112 & and_dcpl_129 & (~ (rem_12cyc_st_6_1_0[1]));
  assign or_874_cse = (rem_12cyc_st_6_1_0!=2'b01) | (rem_12cyc_st_6_3_2!=2'b10);
  assign nor_402_nl = ~(and_dcpl_111 | (~ or_tmp_820));
  assign mux_tmp_315 = MUX_s_1_2_2(nor_402_nl, or_tmp_820, or_874_cse);
  assign and_973_nl = nand_267_cse & mux_tmp_315;
  assign mux_tmp_316 = MUX_s_1_2_2(and_973_nl, mux_tmp_315, or_863_cse);
  assign and_974_nl = nand_79_cse & mux_tmp_316;
  assign mux_tmp_317 = MUX_s_1_2_2(and_974_nl, mux_tmp_316, or_854_cse);
  assign and_975_nl = nand_274_cse & mux_tmp_317;
  assign mux_tmp_318 = MUX_s_1_2_2(and_975_nl, mux_tmp_317, or_847_cse);
  assign and_976_nl = nand_84_cse & mux_tmp_318;
  assign mux_tmp_319 = MUX_s_1_2_2(and_976_nl, mux_tmp_318, or_842_cse);
  assign nor_403_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_319));
  assign mux_322_nl = MUX_s_1_2_2(nor_403_nl, mux_tmp_319, or_837_cse);
  assign and_dcpl_625 = mux_322_nl & and_dcpl_85 & and_dcpl_99 & (rem_12cyc_st_7_1_0[0]);
  assign or_887_cse = (rem_12cyc_st_7_1_0!=2'b01) | (rem_12cyc_st_7_3_2!=2'b10);
  assign nor_399_nl = ~(and_dcpl_84 | (~ or_tmp_820));
  assign mux_tmp_321 = MUX_s_1_2_2(nor_399_nl, or_tmp_820, or_887_cse);
  assign nor_400_nl = ~(and_dcpl_111 | (~ mux_tmp_321));
  assign mux_tmp_322 = MUX_s_1_2_2(nor_400_nl, mux_tmp_321, or_874_cse);
  assign and_969_nl = nand_267_cse & mux_tmp_322;
  assign mux_tmp_323 = MUX_s_1_2_2(and_969_nl, mux_tmp_322, or_863_cse);
  assign and_970_nl = nand_79_cse & mux_tmp_323;
  assign mux_tmp_324 = MUX_s_1_2_2(and_970_nl, mux_tmp_323, or_854_cse);
  assign and_971_nl = nand_274_cse & mux_tmp_324;
  assign mux_tmp_325 = MUX_s_1_2_2(and_971_nl, mux_tmp_324, or_847_cse);
  assign and_972_nl = nand_84_cse & mux_tmp_325;
  assign mux_tmp_326 = MUX_s_1_2_2(and_972_nl, mux_tmp_325, or_842_cse);
  assign nor_401_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_326));
  assign mux_329_nl = MUX_s_1_2_2(nor_401_nl, mux_tmp_326, or_837_cse);
  assign and_dcpl_628 = mux_329_nl & and_dcpl_58 & and_dcpl_72 & (rem_12cyc_st_8_1_0[0]);
  assign or_902_cse = (rem_12cyc_st_8_1_0!=2'b01) | (rem_12cyc_st_8_3_2!=2'b10);
  assign nor_395_nl = ~(and_dcpl_57 | (~ or_tmp_820));
  assign mux_tmp_328 = MUX_s_1_2_2(nor_395_nl, or_tmp_820, or_902_cse);
  assign nor_396_nl = ~(and_dcpl_84 | (~ mux_tmp_328));
  assign mux_tmp_329 = MUX_s_1_2_2(nor_396_nl, mux_tmp_328, or_887_cse);
  assign nor_397_nl = ~(and_dcpl_111 | (~ mux_tmp_329));
  assign mux_tmp_330 = MUX_s_1_2_2(nor_397_nl, mux_tmp_329, or_874_cse);
  assign and_965_nl = nand_267_cse & mux_tmp_330;
  assign mux_tmp_331 = MUX_s_1_2_2(and_965_nl, mux_tmp_330, or_863_cse);
  assign and_966_nl = nand_79_cse & mux_tmp_331;
  assign mux_tmp_332 = MUX_s_1_2_2(and_966_nl, mux_tmp_331, or_854_cse);
  assign and_967_nl = nand_274_cse & mux_tmp_332;
  assign mux_tmp_333 = MUX_s_1_2_2(and_967_nl, mux_tmp_332, or_847_cse);
  assign and_968_nl = nand_84_cse & mux_tmp_333;
  assign mux_tmp_334 = MUX_s_1_2_2(and_968_nl, mux_tmp_333, or_842_cse);
  assign nor_398_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_334));
  assign mux_337_nl = MUX_s_1_2_2(nor_398_nl, mux_tmp_334, or_837_cse);
  assign and_dcpl_631 = mux_337_nl & and_dcpl_31 & and_dcpl_45 & (rem_12cyc_st_9_1_0[0]);
  assign nor_390_nl = ~(and_dcpl_30 | (~ or_tmp_820));
  assign or_919_nl = (rem_12cyc_st_9_1_0!=2'b01) | (rem_12cyc_st_9_3_2!=2'b10);
  assign mux_tmp_336 = MUX_s_1_2_2(nor_390_nl, or_tmp_820, or_919_nl);
  assign nor_391_nl = ~(and_dcpl_57 | (~ mux_tmp_336));
  assign mux_tmp_337 = MUX_s_1_2_2(nor_391_nl, mux_tmp_336, or_902_cse);
  assign nor_392_nl = ~(and_dcpl_84 | (~ mux_tmp_337));
  assign mux_tmp_338 = MUX_s_1_2_2(nor_392_nl, mux_tmp_337, or_887_cse);
  assign nor_393_nl = ~(and_dcpl_111 | (~ mux_tmp_338));
  assign mux_tmp_339 = MUX_s_1_2_2(nor_393_nl, mux_tmp_338, or_874_cse);
  assign and_961_nl = nand_267_cse & mux_tmp_339;
  assign mux_tmp_340 = MUX_s_1_2_2(and_961_nl, mux_tmp_339, or_863_cse);
  assign and_962_nl = nand_79_cse & mux_tmp_340;
  assign mux_tmp_341 = MUX_s_1_2_2(and_962_nl, mux_tmp_340, or_854_cse);
  assign and_963_nl = nand_274_cse & mux_tmp_341;
  assign mux_tmp_342 = MUX_s_1_2_2(and_963_nl, mux_tmp_341, or_847_cse);
  assign and_964_nl = nand_84_cse & mux_tmp_342;
  assign mux_tmp_343 = MUX_s_1_2_2(and_964_nl, mux_tmp_342, or_842_cse);
  assign nor_394_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_343));
  assign mux_346_nl = MUX_s_1_2_2(nor_394_nl, mux_tmp_343, or_837_cse);
  assign and_dcpl_634 = mux_346_nl & and_dcpl_4 & and_dcpl_18 & (rem_12cyc_st_10_1_0[0]);
  assign or_tmp_921 = (acc_tmp!=2'b10) | (acc_1_tmp[1]) | nand_250_cse;
  assign nor_380_nl = ~((rem_12cyc_st_10_3_2[1]) | (~ or_tmp_921));
  assign or_938_nl = (~ main_stage_0_11) | (~ asn_itm_10) | (rem_12cyc_st_10_1_0!=2'b01)
      | (rem_12cyc_st_10_3_2[0]);
  assign mux_tmp_345 = MUX_s_1_2_2(nor_380_nl, or_tmp_921, or_938_nl);
  assign nor_381_nl = ~((rem_12cyc_st_6_3_2[1]) | (~ mux_tmp_345));
  assign or_937_nl = (~ main_stage_0_7) | (~ asn_itm_6) | (rem_12cyc_st_6_1_0!=2'b01)
      | (rem_12cyc_st_6_3_2[0]);
  assign mux_tmp_346 = MUX_s_1_2_2(nor_381_nl, mux_tmp_345, or_937_nl);
  assign nor_382_nl = ~((rem_12cyc_st_5_3_2[1]) | (~ mux_tmp_346));
  assign or_936_nl = (~ main_stage_0_6) | (~ asn_itm_5) | (rem_12cyc_st_5_1_0!=2'b01)
      | (rem_12cyc_st_5_3_2[0]);
  assign mux_tmp_347 = MUX_s_1_2_2(nor_382_nl, mux_tmp_346, or_936_nl);
  assign nor_383_nl = ~((rem_12cyc_st_4_3_2[1]) | (~ mux_tmp_347));
  assign or_935_nl = (~ main_stage_0_5) | (~ asn_itm_4) | (rem_12cyc_st_4_1_0!=2'b01)
      | (rem_12cyc_st_4_3_2[0]);
  assign mux_tmp_348 = MUX_s_1_2_2(nor_383_nl, mux_tmp_347, or_935_nl);
  assign nor_384_nl = ~((rem_12cyc_st_3_3_2[1]) | (~ mux_tmp_348));
  assign or_934_nl = (~ main_stage_0_4) | (~ asn_itm_3) | (rem_12cyc_st_3_1_0!=2'b01)
      | (rem_12cyc_st_3_3_2[0]);
  assign mux_tmp_349 = MUX_s_1_2_2(nor_384_nl, mux_tmp_348, or_934_nl);
  assign nor_385_nl = ~((rem_12cyc_st_2_3_2[1]) | (~ mux_tmp_349));
  assign or_933_nl = (~ main_stage_0_3) | (~ asn_itm_2) | (rem_12cyc_st_2_1_0!=2'b01)
      | (rem_12cyc_st_2_3_2[0]);
  assign mux_tmp_350 = MUX_s_1_2_2(nor_385_nl, mux_tmp_349, or_933_nl);
  assign nor_386_nl = ~((rem_12cyc_st_9_3_2[1]) | (~ mux_tmp_350));
  assign or_932_nl = (~ main_stage_0_10) | (~ asn_itm_9) | (rem_12cyc_st_9_1_0!=2'b01)
      | (rem_12cyc_st_9_3_2[0]);
  assign mux_tmp_351 = MUX_s_1_2_2(nor_386_nl, mux_tmp_350, or_932_nl);
  assign nor_387_nl = ~((rem_12cyc_st_8_3_2[1]) | (~ mux_tmp_351));
  assign or_931_nl = (~ main_stage_0_9) | (~ asn_itm_8) | (rem_12cyc_st_8_1_0!=2'b01)
      | (rem_12cyc_st_8_3_2[0]);
  assign mux_tmp_352 = MUX_s_1_2_2(nor_387_nl, mux_tmp_351, or_931_nl);
  assign nor_388_nl = ~((rem_12cyc_st_7_3_2[1]) | (~ mux_tmp_352));
  assign or_930_nl = (~ main_stage_0_8) | (~ asn_itm_7) | (rem_12cyc_st_7_1_0!=2'b01)
      | (rem_12cyc_st_7_3_2[0]);
  assign mux_tmp_353 = MUX_s_1_2_2(nor_388_nl, mux_tmp_352, or_930_nl);
  assign nor_389_nl = ~((rem_12cyc_1_0[0]) | (~ mux_tmp_353));
  assign or_929_nl = (~ main_stage_0_2) | (~ asn_itm_1) | (rem_12cyc_3_2!=2'b10)
      | (rem_12cyc_1_0[1]);
  assign mux_tmp_354 = MUX_s_1_2_2(nor_389_nl, mux_tmp_353, or_929_nl);
  assign and_dcpl_638 = and_dcpl_568 & and_dcpl_393;
  assign and_dcpl_639 = and_dcpl_570 & (rem_12cyc_st_2_1_0[1]);
  assign or_tmp_934 = (rem_12cyc_1_0!=2'b10) | (rem_12cyc_3_2!=2'b10) | not_tmp_54;
  assign or_952_cse = (acc_1_tmp[1:0]!=2'b10) | (acc_tmp!=2'b10);
  assign nor_379_nl = ~(ccs_ccore_start_rsci_idat | (~ or_tmp_934));
  assign mux_357_nl = MUX_s_1_2_2(nor_379_nl, or_tmp_934, or_952_cse);
  assign and_dcpl_641 = mux_357_nl & and_dcpl_298 & and_dcpl_639;
  assign and_dcpl_642 = and_dcpl_574 & (rem_12cyc_st_3_1_0[1]);
  assign or_957_cse = (~ (rem_12cyc_st_2_1_0[1])) | (rem_12cyc_st_2_3_2!=2'b10) |
      (~ asn_itm_2) | (~ main_stage_0_3) | (rem_12cyc_st_2_1_0[0]);
  assign and_tmp_207 = or_957_cse & or_tmp_934;
  assign nor_378_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_207));
  assign mux_358_nl = MUX_s_1_2_2(nor_378_nl, and_tmp_207, or_952_cse);
  assign and_dcpl_644 = mux_358_nl & and_dcpl_304 & and_dcpl_642;
  assign and_dcpl_645 = and_dcpl_578 & (rem_12cyc_st_4_1_0[1]);
  assign or_961_cse = (~ (rem_12cyc_st_3_1_0[1])) | (rem_12cyc_st_3_3_2!=2'b10) |
      (~ asn_itm_3) | (~ main_stage_0_4) | (rem_12cyc_st_3_1_0[0]);
  assign and_tmp_209 = or_957_cse & or_961_cse & or_tmp_934;
  assign nor_377_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_209));
  assign mux_359_nl = MUX_s_1_2_2(nor_377_nl, and_tmp_209, or_952_cse);
  assign and_dcpl_647 = mux_359_nl & and_dcpl_310 & and_dcpl_645;
  assign and_dcpl_648 = and_dcpl_582 & (rem_12cyc_st_5_1_0[1]);
  assign or_966_cse = (~ (rem_12cyc_st_4_1_0[1])) | (rem_12cyc_st_4_3_2!=2'b10) |
      (~ asn_itm_4) | (~ main_stage_0_5) | (rem_12cyc_st_4_1_0[0]);
  assign and_tmp_212 = or_957_cse & or_961_cse & or_966_cse & or_tmp_934;
  assign nor_376_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_212));
  assign mux_360_nl = MUX_s_1_2_2(nor_376_nl, and_tmp_212, or_952_cse);
  assign and_dcpl_650 = mux_360_nl & and_dcpl_316 & and_dcpl_648;
  assign or_972_cse = (~ (rem_12cyc_st_5_1_0[1])) | (rem_12cyc_st_5_3_2!=2'b10) |
      (~ asn_itm_5) | (~ main_stage_0_6) | (rem_12cyc_st_5_1_0[0]);
  assign and_tmp_216 = or_957_cse & or_961_cse & or_966_cse & or_972_cse & or_tmp_934;
  assign nor_375_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_216));
  assign mux_361_nl = MUX_s_1_2_2(nor_375_nl, and_tmp_216, or_952_cse);
  assign and_dcpl_653 = mux_361_nl & and_dcpl_112 & and_dcpl_126 & (rem_12cyc_st_6_1_0[1]);
  assign or_979_cse = (rem_12cyc_st_6_1_0!=2'b10) | (rem_12cyc_st_6_3_2!=2'b10);
  assign nor_373_nl = ~(and_dcpl_111 | (~ or_tmp_934));
  assign mux_362_nl = MUX_s_1_2_2(nor_373_nl, or_tmp_934, or_979_cse);
  assign and_tmp_220 = or_957_cse & or_961_cse & or_966_cse & or_972_cse & mux_362_nl;
  assign nor_374_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_220));
  assign mux_363_nl = MUX_s_1_2_2(nor_374_nl, and_tmp_220, or_952_cse);
  assign and_dcpl_657 = mux_363_nl & and_dcpl_85 & and_dcpl_104 & (~ (rem_12cyc_st_7_1_0[0]));
  assign or_988_cse = (rem_12cyc_st_7_1_0!=2'b10) | (rem_12cyc_st_7_3_2!=2'b10);
  assign nor_370_nl = ~(and_dcpl_84 | (~ or_tmp_934));
  assign mux_tmp_362 = MUX_s_1_2_2(nor_370_nl, or_tmp_934, or_988_cse);
  assign nor_371_nl = ~(and_dcpl_111 | (~ mux_tmp_362));
  assign mux_365_nl = MUX_s_1_2_2(nor_371_nl, mux_tmp_362, or_979_cse);
  assign and_tmp_224 = or_957_cse & or_961_cse & or_966_cse & or_972_cse & mux_365_nl;
  assign nor_372_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_224));
  assign mux_366_nl = MUX_s_1_2_2(nor_372_nl, and_tmp_224, or_952_cse);
  assign and_dcpl_661 = mux_366_nl & and_dcpl_58 & and_dcpl_77 & (~ (rem_12cyc_st_8_1_0[0]));
  assign or_999_cse = (rem_12cyc_st_8_1_0!=2'b10) | (rem_12cyc_st_8_3_2!=2'b10);
  assign nor_366_nl = ~(and_dcpl_57 | (~ or_tmp_934));
  assign mux_tmp_365 = MUX_s_1_2_2(nor_366_nl, or_tmp_934, or_999_cse);
  assign nor_367_nl = ~(and_dcpl_84 | (~ mux_tmp_365));
  assign mux_tmp_366 = MUX_s_1_2_2(nor_367_nl, mux_tmp_365, or_988_cse);
  assign nor_368_nl = ~(and_dcpl_111 | (~ mux_tmp_366));
  assign mux_369_nl = MUX_s_1_2_2(nor_368_nl, mux_tmp_366, or_979_cse);
  assign and_tmp_228 = or_957_cse & or_961_cse & or_966_cse & or_972_cse & mux_369_nl;
  assign nor_369_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_228));
  assign mux_370_nl = MUX_s_1_2_2(nor_369_nl, and_tmp_228, or_952_cse);
  assign and_dcpl_665 = mux_370_nl & and_dcpl_31 & and_dcpl_50 & (~ (rem_12cyc_st_9_1_0[0]));
  assign nor_361_nl = ~(and_dcpl_30 | (~ or_tmp_934));
  assign or_1012_nl = (rem_12cyc_st_9_1_0!=2'b10) | (rem_12cyc_st_9_3_2!=2'b10);
  assign mux_tmp_369 = MUX_s_1_2_2(nor_361_nl, or_tmp_934, or_1012_nl);
  assign nor_362_nl = ~(and_dcpl_57 | (~ mux_tmp_369));
  assign mux_tmp_370 = MUX_s_1_2_2(nor_362_nl, mux_tmp_369, or_999_cse);
  assign nor_363_nl = ~(and_dcpl_84 | (~ mux_tmp_370));
  assign mux_tmp_371 = MUX_s_1_2_2(nor_363_nl, mux_tmp_370, or_988_cse);
  assign nor_364_nl = ~(and_dcpl_111 | (~ mux_tmp_371));
  assign mux_374_nl = MUX_s_1_2_2(nor_364_nl, mux_tmp_371, or_979_cse);
  assign and_tmp_232 = or_957_cse & or_961_cse & or_966_cse & or_972_cse & mux_374_nl;
  assign nor_365_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_232));
  assign mux_375_nl = MUX_s_1_2_2(nor_365_nl, and_tmp_232, or_952_cse);
  assign and_dcpl_669 = mux_375_nl & and_dcpl_4 & and_dcpl_23 & (~ (rem_12cyc_st_10_1_0[0]));
  assign or_tmp_1009 = (acc_tmp!=2'b10) | (acc_1_tmp[1:0]!=2'b10) | (~ ccs_ccore_start_rsci_idat);
  assign nor_352_nl = ~((rem_12cyc_st_10_3_2[1]) | (~ or_tmp_1009));
  assign or_1027_nl = (~ main_stage_0_11) | (~ asn_itm_10) | (rem_12cyc_st_10_1_0!=2'b10)
      | (rem_12cyc_st_10_3_2[0]);
  assign mux_tmp_374 = MUX_s_1_2_2(nor_352_nl, or_tmp_1009, or_1027_nl);
  assign nor_353_nl = ~((rem_12cyc_st_6_3_2[1]) | (~ mux_tmp_374));
  assign or_1026_nl = (~ main_stage_0_7) | (~ asn_itm_6) | (rem_12cyc_st_6_1_0!=2'b10)
      | (rem_12cyc_st_6_3_2[0]);
  assign mux_tmp_375 = MUX_s_1_2_2(nor_353_nl, mux_tmp_374, or_1026_nl);
  assign nor_354_nl = ~((rem_12cyc_st_5_3_2[1]) | (~ mux_tmp_375));
  assign or_1025_nl = (~ main_stage_0_6) | (~ asn_itm_5) | (rem_12cyc_st_5_1_0!=2'b10)
      | (rem_12cyc_st_5_3_2[0]);
  assign mux_tmp_376 = MUX_s_1_2_2(nor_354_nl, mux_tmp_375, or_1025_nl);
  assign nor_355_nl = ~((rem_12cyc_st_4_3_2[1]) | (~ mux_tmp_376));
  assign or_1024_nl = (~ main_stage_0_5) | (~ asn_itm_4) | (rem_12cyc_st_4_1_0!=2'b10)
      | (rem_12cyc_st_4_3_2[0]);
  assign mux_tmp_377 = MUX_s_1_2_2(nor_355_nl, mux_tmp_376, or_1024_nl);
  assign nor_356_nl = ~((rem_12cyc_st_3_3_2[1]) | (~ mux_tmp_377));
  assign or_1023_nl = (~ main_stage_0_4) | (~ asn_itm_3) | (rem_12cyc_st_3_1_0!=2'b10)
      | (rem_12cyc_st_3_3_2[0]);
  assign mux_tmp_378 = MUX_s_1_2_2(nor_356_nl, mux_tmp_377, or_1023_nl);
  assign nor_357_nl = ~((rem_12cyc_st_2_3_2[1]) | (~ mux_tmp_378));
  assign or_1022_nl = (~ main_stage_0_3) | (~ asn_itm_2) | (rem_12cyc_st_2_1_0!=2'b10)
      | (rem_12cyc_st_2_3_2[0]);
  assign mux_tmp_379 = MUX_s_1_2_2(nor_357_nl, mux_tmp_378, or_1022_nl);
  assign nor_358_nl = ~((rem_12cyc_st_9_3_2[1]) | (~ mux_tmp_379));
  assign or_1021_nl = (~ main_stage_0_10) | (~ asn_itm_9) | (rem_12cyc_st_9_1_0!=2'b10)
      | (rem_12cyc_st_9_3_2[0]);
  assign mux_tmp_380 = MUX_s_1_2_2(nor_358_nl, mux_tmp_379, or_1021_nl);
  assign nor_359_nl = ~((rem_12cyc_st_8_3_2[1]) | (~ mux_tmp_380));
  assign or_1020_nl = (~ main_stage_0_9) | (~ asn_itm_8) | (rem_12cyc_st_8_1_0!=2'b10)
      | (rem_12cyc_st_8_3_2[0]);
  assign mux_tmp_381 = MUX_s_1_2_2(nor_359_nl, mux_tmp_380, or_1020_nl);
  assign nor_360_nl = ~((rem_12cyc_st_7_3_2[1]) | (~ mux_tmp_381));
  assign or_1019_nl = (~ main_stage_0_8) | (~ asn_itm_7) | (rem_12cyc_st_7_1_0!=2'b10)
      | (rem_12cyc_st_7_3_2[0]);
  assign mux_384_nl = MUX_s_1_2_2(nor_360_nl, mux_tmp_381, or_1019_nl);
  assign and_tmp_233 = ((~ main_stage_0_2) | (~ asn_itm_1) | (rem_12cyc_3_2!=2'b10)
      | (rem_12cyc_1_0!=2'b10)) & mux_384_nl;
  assign and_dcpl_673 = and_dcpl_568 & and_dcpl_430;
  assign or_tmp_1021 = (~((rem_12cyc_1_0==2'b11) & (rem_12cyc_3_2==2'b10))) | not_tmp_54;
  assign nand_57_cse = ~((acc_1_tmp[1:0]==2'b11) & (acc_tmp==2'b10));
  assign nor_351_nl = ~(ccs_ccore_start_rsci_idat | (~ or_tmp_1021));
  assign mux_385_nl = MUX_s_1_2_2(nor_351_nl, or_tmp_1021, nand_57_cse);
  assign and_dcpl_675 = mux_385_nl & and_dcpl_358 & and_dcpl_639;
  assign or_1045_cse = (~ (rem_12cyc_st_2_1_0[1])) | (rem_12cyc_st_2_3_2[0]);
  assign and_960_nl = nand_84_cse & or_tmp_1021;
  assign mux_tmp_384 = MUX_s_1_2_2(and_960_nl, or_tmp_1021, or_1045_cse);
  assign nor_350_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_384));
  assign mux_387_nl = MUX_s_1_2_2(nor_350_nl, mux_tmp_384, nand_57_cse);
  assign and_dcpl_677 = mux_387_nl & and_dcpl_362 & and_dcpl_642;
  assign or_1050_cse = (~ (rem_12cyc_st_3_1_0[1])) | (rem_12cyc_st_3_3_2!=2'b10);
  assign and_958_nl = nand_274_cse & or_tmp_1021;
  assign mux_tmp_386 = MUX_s_1_2_2(and_958_nl, or_tmp_1021, or_1050_cse);
  assign and_959_nl = nand_84_cse & mux_tmp_386;
  assign mux_tmp_387 = MUX_s_1_2_2(and_959_nl, mux_tmp_386, or_1045_cse);
  assign nor_349_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_387));
  assign mux_390_nl = MUX_s_1_2_2(nor_349_nl, mux_tmp_387, nand_57_cse);
  assign and_dcpl_679 = mux_390_nl & and_dcpl_366 & and_dcpl_645;
  assign or_1057_cse = (~ (rem_12cyc_st_4_1_0[1])) | (rem_12cyc_st_4_3_2[0]);
  assign and_955_nl = nand_79_cse & or_tmp_1021;
  assign mux_tmp_389 = MUX_s_1_2_2(and_955_nl, or_tmp_1021, or_1057_cse);
  assign and_956_nl = nand_274_cse & mux_tmp_389;
  assign mux_tmp_390 = MUX_s_1_2_2(and_956_nl, mux_tmp_389, or_1050_cse);
  assign and_957_nl = nand_84_cse & mux_tmp_390;
  assign mux_tmp_391 = MUX_s_1_2_2(and_957_nl, mux_tmp_390, or_1045_cse);
  assign nor_348_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_391));
  assign mux_394_nl = MUX_s_1_2_2(nor_348_nl, mux_tmp_391, nand_57_cse);
  assign and_dcpl_681 = mux_394_nl & and_dcpl_370 & and_dcpl_648;
  assign or_1066_cse = (~ (rem_12cyc_st_5_1_0[1])) | (rem_12cyc_st_5_3_2!=2'b10);
  assign and_951_nl = nand_267_cse & or_tmp_1021;
  assign mux_tmp_393 = MUX_s_1_2_2(and_951_nl, or_tmp_1021, or_1066_cse);
  assign and_952_nl = nand_79_cse & mux_tmp_393;
  assign mux_tmp_394 = MUX_s_1_2_2(and_952_nl, mux_tmp_393, or_1057_cse);
  assign and_953_nl = nand_274_cse & mux_tmp_394;
  assign mux_tmp_395 = MUX_s_1_2_2(and_953_nl, mux_tmp_394, or_1050_cse);
  assign and_954_nl = nand_84_cse & mux_tmp_395;
  assign mux_tmp_396 = MUX_s_1_2_2(and_954_nl, mux_tmp_395, or_1045_cse);
  assign nor_347_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_396));
  assign mux_399_nl = MUX_s_1_2_2(nor_347_nl, mux_tmp_396, nand_57_cse);
  assign and_dcpl_684 = mux_399_nl & and_dcpl_112 & and_dcpl_129 & (rem_12cyc_st_6_1_0[1]);
  assign nand_36_cse = ~((rem_12cyc_st_6_1_0==2'b11) & (rem_12cyc_st_6_3_2==2'b10));
  assign nor_345_nl = ~(and_dcpl_111 | (~ or_tmp_1021));
  assign mux_tmp_398 = MUX_s_1_2_2(nor_345_nl, or_tmp_1021, nand_36_cse);
  assign and_947_nl = nand_267_cse & mux_tmp_398;
  assign mux_tmp_399 = MUX_s_1_2_2(and_947_nl, mux_tmp_398, or_1066_cse);
  assign and_948_nl = nand_79_cse & mux_tmp_399;
  assign mux_tmp_400 = MUX_s_1_2_2(and_948_nl, mux_tmp_399, or_1057_cse);
  assign and_949_nl = nand_274_cse & mux_tmp_400;
  assign mux_tmp_401 = MUX_s_1_2_2(and_949_nl, mux_tmp_400, or_1050_cse);
  assign and_950_nl = nand_84_cse & mux_tmp_401;
  assign mux_tmp_402 = MUX_s_1_2_2(and_950_nl, mux_tmp_401, or_1045_cse);
  assign nor_346_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_402));
  assign mux_405_nl = MUX_s_1_2_2(nor_346_nl, mux_tmp_402, nand_57_cse);
  assign and_dcpl_687 = mux_405_nl & and_dcpl_85 & and_dcpl_104 & (rem_12cyc_st_7_1_0[0]);
  assign nand_29_cse = ~((rem_12cyc_st_7_1_0==2'b11) & (rem_12cyc_st_7_3_2==2'b10));
  assign nor_342_nl = ~(and_dcpl_84 | (~ or_tmp_1021));
  assign mux_tmp_404 = MUX_s_1_2_2(nor_342_nl, or_tmp_1021, nand_29_cse);
  assign nor_343_nl = ~(and_dcpl_111 | (~ mux_tmp_404));
  assign mux_tmp_405 = MUX_s_1_2_2(nor_343_nl, mux_tmp_404, nand_36_cse);
  assign and_943_nl = nand_267_cse & mux_tmp_405;
  assign mux_tmp_406 = MUX_s_1_2_2(and_943_nl, mux_tmp_405, or_1066_cse);
  assign and_944_nl = nand_79_cse & mux_tmp_406;
  assign mux_tmp_407 = MUX_s_1_2_2(and_944_nl, mux_tmp_406, or_1057_cse);
  assign and_945_nl = nand_274_cse & mux_tmp_407;
  assign mux_tmp_408 = MUX_s_1_2_2(and_945_nl, mux_tmp_407, or_1050_cse);
  assign and_946_nl = nand_84_cse & mux_tmp_408;
  assign mux_tmp_409 = MUX_s_1_2_2(and_946_nl, mux_tmp_408, or_1045_cse);
  assign nor_344_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_409));
  assign mux_412_nl = MUX_s_1_2_2(nor_344_nl, mux_tmp_409, nand_57_cse);
  assign and_dcpl_690 = mux_412_nl & and_dcpl_58 & and_dcpl_77 & (rem_12cyc_st_8_1_0[0]);
  assign nand_21_cse = ~((rem_12cyc_st_8_1_0==2'b11) & (rem_12cyc_st_8_3_2==2'b10));
  assign nor_338_nl = ~(and_dcpl_57 | (~ or_tmp_1021));
  assign mux_tmp_411 = MUX_s_1_2_2(nor_338_nl, or_tmp_1021, nand_21_cse);
  assign nor_339_nl = ~(and_dcpl_84 | (~ mux_tmp_411));
  assign mux_tmp_412 = MUX_s_1_2_2(nor_339_nl, mux_tmp_411, nand_29_cse);
  assign nor_340_nl = ~(and_dcpl_111 | (~ mux_tmp_412));
  assign mux_tmp_413 = MUX_s_1_2_2(nor_340_nl, mux_tmp_412, nand_36_cse);
  assign and_939_nl = nand_267_cse & mux_tmp_413;
  assign mux_tmp_414 = MUX_s_1_2_2(and_939_nl, mux_tmp_413, or_1066_cse);
  assign and_940_nl = nand_79_cse & mux_tmp_414;
  assign mux_tmp_415 = MUX_s_1_2_2(and_940_nl, mux_tmp_414, or_1057_cse);
  assign and_941_nl = nand_274_cse & mux_tmp_415;
  assign mux_tmp_416 = MUX_s_1_2_2(and_941_nl, mux_tmp_415, or_1050_cse);
  assign and_942_nl = nand_84_cse & mux_tmp_416;
  assign mux_tmp_417 = MUX_s_1_2_2(and_942_nl, mux_tmp_416, or_1045_cse);
  assign nor_341_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_417));
  assign mux_420_nl = MUX_s_1_2_2(nor_341_nl, mux_tmp_417, nand_57_cse);
  assign and_dcpl_693 = mux_420_nl & and_dcpl_31 & and_dcpl_50 & (rem_12cyc_st_9_1_0[0]);
  assign nor_333_nl = ~(and_dcpl_30 | (~ or_tmp_1021));
  assign nand_12_nl = ~((rem_12cyc_st_9_1_0==2'b11) & (rem_12cyc_st_9_3_2==2'b10));
  assign mux_tmp_419 = MUX_s_1_2_2(nor_333_nl, or_tmp_1021, nand_12_nl);
  assign nor_334_nl = ~(and_dcpl_57 | (~ mux_tmp_419));
  assign mux_tmp_420 = MUX_s_1_2_2(nor_334_nl, mux_tmp_419, nand_21_cse);
  assign nor_335_nl = ~(and_dcpl_84 | (~ mux_tmp_420));
  assign mux_tmp_421 = MUX_s_1_2_2(nor_335_nl, mux_tmp_420, nand_29_cse);
  assign nor_336_nl = ~(and_dcpl_111 | (~ mux_tmp_421));
  assign mux_tmp_422 = MUX_s_1_2_2(nor_336_nl, mux_tmp_421, nand_36_cse);
  assign and_935_nl = nand_267_cse & mux_tmp_422;
  assign mux_tmp_423 = MUX_s_1_2_2(and_935_nl, mux_tmp_422, or_1066_cse);
  assign and_936_nl = nand_79_cse & mux_tmp_423;
  assign mux_tmp_424 = MUX_s_1_2_2(and_936_nl, mux_tmp_423, or_1057_cse);
  assign and_937_nl = nand_274_cse & mux_tmp_424;
  assign mux_tmp_425 = MUX_s_1_2_2(and_937_nl, mux_tmp_424, or_1050_cse);
  assign and_938_nl = nand_84_cse & mux_tmp_425;
  assign mux_tmp_426 = MUX_s_1_2_2(and_938_nl, mux_tmp_425, or_1045_cse);
  assign nor_337_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_426));
  assign mux_429_nl = MUX_s_1_2_2(nor_337_nl, mux_tmp_426, nand_57_cse);
  assign and_dcpl_696 = mux_429_nl & and_dcpl_4 & and_dcpl_23 & (rem_12cyc_st_10_1_0[0]);
  assign or_tmp_1122 = (acc_tmp!=2'b10) | nand_222_cse;
  assign nor_324_nl = ~((rem_12cyc_st_10_3_2[1]) | (~ or_tmp_1122));
  assign nand_1_nl = ~(main_stage_0_11 & asn_itm_10 & (rem_12cyc_st_10_1_0==2'b11)
      & (~ (rem_12cyc_st_10_3_2[0])));
  assign mux_tmp_428 = MUX_s_1_2_2(nor_324_nl, or_tmp_1122, nand_1_nl);
  assign nor_325_nl = ~((rem_12cyc_st_6_3_2[1]) | (~ mux_tmp_428));
  assign nand_2_nl = ~(main_stage_0_7 & asn_itm_6 & (rem_12cyc_st_6_1_0==2'b11) &
      (~ (rem_12cyc_st_6_3_2[0])));
  assign mux_tmp_429 = MUX_s_1_2_2(nor_325_nl, mux_tmp_428, nand_2_nl);
  assign nor_326_nl = ~((rem_12cyc_st_5_3_2[1]) | (~ mux_tmp_429));
  assign nand_3_nl = ~(main_stage_0_6 & asn_itm_5 & (rem_12cyc_st_5_1_0==2'b11) &
      (~ (rem_12cyc_st_5_3_2[0])));
  assign mux_tmp_430 = MUX_s_1_2_2(nor_326_nl, mux_tmp_429, nand_3_nl);
  assign nor_327_nl = ~((rem_12cyc_st_4_3_2[1]) | (~ mux_tmp_430));
  assign nand_4_nl = ~(main_stage_0_5 & asn_itm_4 & (rem_12cyc_st_4_1_0==2'b11) &
      (~ (rem_12cyc_st_4_3_2[0])));
  assign mux_tmp_431 = MUX_s_1_2_2(nor_327_nl, mux_tmp_430, nand_4_nl);
  assign nor_328_nl = ~((rem_12cyc_st_3_3_2[1]) | (~ mux_tmp_431));
  assign nand_5_nl = ~(main_stage_0_4 & asn_itm_3 & (rem_12cyc_st_3_1_0==2'b11) &
      (~ (rem_12cyc_st_3_3_2[0])));
  assign mux_tmp_432 = MUX_s_1_2_2(nor_328_nl, mux_tmp_431, nand_5_nl);
  assign nor_329_nl = ~((rem_12cyc_st_2_3_2[1]) | (~ mux_tmp_432));
  assign nand_6_nl = ~(main_stage_0_3 & asn_itm_2 & (rem_12cyc_st_2_1_0==2'b11) &
      (~ (rem_12cyc_st_2_3_2[0])));
  assign mux_tmp_433 = MUX_s_1_2_2(nor_329_nl, mux_tmp_432, nand_6_nl);
  assign nor_330_nl = ~((rem_12cyc_st_9_3_2[1]) | (~ mux_tmp_433));
  assign nand_7_nl = ~(main_stage_0_10 & asn_itm_9 & (rem_12cyc_st_9_1_0==2'b11)
      & (~ (rem_12cyc_st_9_3_2[0])));
  assign mux_tmp_434 = MUX_s_1_2_2(nor_330_nl, mux_tmp_433, nand_7_nl);
  assign nor_331_nl = ~((rem_12cyc_st_8_3_2[1]) | (~ mux_tmp_434));
  assign nand_8_nl = ~(main_stage_0_9 & asn_itm_8 & (rem_12cyc_st_8_1_0==2'b11) &
      (~ (rem_12cyc_st_8_3_2[0])));
  assign mux_tmp_435 = MUX_s_1_2_2(nor_331_nl, mux_tmp_434, nand_8_nl);
  assign nor_332_nl = ~((rem_12cyc_st_7_3_2[1]) | (~ mux_tmp_435));
  assign nand_9_nl = ~(main_stage_0_8 & asn_itm_7 & (rem_12cyc_st_7_1_0==2'b11) &
      (~ (rem_12cyc_st_7_3_2[0])));
  assign mux_tmp_436 = MUX_s_1_2_2(nor_332_nl, mux_tmp_435, nand_9_nl);
  assign and_934_nl = nand_223_cse & mux_tmp_436;
  assign nand_11_nl = ~(main_stage_0_2 & asn_itm_1 & (rem_12cyc_3_2==2'b10));
  assign mux_tmp_437 = MUX_s_1_2_2(and_934_nl, mux_tmp_436, nand_11_nl);
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_en ) begin
      return_rsci_d <= MUX_v_64_2_2(result_sva_duc_mx0, qelse_acc_nl, mux_13_nl);
      m_buf_sva_12 <= m_buf_sva_11;
      m_buf_sva_11 <= m_buf_sva_10;
      m_buf_sva_10 <= m_buf_sva_9;
      m_buf_sva_9 <= m_buf_sva_8;
      m_buf_sva_8 <= m_buf_sva_7;
      m_buf_sva_7 <= m_buf_sva_6;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      asn_itm_12 <= 1'b0;
      asn_itm_11 <= 1'b0;
      asn_itm_10 <= 1'b0;
      asn_itm_9 <= 1'b0;
      asn_itm_8 <= 1'b0;
      asn_itm_7 <= 1'b0;
      asn_itm_6 <= 1'b0;
      asn_itm_5 <= 1'b0;
      asn_itm_4 <= 1'b0;
      asn_itm_3 <= 1'b0;
      asn_itm_2 <= 1'b0;
      asn_itm_1 <= 1'b0;
      main_stage_0_2 <= 1'b0;
      main_stage_0_3 <= 1'b0;
      main_stage_0_4 <= 1'b0;
      main_stage_0_5 <= 1'b0;
      main_stage_0_6 <= 1'b0;
      main_stage_0_7 <= 1'b0;
      main_stage_0_8 <= 1'b0;
      main_stage_0_9 <= 1'b0;
      main_stage_0_10 <= 1'b0;
      main_stage_0_11 <= 1'b0;
      main_stage_0_12 <= 1'b0;
      main_stage_0_13 <= 1'b0;
    end
    else if ( ccs_ccore_en ) begin
      asn_itm_12 <= asn_itm_11;
      asn_itm_11 <= asn_itm_10;
      asn_itm_10 <= asn_itm_9;
      asn_itm_9 <= asn_itm_8;
      asn_itm_8 <= asn_itm_7;
      asn_itm_7 <= asn_itm_6;
      asn_itm_6 <= asn_itm_5;
      asn_itm_5 <= asn_itm_4;
      asn_itm_4 <= asn_itm_3;
      asn_itm_3 <= asn_itm_2;
      asn_itm_2 <= asn_itm_1;
      asn_itm_1 <= ccs_ccore_start_rsci_idat;
      main_stage_0_2 <= 1'b1;
      main_stage_0_3 <= main_stage_0_2;
      main_stage_0_4 <= main_stage_0_3;
      main_stage_0_5 <= main_stage_0_4;
      main_stage_0_6 <= main_stage_0_5;
      main_stage_0_7 <= main_stage_0_6;
      main_stage_0_8 <= main_stage_0_7;
      main_stage_0_9 <= main_stage_0_8;
      main_stage_0_10 <= main_stage_0_9;
      main_stage_0_11 <= main_stage_0_10;
      main_stage_0_12 <= main_stage_0_11;
      main_stage_0_13 <= main_stage_0_12;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      result_sva_duc <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( asn_itm_12 & main_stage_0_13 & ccs_ccore_en & (~((rem_12cyc_st_12_3_2==2'b11)))
        ) begin
      result_sva_duc <= result_sva_duc_mx0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      rem_12cyc_st_12_3_2 <= 2'b00;
      rem_12cyc_st_12_1_0 <= 2'b00;
    end
    else if ( and_1203_cse ) begin
      rem_12cyc_st_12_3_2 <= rem_12cyc_st_11_3_2;
      rem_12cyc_st_12_1_0 <= rem_12cyc_st_11_1_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1173_cse ) begin
      rem_13_cmp_1_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_3_2_63_0, mut_3_3_63_0,
          mut_3_4_63_0, mut_3_5_63_0, mut_3_6_63_0, mut_3_7_63_0, mut_3_8_63_0, mut_3_9_63_0,
          mut_3_10_63_0, mut_3_11_63_0, {and_dcpl_294 , and_dcpl_300 , and_dcpl_306
          , and_dcpl_312 , and_dcpl_318 , and_dcpl_324 , and_dcpl_330 , and_dcpl_336
          , and_dcpl_342 , and_dcpl_348 , and_tmp_35});
      rem_13_cmp_1_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_2_2_63_0, mut_2_3_63_0,
          mut_2_4_63_0, mut_2_5_63_0, mut_2_6_63_0, mut_2_7_63_0, mut_2_8_63_0, mut_2_9_63_0,
          mut_2_10_63_0, mut_2_11_63_0, {and_dcpl_294 , and_dcpl_300 , and_dcpl_306
          , and_dcpl_312 , and_dcpl_318 , and_dcpl_324 , and_dcpl_330 , and_dcpl_336
          , and_dcpl_342 , and_dcpl_348 , and_tmp_35});
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1175_cse ) begin
      rem_13_cmp_2_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_5_2_63_0, mut_5_3_63_0,
          mut_5_4_63_0, mut_5_5_63_0, mut_5_6_63_0, mut_5_7_63_0, mut_5_8_63_0, mut_5_9_63_0,
          mut_5_10_63_0, mut_5_11_63_0, {and_dcpl_356 , and_dcpl_360 , and_dcpl_364
          , and_dcpl_368 , and_dcpl_372 , and_dcpl_376 , and_dcpl_379 , and_dcpl_382
          , and_dcpl_385 , and_dcpl_388 , mux_tmp_76});
      rem_13_cmp_2_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_4_2_63_0, mut_4_3_63_0,
          mut_4_4_63_0, mut_4_5_63_0, mut_4_6_63_0, mut_4_7_63_0, mut_4_8_63_0, mut_4_9_63_0,
          mut_4_10_63_0, mut_4_11_63_0, {and_dcpl_356 , and_dcpl_360 , and_dcpl_364
          , and_dcpl_368 , and_dcpl_372 , and_dcpl_376 , and_dcpl_379 , and_dcpl_382
          , and_dcpl_385 , and_dcpl_388 , mux_tmp_76});
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1177_cse ) begin
      rem_13_cmp_3_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_7_2_63_0, mut_7_3_63_0,
          mut_7_4_63_0, mut_7_5_63_0, mut_7_6_63_0, mut_7_7_63_0, mut_7_8_63_0, mut_7_9_63_0,
          mut_7_10_63_0, mut_7_11_63_0, {and_dcpl_394 , and_dcpl_397 , and_dcpl_400
          , and_dcpl_403 , and_dcpl_406 , and_dcpl_409 , and_dcpl_413 , and_dcpl_417
          , and_dcpl_421 , and_dcpl_425 , and_tmp_80});
      rem_13_cmp_3_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_6_2_63_0, mut_6_3_63_0,
          mut_6_4_63_0, mut_6_5_63_0, mut_6_6_63_0, mut_6_7_63_0, mut_6_8_63_0, mut_6_9_63_0,
          mut_6_10_63_0, mut_6_11_63_0, {and_dcpl_394 , and_dcpl_397 , and_dcpl_400
          , and_dcpl_403 , and_dcpl_406 , and_dcpl_409 , and_dcpl_413 , and_dcpl_417
          , and_dcpl_421 , and_dcpl_425 , and_tmp_80});
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1179_cse ) begin
      rem_13_cmp_4_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_9_2_63_0, mut_9_3_63_0,
          mut_9_4_63_0, mut_9_5_63_0, mut_9_6_63_0, mut_9_7_63_0, mut_9_8_63_0, mut_9_9_63_0,
          mut_9_10_63_0, mut_9_11_63_0, {and_dcpl_431 , and_dcpl_433 , and_dcpl_435
          , and_dcpl_437 , and_dcpl_439 , and_dcpl_442 , and_dcpl_445 , and_dcpl_448
          , and_dcpl_451 , and_dcpl_454 , mux_tmp_141});
      rem_13_cmp_4_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_8_2_63_0, mut_8_3_63_0,
          mut_8_4_63_0, mut_8_5_63_0, mut_8_6_63_0, mut_8_7_63_0, mut_8_8_63_0, mut_8_9_63_0,
          mut_8_10_63_0, mut_8_11_63_0, {and_dcpl_431 , and_dcpl_433 , and_dcpl_435
          , and_dcpl_437 , and_dcpl_439 , and_dcpl_442 , and_dcpl_445 , and_dcpl_448
          , and_dcpl_451 , and_dcpl_454 , mux_tmp_141});
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1181_cse ) begin
      rem_13_cmp_5_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_11_2_63_0, mut_11_3_63_0,
          mut_11_4_63_0, mut_11_5_63_0, mut_11_6_63_0, mut_11_7_63_0, mut_11_8_63_0,
          mut_11_9_63_0, mut_11_10_63_0, mut_11_11_63_0, {and_dcpl_461 , and_dcpl_465
          , and_dcpl_469 , and_dcpl_473 , and_dcpl_477 , and_dcpl_480 , and_dcpl_483
          , and_dcpl_486 , and_dcpl_489 , and_dcpl_492 , and_tmp_125});
      rem_13_cmp_5_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_10_2_63_0, mut_10_3_63_0,
          mut_10_4_63_0, mut_10_5_63_0, mut_10_6_63_0, mut_10_7_63_0, mut_10_8_63_0,
          mut_10_9_63_0, mut_10_10_63_0, mut_10_11_63_0, {and_dcpl_461 , and_dcpl_465
          , and_dcpl_469 , and_dcpl_473 , and_dcpl_477 , and_dcpl_480 , and_dcpl_483
          , and_dcpl_486 , and_dcpl_489 , and_dcpl_492 , and_tmp_125});
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1183_cse ) begin
      rem_13_cmp_6_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_13_2_63_0, mut_13_3_63_0,
          mut_13_4_63_0, mut_13_5_63_0, mut_13_6_63_0, mut_13_7_63_0, mut_13_8_63_0,
          mut_13_9_63_0, mut_13_10_63_0, mut_13_11_63_0, {and_dcpl_498 , and_dcpl_500
          , and_dcpl_502 , and_dcpl_504 , and_dcpl_506 , and_dcpl_508 , and_dcpl_510
          , and_dcpl_512 , and_dcpl_514 , and_dcpl_516 , mux_tmp_206});
      rem_13_cmp_6_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_12_2_63_0, mut_12_3_63_0,
          mut_12_4_63_0, mut_12_5_63_0, mut_12_6_63_0, mut_12_7_63_0, mut_12_8_63_0,
          mut_12_9_63_0, mut_12_10_63_0, mut_12_11_63_0, {and_dcpl_498 , and_dcpl_500
          , and_dcpl_502 , and_dcpl_504 , and_dcpl_506 , and_dcpl_508 , and_dcpl_510
          , and_dcpl_512 , and_dcpl_514 , and_dcpl_516 , mux_tmp_206});
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1185_cse ) begin
      rem_13_cmp_7_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_15_2_63_0, mut_15_3_63_0,
          mut_15_4_63_0, mut_15_5_63_0, mut_15_6_63_0, mut_15_7_63_0, mut_15_8_63_0,
          mut_15_9_63_0, mut_15_10_63_0, mut_15_11_63_0, {and_dcpl_520 , and_dcpl_523
          , and_dcpl_526 , and_dcpl_529 , and_dcpl_532 , and_dcpl_534 , and_dcpl_536
          , and_dcpl_538 , and_dcpl_540 , and_dcpl_542 , and_tmp_170});
      rem_13_cmp_7_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_14_2_63_0, mut_14_3_63_0,
          mut_14_4_63_0, mut_14_5_63_0, mut_14_6_63_0, mut_14_7_63_0, mut_14_8_63_0,
          mut_14_9_63_0, mut_14_10_63_0, mut_14_11_63_0, {and_dcpl_520 , and_dcpl_523
          , and_dcpl_526 , and_dcpl_529 , and_dcpl_532 , and_dcpl_534 , and_dcpl_536
          , and_dcpl_538 , and_dcpl_540 , and_dcpl_542 , and_tmp_170});
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1187_cse ) begin
      rem_13_cmp_8_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_17_2_63_0, mut_17_3_63_0,
          mut_17_4_63_0, mut_17_5_63_0, mut_17_6_63_0, mut_17_7_63_0, mut_17_8_63_0,
          mut_17_9_63_0, mut_17_10_63_0, mut_17_11_63_0, {and_dcpl_546 , and_dcpl_548
          , and_dcpl_550 , and_dcpl_552 , and_dcpl_554 , and_dcpl_556 , and_dcpl_558
          , and_dcpl_560 , and_dcpl_562 , and_dcpl_564 , mux_tmp_271});
      rem_13_cmp_8_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_16_2_63_0, mut_16_3_63_0,
          mut_16_4_63_0, mut_16_5_63_0, mut_16_6_63_0, mut_16_7_63_0, mut_16_8_63_0,
          mut_16_9_63_0, mut_16_10_63_0, mut_16_11_63_0, {and_dcpl_546 , and_dcpl_548
          , and_dcpl_550 , and_dcpl_552 , and_dcpl_554 , and_dcpl_556 , and_dcpl_558
          , and_dcpl_560 , and_dcpl_562 , and_dcpl_564 , mux_tmp_271});
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1189_cse ) begin
      rem_13_cmp_9_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_19_2_63_0, mut_19_3_63_0,
          mut_19_4_63_0, mut_19_5_63_0, mut_19_6_63_0, mut_19_7_63_0, mut_19_8_63_0,
          mut_19_9_63_0, mut_19_10_63_0, mut_19_11_63_0, {and_dcpl_569 , and_dcpl_573
          , and_dcpl_577 , and_dcpl_581 , and_dcpl_585 , and_dcpl_589 , and_dcpl_593
          , and_dcpl_597 , and_dcpl_601 , and_dcpl_605 , and_tmp_206});
      rem_13_cmp_9_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_18_2_63_0, mut_18_3_63_0,
          mut_18_4_63_0, mut_18_5_63_0, mut_18_6_63_0, mut_18_7_63_0, mut_18_8_63_0,
          mut_18_9_63_0, mut_18_10_63_0, mut_18_11_63_0, {and_dcpl_569 , and_dcpl_573
          , and_dcpl_577 , and_dcpl_581 , and_dcpl_585 , and_dcpl_589 , and_dcpl_593
          , and_dcpl_597 , and_dcpl_601 , and_dcpl_605 , and_tmp_206});
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1191_cse ) begin
      rem_13_cmp_10_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_21_2_63_0, mut_21_3_63_0,
          mut_21_4_63_0, mut_21_5_63_0, mut_21_6_63_0, mut_21_7_63_0, mut_21_8_63_0,
          mut_21_9_63_0, mut_21_10_63_0, mut_21_11_63_0, {and_dcpl_610 , and_dcpl_612
          , and_dcpl_614 , and_dcpl_616 , and_dcpl_618 , and_dcpl_622 , and_dcpl_625
          , and_dcpl_628 , and_dcpl_631 , and_dcpl_634 , mux_tmp_354});
      rem_13_cmp_10_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_20_2_63_0, mut_20_3_63_0,
          mut_20_4_63_0, mut_20_5_63_0, mut_20_6_63_0, mut_20_7_63_0, mut_20_8_63_0,
          mut_20_9_63_0, mut_20_10_63_0, mut_20_11_63_0, {and_dcpl_610 , and_dcpl_612
          , and_dcpl_614 , and_dcpl_616 , and_dcpl_618 , and_dcpl_622 , and_dcpl_625
          , and_dcpl_628 , and_dcpl_631 , and_dcpl_634 , mux_tmp_354});
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1193_cse ) begin
      rem_13_cmp_11_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_23_2_63_0, mut_23_3_63_0,
          mut_23_4_63_0, mut_23_5_63_0, mut_23_6_63_0, mut_23_7_63_0, mut_23_8_63_0,
          mut_23_9_63_0, mut_23_10_63_0, mut_23_11_63_0, {and_dcpl_638 , and_dcpl_641
          , and_dcpl_644 , and_dcpl_647 , and_dcpl_650 , and_dcpl_653 , and_dcpl_657
          , and_dcpl_661 , and_dcpl_665 , and_dcpl_669 , and_tmp_233});
      rem_13_cmp_11_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_22_2_63_0, mut_22_3_63_0,
          mut_22_4_63_0, mut_22_5_63_0, mut_22_6_63_0, mut_22_7_63_0, mut_22_8_63_0,
          mut_22_9_63_0, mut_22_10_63_0, mut_22_11_63_0, {and_dcpl_638 , and_dcpl_641
          , and_dcpl_644 , and_dcpl_647 , and_dcpl_650 , and_dcpl_653 , and_dcpl_657
          , and_dcpl_661 , and_dcpl_665 , and_dcpl_669 , and_tmp_233});
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1195_cse ) begin
      rem_13_cmp_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_1_2_63_0, mut_1_3_63_0,
          mut_1_4_63_0, mut_1_5_63_0, mut_1_6_63_0, mut_1_7_63_0, mut_1_8_63_0, mut_1_9_63_0,
          mut_1_10_63_0, mut_1_11_63_0, {and_dcpl_673 , and_dcpl_675 , and_dcpl_677
          , and_dcpl_679 , and_dcpl_681 , and_dcpl_684 , and_dcpl_687 , and_dcpl_690
          , and_dcpl_693 , and_dcpl_696 , mux_tmp_437});
      rem_13_cmp_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_2_63_0, mut_3_63_0,
          mut_4_63_0, mut_5_63_0, mut_6_63_0, mut_7_63_0, mut_8_63_0, mut_9_63_0,
          mut_10_63_0, mut_11_63_0, {and_dcpl_673 , and_dcpl_675 , and_dcpl_677 ,
          and_dcpl_679 , and_dcpl_681 , and_dcpl_684 , and_dcpl_687 , and_dcpl_690
          , and_dcpl_693 , and_dcpl_696 , mux_tmp_437});
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1205_cse ) begin
      mut_3_11_63_0 <= mut_3_10_63_0;
      mut_2_11_63_0 <= mut_2_10_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1207_cse ) begin
      mut_5_11_63_0 <= mut_5_10_63_0;
      mut_4_11_63_0 <= mut_4_10_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1209_cse ) begin
      mut_7_11_63_0 <= mut_7_10_63_0;
      mut_6_11_63_0 <= mut_6_10_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1211_cse ) begin
      mut_9_11_63_0 <= mut_9_10_63_0;
      mut_8_11_63_0 <= mut_8_10_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1213_cse ) begin
      mut_11_11_63_0 <= mut_11_10_63_0;
      mut_10_11_63_0 <= mut_10_10_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1215_cse ) begin
      mut_13_11_63_0 <= mut_13_10_63_0;
      mut_12_11_63_0 <= mut_12_10_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1217_cse ) begin
      mut_15_11_63_0 <= mut_15_10_63_0;
      mut_14_11_63_0 <= mut_14_10_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1219_cse ) begin
      mut_17_11_63_0 <= mut_17_10_63_0;
      mut_16_11_63_0 <= mut_16_10_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1221_cse ) begin
      mut_19_11_63_0 <= mut_19_10_63_0;
      mut_18_11_63_0 <= mut_18_10_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1223_cse ) begin
      mut_21_11_63_0 <= mut_21_10_63_0;
      mut_20_11_63_0 <= mut_20_10_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1225_cse ) begin
      mut_23_11_63_0 <= mut_23_10_63_0;
      mut_22_11_63_0 <= mut_22_10_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1227_cse ) begin
      mut_1_11_63_0 <= mut_1_10_63_0;
      mut_11_63_0 <= mut_10_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      rem_12cyc_st_11_3_2 <= 2'b00;
      rem_12cyc_st_11_1_0 <= 2'b00;
    end
    else if ( and_1229_cse ) begin
      rem_12cyc_st_11_3_2 <= rem_12cyc_st_10_3_2;
      rem_12cyc_st_11_1_0 <= rem_12cyc_st_10_1_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1231_cse ) begin
      mut_3_10_63_0 <= mut_3_9_63_0;
      mut_2_10_63_0 <= mut_2_9_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1233_cse ) begin
      mut_5_10_63_0 <= mut_5_9_63_0;
      mut_4_10_63_0 <= mut_4_9_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1235_cse ) begin
      mut_7_10_63_0 <= mut_7_9_63_0;
      mut_6_10_63_0 <= mut_6_9_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1237_cse ) begin
      mut_9_10_63_0 <= mut_9_9_63_0;
      mut_8_10_63_0 <= mut_8_9_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1239_cse ) begin
      mut_11_10_63_0 <= mut_11_9_63_0;
      mut_10_10_63_0 <= mut_10_9_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1241_cse ) begin
      mut_13_10_63_0 <= mut_13_9_63_0;
      mut_12_10_63_0 <= mut_12_9_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1243_cse ) begin
      mut_15_10_63_0 <= mut_15_9_63_0;
      mut_14_10_63_0 <= mut_14_9_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1245_cse ) begin
      mut_17_10_63_0 <= mut_17_9_63_0;
      mut_16_10_63_0 <= mut_16_9_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1247_cse ) begin
      mut_19_10_63_0 <= mut_19_9_63_0;
      mut_18_10_63_0 <= mut_18_9_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1249_cse ) begin
      mut_21_10_63_0 <= mut_21_9_63_0;
      mut_20_10_63_0 <= mut_20_9_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1251_cse ) begin
      mut_23_10_63_0 <= mut_23_9_63_0;
      mut_22_10_63_0 <= mut_22_9_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1253_cse ) begin
      mut_1_10_63_0 <= mut_1_9_63_0;
      mut_10_63_0 <= mut_9_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      rem_12cyc_st_10_3_2 <= 2'b00;
      rem_12cyc_st_10_1_0 <= 2'b00;
    end
    else if ( and_1255_cse ) begin
      rem_12cyc_st_10_3_2 <= rem_12cyc_st_9_3_2;
      rem_12cyc_st_10_1_0 <= rem_12cyc_st_9_1_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1257_cse ) begin
      mut_3_9_63_0 <= mut_3_8_63_0;
      mut_2_9_63_0 <= mut_2_8_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1259_cse ) begin
      mut_5_9_63_0 <= mut_5_8_63_0;
      mut_4_9_63_0 <= mut_4_8_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1261_cse ) begin
      mut_7_9_63_0 <= mut_7_8_63_0;
      mut_6_9_63_0 <= mut_6_8_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1263_cse ) begin
      mut_9_9_63_0 <= mut_9_8_63_0;
      mut_8_9_63_0 <= mut_8_8_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1265_cse ) begin
      mut_11_9_63_0 <= mut_11_8_63_0;
      mut_10_9_63_0 <= mut_10_8_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1267_cse ) begin
      mut_13_9_63_0 <= mut_13_8_63_0;
      mut_12_9_63_0 <= mut_12_8_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1269_cse ) begin
      mut_15_9_63_0 <= mut_15_8_63_0;
      mut_14_9_63_0 <= mut_14_8_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1271_cse ) begin
      mut_17_9_63_0 <= mut_17_8_63_0;
      mut_16_9_63_0 <= mut_16_8_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1273_cse ) begin
      mut_19_9_63_0 <= mut_19_8_63_0;
      mut_18_9_63_0 <= mut_18_8_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1275_cse ) begin
      mut_21_9_63_0 <= mut_21_8_63_0;
      mut_20_9_63_0 <= mut_20_8_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1277_cse ) begin
      mut_23_9_63_0 <= mut_23_8_63_0;
      mut_22_9_63_0 <= mut_22_8_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1279_cse ) begin
      mut_1_9_63_0 <= mut_1_8_63_0;
      mut_9_63_0 <= mut_8_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      rem_12cyc_st_9_3_2 <= 2'b00;
      rem_12cyc_st_9_1_0 <= 2'b00;
    end
    else if ( and_1281_cse ) begin
      rem_12cyc_st_9_3_2 <= rem_12cyc_st_8_3_2;
      rem_12cyc_st_9_1_0 <= rem_12cyc_st_8_1_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1283_cse ) begin
      mut_3_8_63_0 <= mut_3_7_63_0;
      mut_2_8_63_0 <= mut_2_7_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1285_cse ) begin
      mut_5_8_63_0 <= mut_5_7_63_0;
      mut_4_8_63_0 <= mut_4_7_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1287_cse ) begin
      mut_7_8_63_0 <= mut_7_7_63_0;
      mut_6_8_63_0 <= mut_6_7_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1289_cse ) begin
      mut_9_8_63_0 <= mut_9_7_63_0;
      mut_8_8_63_0 <= mut_8_7_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1291_cse ) begin
      mut_11_8_63_0 <= mut_11_7_63_0;
      mut_10_8_63_0 <= mut_10_7_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1293_cse ) begin
      mut_13_8_63_0 <= mut_13_7_63_0;
      mut_12_8_63_0 <= mut_12_7_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1295_cse ) begin
      mut_15_8_63_0 <= mut_15_7_63_0;
      mut_14_8_63_0 <= mut_14_7_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1297_cse ) begin
      mut_17_8_63_0 <= mut_17_7_63_0;
      mut_16_8_63_0 <= mut_16_7_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1299_cse ) begin
      mut_19_8_63_0 <= mut_19_7_63_0;
      mut_18_8_63_0 <= mut_18_7_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1301_cse ) begin
      mut_21_8_63_0 <= mut_21_7_63_0;
      mut_20_8_63_0 <= mut_20_7_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1303_cse ) begin
      mut_23_8_63_0 <= mut_23_7_63_0;
      mut_22_8_63_0 <= mut_22_7_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1305_cse ) begin
      mut_1_8_63_0 <= mut_1_7_63_0;
      mut_8_63_0 <= mut_7_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      rem_12cyc_st_8_3_2 <= 2'b00;
      rem_12cyc_st_8_1_0 <= 2'b00;
    end
    else if ( and_1307_cse ) begin
      rem_12cyc_st_8_3_2 <= rem_12cyc_st_7_3_2;
      rem_12cyc_st_8_1_0 <= rem_12cyc_st_7_1_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1309_cse ) begin
      mut_3_7_63_0 <= mut_3_6_63_0;
      mut_2_7_63_0 <= mut_2_6_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1311_cse ) begin
      mut_5_7_63_0 <= mut_5_6_63_0;
      mut_4_7_63_0 <= mut_4_6_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1313_cse ) begin
      mut_7_7_63_0 <= mut_7_6_63_0;
      mut_6_7_63_0 <= mut_6_6_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1315_cse ) begin
      mut_9_7_63_0 <= mut_9_6_63_0;
      mut_8_7_63_0 <= mut_8_6_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1317_cse ) begin
      mut_11_7_63_0 <= mut_11_6_63_0;
      mut_10_7_63_0 <= mut_10_6_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1319_cse ) begin
      mut_13_7_63_0 <= mut_13_6_63_0;
      mut_12_7_63_0 <= mut_12_6_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1321_cse ) begin
      mut_15_7_63_0 <= mut_15_6_63_0;
      mut_14_7_63_0 <= mut_14_6_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1323_cse ) begin
      mut_17_7_63_0 <= mut_17_6_63_0;
      mut_16_7_63_0 <= mut_16_6_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1325_cse ) begin
      mut_19_7_63_0 <= mut_19_6_63_0;
      mut_18_7_63_0 <= mut_18_6_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1327_cse ) begin
      mut_21_7_63_0 <= mut_21_6_63_0;
      mut_20_7_63_0 <= mut_20_6_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1329_cse ) begin
      mut_23_7_63_0 <= mut_23_6_63_0;
      mut_22_7_63_0 <= mut_22_6_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1331_cse ) begin
      mut_1_7_63_0 <= mut_1_6_63_0;
      mut_7_63_0 <= mut_6_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      rem_12cyc_st_7_3_2 <= 2'b00;
      rem_12cyc_st_7_1_0 <= 2'b00;
    end
    else if ( and_1333_cse ) begin
      rem_12cyc_st_7_3_2 <= rem_12cyc_st_6_3_2;
      rem_12cyc_st_7_1_0 <= rem_12cyc_st_6_1_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1335_cse ) begin
      mut_3_6_63_0 <= mut_3_5_63_0;
      mut_2_6_63_0 <= mut_2_5_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1337_cse ) begin
      mut_5_6_63_0 <= mut_5_5_63_0;
      mut_4_6_63_0 <= mut_4_5_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1339_cse ) begin
      mut_7_6_63_0 <= mut_7_5_63_0;
      mut_6_6_63_0 <= mut_6_5_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1341_cse ) begin
      mut_9_6_63_0 <= mut_9_5_63_0;
      mut_8_6_63_0 <= mut_8_5_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1343_cse ) begin
      mut_11_6_63_0 <= mut_11_5_63_0;
      mut_10_6_63_0 <= mut_10_5_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1345_cse ) begin
      mut_13_6_63_0 <= mut_13_5_63_0;
      mut_12_6_63_0 <= mut_12_5_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1347_cse ) begin
      mut_15_6_63_0 <= mut_15_5_63_0;
      mut_14_6_63_0 <= mut_14_5_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1349_cse ) begin
      mut_17_6_63_0 <= mut_17_5_63_0;
      mut_16_6_63_0 <= mut_16_5_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1351_cse ) begin
      mut_19_6_63_0 <= mut_19_5_63_0;
      mut_18_6_63_0 <= mut_18_5_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1353_cse ) begin
      mut_21_6_63_0 <= mut_21_5_63_0;
      mut_20_6_63_0 <= mut_20_5_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1355_cse ) begin
      mut_23_6_63_0 <= mut_23_5_63_0;
      mut_22_6_63_0 <= mut_22_5_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1357_cse ) begin
      mut_1_6_63_0 <= mut_1_5_63_0;
      mut_6_63_0 <= mut_5_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1359_cse ) begin
      m_buf_sva_6 <= m_buf_sva_5;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      rem_12cyc_st_6_3_2 <= 2'b00;
      rem_12cyc_st_6_1_0 <= 2'b00;
    end
    else if ( and_1359_cse ) begin
      rem_12cyc_st_6_3_2 <= rem_12cyc_st_5_3_2;
      rem_12cyc_st_6_1_0 <= rem_12cyc_st_5_1_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1361_cse ) begin
      mut_3_5_63_0 <= mut_3_4_63_0;
      mut_2_5_63_0 <= mut_2_4_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1363_cse ) begin
      mut_5_5_63_0 <= mut_5_4_63_0;
      mut_4_5_63_0 <= mut_4_4_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1365_cse ) begin
      mut_7_5_63_0 <= mut_7_4_63_0;
      mut_6_5_63_0 <= mut_6_4_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1367_cse ) begin
      mut_9_5_63_0 <= mut_9_4_63_0;
      mut_8_5_63_0 <= mut_8_4_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1369_cse ) begin
      mut_11_5_63_0 <= mut_11_4_63_0;
      mut_10_5_63_0 <= mut_10_4_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1371_cse ) begin
      mut_13_5_63_0 <= mut_13_4_63_0;
      mut_12_5_63_0 <= mut_12_4_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1373_cse ) begin
      mut_15_5_63_0 <= mut_15_4_63_0;
      mut_14_5_63_0 <= mut_14_4_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1375_cse ) begin
      mut_17_5_63_0 <= mut_17_4_63_0;
      mut_16_5_63_0 <= mut_16_4_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1377_cse ) begin
      mut_19_5_63_0 <= mut_19_4_63_0;
      mut_18_5_63_0 <= mut_18_4_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1379_cse ) begin
      mut_21_5_63_0 <= mut_21_4_63_0;
      mut_20_5_63_0 <= mut_20_4_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1381_cse ) begin
      mut_23_5_63_0 <= mut_23_4_63_0;
      mut_22_5_63_0 <= mut_22_4_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1383_cse ) begin
      mut_1_5_63_0 <= mut_1_4_63_0;
      mut_5_63_0 <= mut_4_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1385_cse ) begin
      m_buf_sva_5 <= m_buf_sva_4;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      rem_12cyc_st_5_3_2 <= 2'b00;
      rem_12cyc_st_5_1_0 <= 2'b00;
    end
    else if ( and_1385_cse ) begin
      rem_12cyc_st_5_3_2 <= rem_12cyc_st_4_3_2;
      rem_12cyc_st_5_1_0 <= rem_12cyc_st_4_1_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1387_cse ) begin
      mut_3_4_63_0 <= mut_3_3_63_0;
      mut_2_4_63_0 <= mut_2_3_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1389_cse ) begin
      mut_5_4_63_0 <= mut_5_3_63_0;
      mut_4_4_63_0 <= mut_4_3_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1391_cse ) begin
      mut_7_4_63_0 <= mut_7_3_63_0;
      mut_6_4_63_0 <= mut_6_3_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1393_cse ) begin
      mut_9_4_63_0 <= mut_9_3_63_0;
      mut_8_4_63_0 <= mut_8_3_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1395_cse ) begin
      mut_11_4_63_0 <= mut_11_3_63_0;
      mut_10_4_63_0 <= mut_10_3_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1397_cse ) begin
      mut_13_4_63_0 <= mut_13_3_63_0;
      mut_12_4_63_0 <= mut_12_3_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1399_cse ) begin
      mut_15_4_63_0 <= mut_15_3_63_0;
      mut_14_4_63_0 <= mut_14_3_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1401_cse ) begin
      mut_17_4_63_0 <= mut_17_3_63_0;
      mut_16_4_63_0 <= mut_16_3_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1403_cse ) begin
      mut_19_4_63_0 <= mut_19_3_63_0;
      mut_18_4_63_0 <= mut_18_3_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1405_cse ) begin
      mut_21_4_63_0 <= mut_21_3_63_0;
      mut_20_4_63_0 <= mut_20_3_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1407_cse ) begin
      mut_23_4_63_0 <= mut_23_3_63_0;
      mut_22_4_63_0 <= mut_22_3_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1409_cse ) begin
      mut_1_4_63_0 <= mut_1_3_63_0;
      mut_4_63_0 <= mut_3_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1411_cse ) begin
      m_buf_sva_4 <= m_buf_sva_3;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      rem_12cyc_st_4_3_2 <= 2'b00;
      rem_12cyc_st_4_1_0 <= 2'b00;
    end
    else if ( and_1411_cse ) begin
      rem_12cyc_st_4_3_2 <= rem_12cyc_st_3_3_2;
      rem_12cyc_st_4_1_0 <= rem_12cyc_st_3_1_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1413_cse ) begin
      mut_3_3_63_0 <= mut_3_2_63_0;
      mut_2_3_63_0 <= mut_2_2_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1415_cse ) begin
      mut_5_3_63_0 <= mut_5_2_63_0;
      mut_4_3_63_0 <= mut_4_2_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1417_cse ) begin
      mut_7_3_63_0 <= mut_7_2_63_0;
      mut_6_3_63_0 <= mut_6_2_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1419_cse ) begin
      mut_9_3_63_0 <= mut_9_2_63_0;
      mut_8_3_63_0 <= mut_8_2_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1421_cse ) begin
      mut_11_3_63_0 <= mut_11_2_63_0;
      mut_10_3_63_0 <= mut_10_2_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1423_cse ) begin
      mut_13_3_63_0 <= mut_13_2_63_0;
      mut_12_3_63_0 <= mut_12_2_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1425_cse ) begin
      mut_15_3_63_0 <= mut_15_2_63_0;
      mut_14_3_63_0 <= mut_14_2_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1427_cse ) begin
      mut_17_3_63_0 <= mut_17_2_63_0;
      mut_16_3_63_0 <= mut_16_2_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1429_cse ) begin
      mut_19_3_63_0 <= mut_19_2_63_0;
      mut_18_3_63_0 <= mut_18_2_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1431_cse ) begin
      mut_21_3_63_0 <= mut_21_2_63_0;
      mut_20_3_63_0 <= mut_20_2_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1433_cse ) begin
      mut_23_3_63_0 <= mut_23_2_63_0;
      mut_22_3_63_0 <= mut_22_2_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1435_cse ) begin
      mut_1_3_63_0 <= mut_1_2_63_0;
      mut_3_63_0 <= mut_2_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1437_cse ) begin
      m_buf_sva_3 <= m_buf_sva_2;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      rem_12cyc_st_3_3_2 <= 2'b00;
      rem_12cyc_st_3_1_0 <= 2'b00;
    end
    else if ( and_1437_cse ) begin
      rem_12cyc_st_3_3_2 <= rem_12cyc_st_2_3_2;
      rem_12cyc_st_3_1_0 <= rem_12cyc_st_2_1_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1439_cse ) begin
      mut_3_2_63_0 <= rem_13_cmp_1_b_63_0;
      mut_2_2_63_0 <= rem_13_cmp_1_a_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1441_cse ) begin
      mut_5_2_63_0 <= rem_13_cmp_2_b_63_0;
      mut_4_2_63_0 <= rem_13_cmp_2_a_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1443_cse ) begin
      mut_7_2_63_0 <= rem_13_cmp_3_b_63_0;
      mut_6_2_63_0 <= rem_13_cmp_3_a_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1445_cse ) begin
      mut_9_2_63_0 <= rem_13_cmp_4_b_63_0;
      mut_8_2_63_0 <= rem_13_cmp_4_a_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1447_cse ) begin
      mut_11_2_63_0 <= rem_13_cmp_5_b_63_0;
      mut_10_2_63_0 <= rem_13_cmp_5_a_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1449_cse ) begin
      mut_13_2_63_0 <= rem_13_cmp_6_b_63_0;
      mut_12_2_63_0 <= rem_13_cmp_6_a_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1451_cse ) begin
      mut_15_2_63_0 <= rem_13_cmp_7_b_63_0;
      mut_14_2_63_0 <= rem_13_cmp_7_a_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1453_cse ) begin
      mut_17_2_63_0 <= rem_13_cmp_8_b_63_0;
      mut_16_2_63_0 <= rem_13_cmp_8_a_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1455_cse ) begin
      mut_19_2_63_0 <= rem_13_cmp_9_b_63_0;
      mut_18_2_63_0 <= rem_13_cmp_9_a_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1457_cse ) begin
      mut_21_2_63_0 <= rem_13_cmp_10_b_63_0;
      mut_20_2_63_0 <= rem_13_cmp_10_a_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1459_cse ) begin
      mut_23_2_63_0 <= rem_13_cmp_11_b_63_0;
      mut_22_2_63_0 <= rem_13_cmp_11_a_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1461_cse ) begin
      mut_1_2_63_0 <= rem_13_cmp_b_63_0;
      mut_2_63_0 <= rem_13_cmp_a_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1463_cse ) begin
      m_buf_sva_2 <= m_buf_sva_1;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      rem_12cyc_st_2_3_2 <= 2'b00;
      rem_12cyc_st_2_1_0 <= 2'b00;
    end
    else if ( and_1463_cse ) begin
      rem_12cyc_st_2_3_2 <= rem_12cyc_3_2;
      rem_12cyc_st_2_1_0 <= rem_12cyc_1_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1197_cse ) begin
      m_buf_sva_1 <= m_rsci_idat;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      rem_12cyc_3_2 <= 2'b00;
      rem_12cyc_1_0 <= 2'b00;
    end
    else if ( and_1197_cse ) begin
      rem_12cyc_3_2 <= acc_tmp;
      rem_12cyc_1_0 <= acc_1_tmp[1:0];
    end
  end
  assign nl_qelse_acc_nl = result_sva_duc_mx0 + m_buf_sva_12;
  assign qelse_acc_nl = nl_qelse_acc_nl[63:0];
  assign mux_10_nl = MUX_s_1_2_2((rem_13_cmp_1_z[63]), (rem_13_cmp_3_z[63]), rem_12cyc_st_12_1_0[1]);
  assign mux_9_nl = MUX_s_1_2_2((rem_13_cmp_2_z[63]), (rem_13_cmp_4_z[63]), rem_12cyc_st_12_1_0[1]);
  assign mux_11_nl = MUX_s_1_2_2(mux_10_nl, mux_9_nl, rem_12cyc_st_12_1_0[0]);
  assign mux_7_nl = MUX_s_1_2_2((rem_13_cmp_9_z[63]), (rem_13_cmp_11_z[63]), rem_12cyc_st_12_1_0[1]);
  assign mux_6_nl = MUX_s_1_2_2((rem_13_cmp_10_z[63]), (rem_13_cmp_z[63]), rem_12cyc_st_12_1_0[1]);
  assign mux_8_nl = MUX_s_1_2_2(mux_7_nl, mux_6_nl, rem_12cyc_st_12_1_0[0]);
  assign mux_12_nl = MUX_s_1_2_2(mux_11_nl, mux_8_nl, rem_12cyc_st_12_3_2[1]);
  assign mux_3_nl = MUX_s_1_2_2((rem_13_cmp_5_z[63]), (rem_13_cmp_7_z[63]), rem_12cyc_st_12_1_0[1]);
  assign mux_2_nl = MUX_s_1_2_2((rem_13_cmp_6_z[63]), (rem_13_cmp_8_z[63]), rem_12cyc_st_12_1_0[1]);
  assign mux_4_nl = MUX_s_1_2_2(mux_3_nl, mux_2_nl, rem_12cyc_st_12_1_0[0]);
  assign mux_5_nl = MUX_s_1_2_2(mux_4_nl, (result_sva_duc[63]), rem_12cyc_st_12_3_2[1]);
  assign mux_13_nl = MUX_s_1_2_2(mux_12_nl, mux_5_nl, rem_12cyc_st_12_3_2[0]);

  function automatic [63:0] MUX1HOT_v_64_11_2;
    input [63:0] input_10;
    input [63:0] input_9;
    input [63:0] input_8;
    input [63:0] input_7;
    input [63:0] input_6;
    input [63:0] input_5;
    input [63:0] input_4;
    input [63:0] input_3;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [10:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    result = result | ( input_3 & {64{sel[3]}});
    result = result | ( input_4 & {64{sel[4]}});
    result = result | ( input_5 & {64{sel[5]}});
    result = result | ( input_6 & {64{sel[6]}});
    result = result | ( input_7 & {64{sel[7]}});
    result = result | ( input_8 & {64{sel[8]}});
    result = result | ( input_9 & {64{sel[9]}});
    result = result | ( input_10 & {64{sel[10]}});
    MUX1HOT_v_64_11_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_13_2;
    input [63:0] input_12;
    input [63:0] input_11;
    input [63:0] input_10;
    input [63:0] input_9;
    input [63:0] input_8;
    input [63:0] input_7;
    input [63:0] input_6;
    input [63:0] input_5;
    input [63:0] input_4;
    input [63:0] input_3;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [12:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    result = result | ( input_3 & {64{sel[3]}});
    result = result | ( input_4 & {64{sel[4]}});
    result = result | ( input_5 & {64{sel[5]}});
    result = result | ( input_6 & {64{sel[6]}});
    result = result | ( input_7 & {64{sel[7]}});
    result = result | ( input_8 & {64{sel[8]}});
    result = result | ( input_9 & {64{sel[9]}});
    result = result | ( input_10 & {64{sel[10]}});
    result = result | ( input_11 & {64{sel[11]}});
    result = result | ( input_12 & {64{sel[12]}});
    MUX1HOT_v_64_13_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function automatic [1:0] conv_u2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_2 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    modulo_dev
// ------------------------------------------------------------------


module modulo_dev (
  base_rsc_dat, m_rsc_dat, return_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk,
      ccs_ccore_srst, ccs_ccore_en
);
  input [63:0] base_rsc_dat;
  input [63:0] m_rsc_dat;
  output [63:0] return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_srst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  modulo_dev_core modulo_dev_core_inst (
      .base_rsc_dat(base_rsc_dat),
      .m_rsc_dat(m_rsc_dat),
      .return_rsc_z(return_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_srst(ccs_ccore_srst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_div_beh.v 
module mgc_div(a,b,z);
   parameter width_a = 8;
   parameter width_b = 8;
   parameter signd = 1;
   input [width_a-1:0] a;
   input [width_b-1:0] b; 
   output [width_a-1:0] z;  
   reg  [width_a-1:0] z;

   always@(a or b)
     begin
	if(signd)
	  div_s(a,b,z);
	else
          div_u(a,b,z);
     end


//-----------------------------------------------------------------
//     -- Vectorized Overloaded Arithmetic Operators
//-----------------------------------------------------------------
   
   function [width_a-1:0] fabs_l; 
      input [width_a-1:0] arg1;
      begin
         case(arg1[width_a-1])
            1'b1:
               fabs_l = {(width_a){1'b0}} - arg1;
            default: // was: 1'b0:
               fabs_l = arg1;
         endcase
      end
   endfunction
   
   function [width_b-1:0] fabs_r; 
      input [width_b-1:0] arg1;
      begin
         case (arg1[width_b-1])
            1'b1:
               fabs_r =  {(width_b){1'b0}} - arg1;
            default: // was: 1'b0:
               fabs_r = arg1;
         endcase
      end
   endfunction

   function [width_b:0] minus;
     input [width_b:0] in1;
     input [width_b:0] in2;
     reg [width_b+1:0] tmp;
     begin
       tmp = in1 - in2;
       minus = tmp[width_b:0];
     end
   endfunction

   
   task divmod;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      output [width_b-1:0] rmod;
      
      parameter llen = width_a;
      parameter rlen = width_b;
      reg [(llen+rlen)-1:0] lbuf;
      reg [rlen:0] diff;
	  integer i;
      begin
	 lbuf = {(llen+rlen){1'b0}};
//64'b0;
	 lbuf[llen-1:0] = l;
	 for(i=width_a-1;i>=0;i=i-1)
	   begin
              diff = minus(lbuf[(llen+rlen)-1:llen-1], {1'b0,r});
	      rdiv[i] = ~diff[rlen];
	      if(diff[rlen] == 0)
		lbuf[(llen+rlen)-1:llen-1] = diff;
	      lbuf[(llen+rlen)-1:1] = lbuf[(llen+rlen)-2:0];
	   end
	 rmod = lbuf[(llen+rlen)-1:llen];
      end
   endtask
      

   task div_u;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(l, r, rdiv, rmod);
      end
   endtask
   
   task mod_u;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_b-1:0] rmod;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(l, r, rdiv, rmod);
      end
   endtask

   task rem_u; 
      input [width_a-1:0] l;
      input [width_b-1:0] r;    
      output [width_b-1:0] rmod;
      begin
	 mod_u(l,r,rmod);
      end
   endtask // rem_u

   task div_s;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(fabs_l(l), fabs_r(r),rdiv,rmod);
	 if(l[width_a-1] != r[width_b-1])
	   rdiv = {(width_a){1'b0}} - rdiv;
      end
   endtask

   task mod_s;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_b-1:0] rmod;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      reg [width_b-1:0] rnul;
      reg [width_b:0] rmod_t;
      begin
         rnul = {width_b{1'b0}};
	 divmod(fabs_l(l), fabs_r(r), rdiv, rmod);
         if (l[width_a-1])
	   rmod = {(width_b){1'b0}} - rmod;
	 if((rmod != rnul) && (l[width_a-1] != r[width_b-1]))
            begin
               rmod_t = r + rmod;
               rmod = rmod_t[width_b-1:0];
            end
      end
   endtask // mod_s
   
   task rem_s; 
      input [width_a-1:0] l;
      input [width_b-1:0] r;    
      output [width_b-1:0] rmod;   
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(fabs_l(l),fabs_r(r),rdiv,rmod);
	 if(l[width_a-1])
	   rmod = {(width_b){1'b0}} - rmod;
      end
   endtask

  endmodule

//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_shift_l_beh_v5.v 
module mgc_shift_l_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
   if (signd_a)
   begin: SGNED
      assign z = fshl_u(a,s,a[width_a-1]);
   end
   else
   begin: UNSGNED
      assign z = fshl_u(a,s,1'b0);
   end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u

endmodule

//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5c/896140 Production Release
//  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
// 
//  Generated by:   yl7897@newnano.poly.edu
//  Generated date: Wed Jul 21 01:49:29 2021
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_23_6_64_64_64_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_23_6_64_64_64_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [5:0] adra;
  input [5:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_22_6_64_64_64_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_22_6_64_64_64_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [5:0] adra;
  input [5:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_21_6_64_64_64_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_21_6_64_64_64_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [5:0] adra;
  input [5:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_20_6_64_64_64_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_20_6_64_64_64_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [5:0] adra;
  input [5:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_19_6_64_64_64_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_19_6_64_64_64_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [5:0] adra;
  input [5:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_18_6_64_64_64_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_18_6_64_64_64_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [5:0] adra;
  input [5:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_17_6_64_64_64_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_17_6_64_64_64_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [5:0] adra;
  input [5:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_16_6_64_64_64_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_16_6_64_64_64_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [5:0] adra;
  input [5:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_15_6_64_64_64_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_15_6_64_64_64_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [5:0] adra;
  input [5:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_14_6_64_64_64_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_14_6_64_64_64_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [5:0] adra;
  input [5:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_13_6_64_64_64_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_13_6_64_64_64_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [5:0] adra;
  input [5:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_12_6_64_64_64_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_12_6_64_64_64_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [5:0] adra;
  input [5:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_11_6_64_64_64_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_11_6_64_64_64_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [5:0] adra;
  input [5:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_10_6_64_64_64_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_10_6_64_64_64_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [5:0] adra;
  input [5:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_9_6_64_64_64_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_9_6_64_64_64_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [5:0] adra;
  input [5:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_8_6_64_64_64_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_8_6_64_64_64_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [5:0] adra;
  input [5:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module inPlaceNTT_DIF_core_core_fsm (
  clk, rst, fsm_output, STAGE_MAIN_LOOP_C_3_tr0, modExp_dev_while_C_11_tr0, STAGE_VEC_LOOP_C_0_tr0,
      COMP_LOOP_C_16_tr0, COMP_LOOP_1_modExp_dev_1_while_C_11_tr0, COMP_LOOP_C_45_tr0,
      COMP_LOOP_2_modExp_dev_1_while_C_11_tr0, COMP_LOOP_C_90_tr0, COMP_LOOP_3_modExp_dev_1_while_C_11_tr0,
      COMP_LOOP_C_135_tr0, COMP_LOOP_4_modExp_dev_1_while_C_11_tr0, COMP_LOOP_C_180_tr0,
      COMP_LOOP_5_modExp_dev_1_while_C_11_tr0, COMP_LOOP_C_225_tr0, COMP_LOOP_6_modExp_dev_1_while_C_11_tr0,
      COMP_LOOP_C_270_tr0, COMP_LOOP_7_modExp_dev_1_while_C_11_tr0, COMP_LOOP_C_315_tr0,
      COMP_LOOP_8_modExp_dev_1_while_C_11_tr0, COMP_LOOP_C_360_tr0, COMP_LOOP_9_modExp_dev_1_while_C_11_tr0,
      COMP_LOOP_C_405_tr0, COMP_LOOP_10_modExp_dev_1_while_C_11_tr0, COMP_LOOP_C_450_tr0,
      COMP_LOOP_11_modExp_dev_1_while_C_11_tr0, COMP_LOOP_C_495_tr0, COMP_LOOP_12_modExp_dev_1_while_C_11_tr0,
      COMP_LOOP_C_540_tr0, COMP_LOOP_13_modExp_dev_1_while_C_11_tr0, COMP_LOOP_C_585_tr0,
      COMP_LOOP_14_modExp_dev_1_while_C_11_tr0, COMP_LOOP_C_630_tr0, COMP_LOOP_15_modExp_dev_1_while_C_11_tr0,
      COMP_LOOP_C_675_tr0, COMP_LOOP_16_modExp_dev_1_while_C_11_tr0, COMP_LOOP_C_720_tr0,
      STAGE_VEC_LOOP_C_1_tr0, STAGE_MAIN_LOOP_C_4_tr0
);
  input clk;
  input rst;
  output [9:0] fsm_output;
  reg [9:0] fsm_output;
  input STAGE_MAIN_LOOP_C_3_tr0;
  input modExp_dev_while_C_11_tr0;
  input STAGE_VEC_LOOP_C_0_tr0;
  input COMP_LOOP_C_16_tr0;
  input COMP_LOOP_1_modExp_dev_1_while_C_11_tr0;
  input COMP_LOOP_C_45_tr0;
  input COMP_LOOP_2_modExp_dev_1_while_C_11_tr0;
  input COMP_LOOP_C_90_tr0;
  input COMP_LOOP_3_modExp_dev_1_while_C_11_tr0;
  input COMP_LOOP_C_135_tr0;
  input COMP_LOOP_4_modExp_dev_1_while_C_11_tr0;
  input COMP_LOOP_C_180_tr0;
  input COMP_LOOP_5_modExp_dev_1_while_C_11_tr0;
  input COMP_LOOP_C_225_tr0;
  input COMP_LOOP_6_modExp_dev_1_while_C_11_tr0;
  input COMP_LOOP_C_270_tr0;
  input COMP_LOOP_7_modExp_dev_1_while_C_11_tr0;
  input COMP_LOOP_C_315_tr0;
  input COMP_LOOP_8_modExp_dev_1_while_C_11_tr0;
  input COMP_LOOP_C_360_tr0;
  input COMP_LOOP_9_modExp_dev_1_while_C_11_tr0;
  input COMP_LOOP_C_405_tr0;
  input COMP_LOOP_10_modExp_dev_1_while_C_11_tr0;
  input COMP_LOOP_C_450_tr0;
  input COMP_LOOP_11_modExp_dev_1_while_C_11_tr0;
  input COMP_LOOP_C_495_tr0;
  input COMP_LOOP_12_modExp_dev_1_while_C_11_tr0;
  input COMP_LOOP_C_540_tr0;
  input COMP_LOOP_13_modExp_dev_1_while_C_11_tr0;
  input COMP_LOOP_C_585_tr0;
  input COMP_LOOP_14_modExp_dev_1_while_C_11_tr0;
  input COMP_LOOP_C_630_tr0;
  input COMP_LOOP_15_modExp_dev_1_while_C_11_tr0;
  input COMP_LOOP_C_675_tr0;
  input COMP_LOOP_16_modExp_dev_1_while_C_11_tr0;
  input COMP_LOOP_C_720_tr0;
  input STAGE_VEC_LOOP_C_1_tr0;
  input STAGE_MAIN_LOOP_C_4_tr0;


  // FSM State Type Declaration for inPlaceNTT_DIF_core_core_fsm_1
  parameter
    main_C_0 = 10'd0,
    STAGE_MAIN_LOOP_C_0 = 10'd1,
    STAGE_MAIN_LOOP_C_1 = 10'd2,
    STAGE_MAIN_LOOP_C_2 = 10'd3,
    STAGE_MAIN_LOOP_C_3 = 10'd4,
    modExp_dev_while_C_0 = 10'd5,
    modExp_dev_while_C_1 = 10'd6,
    modExp_dev_while_C_2 = 10'd7,
    modExp_dev_while_C_3 = 10'd8,
    modExp_dev_while_C_4 = 10'd9,
    modExp_dev_while_C_5 = 10'd10,
    modExp_dev_while_C_6 = 10'd11,
    modExp_dev_while_C_7 = 10'd12,
    modExp_dev_while_C_8 = 10'd13,
    modExp_dev_while_C_9 = 10'd14,
    modExp_dev_while_C_10 = 10'd15,
    modExp_dev_while_C_11 = 10'd16,
    STAGE_VEC_LOOP_C_0 = 10'd17,
    COMP_LOOP_C_0 = 10'd18,
    COMP_LOOP_C_1 = 10'd19,
    COMP_LOOP_C_2 = 10'd20,
    COMP_LOOP_C_3 = 10'd21,
    COMP_LOOP_C_4 = 10'd22,
    COMP_LOOP_C_5 = 10'd23,
    COMP_LOOP_C_6 = 10'd24,
    COMP_LOOP_C_7 = 10'd25,
    COMP_LOOP_C_8 = 10'd26,
    COMP_LOOP_C_9 = 10'd27,
    COMP_LOOP_C_10 = 10'd28,
    COMP_LOOP_C_11 = 10'd29,
    COMP_LOOP_C_12 = 10'd30,
    COMP_LOOP_C_13 = 10'd31,
    COMP_LOOP_C_14 = 10'd32,
    COMP_LOOP_C_15 = 10'd33,
    COMP_LOOP_C_16 = 10'd34,
    COMP_LOOP_1_modExp_dev_1_while_C_0 = 10'd35,
    COMP_LOOP_1_modExp_dev_1_while_C_1 = 10'd36,
    COMP_LOOP_1_modExp_dev_1_while_C_2 = 10'd37,
    COMP_LOOP_1_modExp_dev_1_while_C_3 = 10'd38,
    COMP_LOOP_1_modExp_dev_1_while_C_4 = 10'd39,
    COMP_LOOP_1_modExp_dev_1_while_C_5 = 10'd40,
    COMP_LOOP_1_modExp_dev_1_while_C_6 = 10'd41,
    COMP_LOOP_1_modExp_dev_1_while_C_7 = 10'd42,
    COMP_LOOP_1_modExp_dev_1_while_C_8 = 10'd43,
    COMP_LOOP_1_modExp_dev_1_while_C_9 = 10'd44,
    COMP_LOOP_1_modExp_dev_1_while_C_10 = 10'd45,
    COMP_LOOP_1_modExp_dev_1_while_C_11 = 10'd46,
    COMP_LOOP_C_17 = 10'd47,
    COMP_LOOP_C_18 = 10'd48,
    COMP_LOOP_C_19 = 10'd49,
    COMP_LOOP_C_20 = 10'd50,
    COMP_LOOP_C_21 = 10'd51,
    COMP_LOOP_C_22 = 10'd52,
    COMP_LOOP_C_23 = 10'd53,
    COMP_LOOP_C_24 = 10'd54,
    COMP_LOOP_C_25 = 10'd55,
    COMP_LOOP_C_26 = 10'd56,
    COMP_LOOP_C_27 = 10'd57,
    COMP_LOOP_C_28 = 10'd58,
    COMP_LOOP_C_29 = 10'd59,
    COMP_LOOP_C_30 = 10'd60,
    COMP_LOOP_C_31 = 10'd61,
    COMP_LOOP_C_32 = 10'd62,
    COMP_LOOP_C_33 = 10'd63,
    COMP_LOOP_C_34 = 10'd64,
    COMP_LOOP_C_35 = 10'd65,
    COMP_LOOP_C_36 = 10'd66,
    COMP_LOOP_C_37 = 10'd67,
    COMP_LOOP_C_38 = 10'd68,
    COMP_LOOP_C_39 = 10'd69,
    COMP_LOOP_C_40 = 10'd70,
    COMP_LOOP_C_41 = 10'd71,
    COMP_LOOP_C_42 = 10'd72,
    COMP_LOOP_C_43 = 10'd73,
    COMP_LOOP_C_44 = 10'd74,
    COMP_LOOP_C_45 = 10'd75,
    COMP_LOOP_C_46 = 10'd76,
    COMP_LOOP_C_47 = 10'd77,
    COMP_LOOP_C_48 = 10'd78,
    COMP_LOOP_C_49 = 10'd79,
    COMP_LOOP_C_50 = 10'd80,
    COMP_LOOP_C_51 = 10'd81,
    COMP_LOOP_C_52 = 10'd82,
    COMP_LOOP_C_53 = 10'd83,
    COMP_LOOP_C_54 = 10'd84,
    COMP_LOOP_C_55 = 10'd85,
    COMP_LOOP_C_56 = 10'd86,
    COMP_LOOP_C_57 = 10'd87,
    COMP_LOOP_C_58 = 10'd88,
    COMP_LOOP_C_59 = 10'd89,
    COMP_LOOP_C_60 = 10'd90,
    COMP_LOOP_C_61 = 10'd91,
    COMP_LOOP_2_modExp_dev_1_while_C_0 = 10'd92,
    COMP_LOOP_2_modExp_dev_1_while_C_1 = 10'd93,
    COMP_LOOP_2_modExp_dev_1_while_C_2 = 10'd94,
    COMP_LOOP_2_modExp_dev_1_while_C_3 = 10'd95,
    COMP_LOOP_2_modExp_dev_1_while_C_4 = 10'd96,
    COMP_LOOP_2_modExp_dev_1_while_C_5 = 10'd97,
    COMP_LOOP_2_modExp_dev_1_while_C_6 = 10'd98,
    COMP_LOOP_2_modExp_dev_1_while_C_7 = 10'd99,
    COMP_LOOP_2_modExp_dev_1_while_C_8 = 10'd100,
    COMP_LOOP_2_modExp_dev_1_while_C_9 = 10'd101,
    COMP_LOOP_2_modExp_dev_1_while_C_10 = 10'd102,
    COMP_LOOP_2_modExp_dev_1_while_C_11 = 10'd103,
    COMP_LOOP_C_62 = 10'd104,
    COMP_LOOP_C_63 = 10'd105,
    COMP_LOOP_C_64 = 10'd106,
    COMP_LOOP_C_65 = 10'd107,
    COMP_LOOP_C_66 = 10'd108,
    COMP_LOOP_C_67 = 10'd109,
    COMP_LOOP_C_68 = 10'd110,
    COMP_LOOP_C_69 = 10'd111,
    COMP_LOOP_C_70 = 10'd112,
    COMP_LOOP_C_71 = 10'd113,
    COMP_LOOP_C_72 = 10'd114,
    COMP_LOOP_C_73 = 10'd115,
    COMP_LOOP_C_74 = 10'd116,
    COMP_LOOP_C_75 = 10'd117,
    COMP_LOOP_C_76 = 10'd118,
    COMP_LOOP_C_77 = 10'd119,
    COMP_LOOP_C_78 = 10'd120,
    COMP_LOOP_C_79 = 10'd121,
    COMP_LOOP_C_80 = 10'd122,
    COMP_LOOP_C_81 = 10'd123,
    COMP_LOOP_C_82 = 10'd124,
    COMP_LOOP_C_83 = 10'd125,
    COMP_LOOP_C_84 = 10'd126,
    COMP_LOOP_C_85 = 10'd127,
    COMP_LOOP_C_86 = 10'd128,
    COMP_LOOP_C_87 = 10'd129,
    COMP_LOOP_C_88 = 10'd130,
    COMP_LOOP_C_89 = 10'd131,
    COMP_LOOP_C_90 = 10'd132,
    COMP_LOOP_C_91 = 10'd133,
    COMP_LOOP_C_92 = 10'd134,
    COMP_LOOP_C_93 = 10'd135,
    COMP_LOOP_C_94 = 10'd136,
    COMP_LOOP_C_95 = 10'd137,
    COMP_LOOP_C_96 = 10'd138,
    COMP_LOOP_C_97 = 10'd139,
    COMP_LOOP_C_98 = 10'd140,
    COMP_LOOP_C_99 = 10'd141,
    COMP_LOOP_C_100 = 10'd142,
    COMP_LOOP_C_101 = 10'd143,
    COMP_LOOP_C_102 = 10'd144,
    COMP_LOOP_C_103 = 10'd145,
    COMP_LOOP_C_104 = 10'd146,
    COMP_LOOP_C_105 = 10'd147,
    COMP_LOOP_C_106 = 10'd148,
    COMP_LOOP_3_modExp_dev_1_while_C_0 = 10'd149,
    COMP_LOOP_3_modExp_dev_1_while_C_1 = 10'd150,
    COMP_LOOP_3_modExp_dev_1_while_C_2 = 10'd151,
    COMP_LOOP_3_modExp_dev_1_while_C_3 = 10'd152,
    COMP_LOOP_3_modExp_dev_1_while_C_4 = 10'd153,
    COMP_LOOP_3_modExp_dev_1_while_C_5 = 10'd154,
    COMP_LOOP_3_modExp_dev_1_while_C_6 = 10'd155,
    COMP_LOOP_3_modExp_dev_1_while_C_7 = 10'd156,
    COMP_LOOP_3_modExp_dev_1_while_C_8 = 10'd157,
    COMP_LOOP_3_modExp_dev_1_while_C_9 = 10'd158,
    COMP_LOOP_3_modExp_dev_1_while_C_10 = 10'd159,
    COMP_LOOP_3_modExp_dev_1_while_C_11 = 10'd160,
    COMP_LOOP_C_107 = 10'd161,
    COMP_LOOP_C_108 = 10'd162,
    COMP_LOOP_C_109 = 10'd163,
    COMP_LOOP_C_110 = 10'd164,
    COMP_LOOP_C_111 = 10'd165,
    COMP_LOOP_C_112 = 10'd166,
    COMP_LOOP_C_113 = 10'd167,
    COMP_LOOP_C_114 = 10'd168,
    COMP_LOOP_C_115 = 10'd169,
    COMP_LOOP_C_116 = 10'd170,
    COMP_LOOP_C_117 = 10'd171,
    COMP_LOOP_C_118 = 10'd172,
    COMP_LOOP_C_119 = 10'd173,
    COMP_LOOP_C_120 = 10'd174,
    COMP_LOOP_C_121 = 10'd175,
    COMP_LOOP_C_122 = 10'd176,
    COMP_LOOP_C_123 = 10'd177,
    COMP_LOOP_C_124 = 10'd178,
    COMP_LOOP_C_125 = 10'd179,
    COMP_LOOP_C_126 = 10'd180,
    COMP_LOOP_C_127 = 10'd181,
    COMP_LOOP_C_128 = 10'd182,
    COMP_LOOP_C_129 = 10'd183,
    COMP_LOOP_C_130 = 10'd184,
    COMP_LOOP_C_131 = 10'd185,
    COMP_LOOP_C_132 = 10'd186,
    COMP_LOOP_C_133 = 10'd187,
    COMP_LOOP_C_134 = 10'd188,
    COMP_LOOP_C_135 = 10'd189,
    COMP_LOOP_C_136 = 10'd190,
    COMP_LOOP_C_137 = 10'd191,
    COMP_LOOP_C_138 = 10'd192,
    COMP_LOOP_C_139 = 10'd193,
    COMP_LOOP_C_140 = 10'd194,
    COMP_LOOP_C_141 = 10'd195,
    COMP_LOOP_C_142 = 10'd196,
    COMP_LOOP_C_143 = 10'd197,
    COMP_LOOP_C_144 = 10'd198,
    COMP_LOOP_C_145 = 10'd199,
    COMP_LOOP_C_146 = 10'd200,
    COMP_LOOP_C_147 = 10'd201,
    COMP_LOOP_C_148 = 10'd202,
    COMP_LOOP_C_149 = 10'd203,
    COMP_LOOP_C_150 = 10'd204,
    COMP_LOOP_C_151 = 10'd205,
    COMP_LOOP_4_modExp_dev_1_while_C_0 = 10'd206,
    COMP_LOOP_4_modExp_dev_1_while_C_1 = 10'd207,
    COMP_LOOP_4_modExp_dev_1_while_C_2 = 10'd208,
    COMP_LOOP_4_modExp_dev_1_while_C_3 = 10'd209,
    COMP_LOOP_4_modExp_dev_1_while_C_4 = 10'd210,
    COMP_LOOP_4_modExp_dev_1_while_C_5 = 10'd211,
    COMP_LOOP_4_modExp_dev_1_while_C_6 = 10'd212,
    COMP_LOOP_4_modExp_dev_1_while_C_7 = 10'd213,
    COMP_LOOP_4_modExp_dev_1_while_C_8 = 10'd214,
    COMP_LOOP_4_modExp_dev_1_while_C_9 = 10'd215,
    COMP_LOOP_4_modExp_dev_1_while_C_10 = 10'd216,
    COMP_LOOP_4_modExp_dev_1_while_C_11 = 10'd217,
    COMP_LOOP_C_152 = 10'd218,
    COMP_LOOP_C_153 = 10'd219,
    COMP_LOOP_C_154 = 10'd220,
    COMP_LOOP_C_155 = 10'd221,
    COMP_LOOP_C_156 = 10'd222,
    COMP_LOOP_C_157 = 10'd223,
    COMP_LOOP_C_158 = 10'd224,
    COMP_LOOP_C_159 = 10'd225,
    COMP_LOOP_C_160 = 10'd226,
    COMP_LOOP_C_161 = 10'd227,
    COMP_LOOP_C_162 = 10'd228,
    COMP_LOOP_C_163 = 10'd229,
    COMP_LOOP_C_164 = 10'd230,
    COMP_LOOP_C_165 = 10'd231,
    COMP_LOOP_C_166 = 10'd232,
    COMP_LOOP_C_167 = 10'd233,
    COMP_LOOP_C_168 = 10'd234,
    COMP_LOOP_C_169 = 10'd235,
    COMP_LOOP_C_170 = 10'd236,
    COMP_LOOP_C_171 = 10'd237,
    COMP_LOOP_C_172 = 10'd238,
    COMP_LOOP_C_173 = 10'd239,
    COMP_LOOP_C_174 = 10'd240,
    COMP_LOOP_C_175 = 10'd241,
    COMP_LOOP_C_176 = 10'd242,
    COMP_LOOP_C_177 = 10'd243,
    COMP_LOOP_C_178 = 10'd244,
    COMP_LOOP_C_179 = 10'd245,
    COMP_LOOP_C_180 = 10'd246,
    COMP_LOOP_C_181 = 10'd247,
    COMP_LOOP_C_182 = 10'd248,
    COMP_LOOP_C_183 = 10'd249,
    COMP_LOOP_C_184 = 10'd250,
    COMP_LOOP_C_185 = 10'd251,
    COMP_LOOP_C_186 = 10'd252,
    COMP_LOOP_C_187 = 10'd253,
    COMP_LOOP_C_188 = 10'd254,
    COMP_LOOP_C_189 = 10'd255,
    COMP_LOOP_C_190 = 10'd256,
    COMP_LOOP_C_191 = 10'd257,
    COMP_LOOP_C_192 = 10'd258,
    COMP_LOOP_C_193 = 10'd259,
    COMP_LOOP_C_194 = 10'd260,
    COMP_LOOP_C_195 = 10'd261,
    COMP_LOOP_C_196 = 10'd262,
    COMP_LOOP_5_modExp_dev_1_while_C_0 = 10'd263,
    COMP_LOOP_5_modExp_dev_1_while_C_1 = 10'd264,
    COMP_LOOP_5_modExp_dev_1_while_C_2 = 10'd265,
    COMP_LOOP_5_modExp_dev_1_while_C_3 = 10'd266,
    COMP_LOOP_5_modExp_dev_1_while_C_4 = 10'd267,
    COMP_LOOP_5_modExp_dev_1_while_C_5 = 10'd268,
    COMP_LOOP_5_modExp_dev_1_while_C_6 = 10'd269,
    COMP_LOOP_5_modExp_dev_1_while_C_7 = 10'd270,
    COMP_LOOP_5_modExp_dev_1_while_C_8 = 10'd271,
    COMP_LOOP_5_modExp_dev_1_while_C_9 = 10'd272,
    COMP_LOOP_5_modExp_dev_1_while_C_10 = 10'd273,
    COMP_LOOP_5_modExp_dev_1_while_C_11 = 10'd274,
    COMP_LOOP_C_197 = 10'd275,
    COMP_LOOP_C_198 = 10'd276,
    COMP_LOOP_C_199 = 10'd277,
    COMP_LOOP_C_200 = 10'd278,
    COMP_LOOP_C_201 = 10'd279,
    COMP_LOOP_C_202 = 10'd280,
    COMP_LOOP_C_203 = 10'd281,
    COMP_LOOP_C_204 = 10'd282,
    COMP_LOOP_C_205 = 10'd283,
    COMP_LOOP_C_206 = 10'd284,
    COMP_LOOP_C_207 = 10'd285,
    COMP_LOOP_C_208 = 10'd286,
    COMP_LOOP_C_209 = 10'd287,
    COMP_LOOP_C_210 = 10'd288,
    COMP_LOOP_C_211 = 10'd289,
    COMP_LOOP_C_212 = 10'd290,
    COMP_LOOP_C_213 = 10'd291,
    COMP_LOOP_C_214 = 10'd292,
    COMP_LOOP_C_215 = 10'd293,
    COMP_LOOP_C_216 = 10'd294,
    COMP_LOOP_C_217 = 10'd295,
    COMP_LOOP_C_218 = 10'd296,
    COMP_LOOP_C_219 = 10'd297,
    COMP_LOOP_C_220 = 10'd298,
    COMP_LOOP_C_221 = 10'd299,
    COMP_LOOP_C_222 = 10'd300,
    COMP_LOOP_C_223 = 10'd301,
    COMP_LOOP_C_224 = 10'd302,
    COMP_LOOP_C_225 = 10'd303,
    COMP_LOOP_C_226 = 10'd304,
    COMP_LOOP_C_227 = 10'd305,
    COMP_LOOP_C_228 = 10'd306,
    COMP_LOOP_C_229 = 10'd307,
    COMP_LOOP_C_230 = 10'd308,
    COMP_LOOP_C_231 = 10'd309,
    COMP_LOOP_C_232 = 10'd310,
    COMP_LOOP_C_233 = 10'd311,
    COMP_LOOP_C_234 = 10'd312,
    COMP_LOOP_C_235 = 10'd313,
    COMP_LOOP_C_236 = 10'd314,
    COMP_LOOP_C_237 = 10'd315,
    COMP_LOOP_C_238 = 10'd316,
    COMP_LOOP_C_239 = 10'd317,
    COMP_LOOP_C_240 = 10'd318,
    COMP_LOOP_C_241 = 10'd319,
    COMP_LOOP_6_modExp_dev_1_while_C_0 = 10'd320,
    COMP_LOOP_6_modExp_dev_1_while_C_1 = 10'd321,
    COMP_LOOP_6_modExp_dev_1_while_C_2 = 10'd322,
    COMP_LOOP_6_modExp_dev_1_while_C_3 = 10'd323,
    COMP_LOOP_6_modExp_dev_1_while_C_4 = 10'd324,
    COMP_LOOP_6_modExp_dev_1_while_C_5 = 10'd325,
    COMP_LOOP_6_modExp_dev_1_while_C_6 = 10'd326,
    COMP_LOOP_6_modExp_dev_1_while_C_7 = 10'd327,
    COMP_LOOP_6_modExp_dev_1_while_C_8 = 10'd328,
    COMP_LOOP_6_modExp_dev_1_while_C_9 = 10'd329,
    COMP_LOOP_6_modExp_dev_1_while_C_10 = 10'd330,
    COMP_LOOP_6_modExp_dev_1_while_C_11 = 10'd331,
    COMP_LOOP_C_242 = 10'd332,
    COMP_LOOP_C_243 = 10'd333,
    COMP_LOOP_C_244 = 10'd334,
    COMP_LOOP_C_245 = 10'd335,
    COMP_LOOP_C_246 = 10'd336,
    COMP_LOOP_C_247 = 10'd337,
    COMP_LOOP_C_248 = 10'd338,
    COMP_LOOP_C_249 = 10'd339,
    COMP_LOOP_C_250 = 10'd340,
    COMP_LOOP_C_251 = 10'd341,
    COMP_LOOP_C_252 = 10'd342,
    COMP_LOOP_C_253 = 10'd343,
    COMP_LOOP_C_254 = 10'd344,
    COMP_LOOP_C_255 = 10'd345,
    COMP_LOOP_C_256 = 10'd346,
    COMP_LOOP_C_257 = 10'd347,
    COMP_LOOP_C_258 = 10'd348,
    COMP_LOOP_C_259 = 10'd349,
    COMP_LOOP_C_260 = 10'd350,
    COMP_LOOP_C_261 = 10'd351,
    COMP_LOOP_C_262 = 10'd352,
    COMP_LOOP_C_263 = 10'd353,
    COMP_LOOP_C_264 = 10'd354,
    COMP_LOOP_C_265 = 10'd355,
    COMP_LOOP_C_266 = 10'd356,
    COMP_LOOP_C_267 = 10'd357,
    COMP_LOOP_C_268 = 10'd358,
    COMP_LOOP_C_269 = 10'd359,
    COMP_LOOP_C_270 = 10'd360,
    COMP_LOOP_C_271 = 10'd361,
    COMP_LOOP_C_272 = 10'd362,
    COMP_LOOP_C_273 = 10'd363,
    COMP_LOOP_C_274 = 10'd364,
    COMP_LOOP_C_275 = 10'd365,
    COMP_LOOP_C_276 = 10'd366,
    COMP_LOOP_C_277 = 10'd367,
    COMP_LOOP_C_278 = 10'd368,
    COMP_LOOP_C_279 = 10'd369,
    COMP_LOOP_C_280 = 10'd370,
    COMP_LOOP_C_281 = 10'd371,
    COMP_LOOP_C_282 = 10'd372,
    COMP_LOOP_C_283 = 10'd373,
    COMP_LOOP_C_284 = 10'd374,
    COMP_LOOP_C_285 = 10'd375,
    COMP_LOOP_C_286 = 10'd376,
    COMP_LOOP_7_modExp_dev_1_while_C_0 = 10'd377,
    COMP_LOOP_7_modExp_dev_1_while_C_1 = 10'd378,
    COMP_LOOP_7_modExp_dev_1_while_C_2 = 10'd379,
    COMP_LOOP_7_modExp_dev_1_while_C_3 = 10'd380,
    COMP_LOOP_7_modExp_dev_1_while_C_4 = 10'd381,
    COMP_LOOP_7_modExp_dev_1_while_C_5 = 10'd382,
    COMP_LOOP_7_modExp_dev_1_while_C_6 = 10'd383,
    COMP_LOOP_7_modExp_dev_1_while_C_7 = 10'd384,
    COMP_LOOP_7_modExp_dev_1_while_C_8 = 10'd385,
    COMP_LOOP_7_modExp_dev_1_while_C_9 = 10'd386,
    COMP_LOOP_7_modExp_dev_1_while_C_10 = 10'd387,
    COMP_LOOP_7_modExp_dev_1_while_C_11 = 10'd388,
    COMP_LOOP_C_287 = 10'd389,
    COMP_LOOP_C_288 = 10'd390,
    COMP_LOOP_C_289 = 10'd391,
    COMP_LOOP_C_290 = 10'd392,
    COMP_LOOP_C_291 = 10'd393,
    COMP_LOOP_C_292 = 10'd394,
    COMP_LOOP_C_293 = 10'd395,
    COMP_LOOP_C_294 = 10'd396,
    COMP_LOOP_C_295 = 10'd397,
    COMP_LOOP_C_296 = 10'd398,
    COMP_LOOP_C_297 = 10'd399,
    COMP_LOOP_C_298 = 10'd400,
    COMP_LOOP_C_299 = 10'd401,
    COMP_LOOP_C_300 = 10'd402,
    COMP_LOOP_C_301 = 10'd403,
    COMP_LOOP_C_302 = 10'd404,
    COMP_LOOP_C_303 = 10'd405,
    COMP_LOOP_C_304 = 10'd406,
    COMP_LOOP_C_305 = 10'd407,
    COMP_LOOP_C_306 = 10'd408,
    COMP_LOOP_C_307 = 10'd409,
    COMP_LOOP_C_308 = 10'd410,
    COMP_LOOP_C_309 = 10'd411,
    COMP_LOOP_C_310 = 10'd412,
    COMP_LOOP_C_311 = 10'd413,
    COMP_LOOP_C_312 = 10'd414,
    COMP_LOOP_C_313 = 10'd415,
    COMP_LOOP_C_314 = 10'd416,
    COMP_LOOP_C_315 = 10'd417,
    COMP_LOOP_C_316 = 10'd418,
    COMP_LOOP_C_317 = 10'd419,
    COMP_LOOP_C_318 = 10'd420,
    COMP_LOOP_C_319 = 10'd421,
    COMP_LOOP_C_320 = 10'd422,
    COMP_LOOP_C_321 = 10'd423,
    COMP_LOOP_C_322 = 10'd424,
    COMP_LOOP_C_323 = 10'd425,
    COMP_LOOP_C_324 = 10'd426,
    COMP_LOOP_C_325 = 10'd427,
    COMP_LOOP_C_326 = 10'd428,
    COMP_LOOP_C_327 = 10'd429,
    COMP_LOOP_C_328 = 10'd430,
    COMP_LOOP_C_329 = 10'd431,
    COMP_LOOP_C_330 = 10'd432,
    COMP_LOOP_C_331 = 10'd433,
    COMP_LOOP_8_modExp_dev_1_while_C_0 = 10'd434,
    COMP_LOOP_8_modExp_dev_1_while_C_1 = 10'd435,
    COMP_LOOP_8_modExp_dev_1_while_C_2 = 10'd436,
    COMP_LOOP_8_modExp_dev_1_while_C_3 = 10'd437,
    COMP_LOOP_8_modExp_dev_1_while_C_4 = 10'd438,
    COMP_LOOP_8_modExp_dev_1_while_C_5 = 10'd439,
    COMP_LOOP_8_modExp_dev_1_while_C_6 = 10'd440,
    COMP_LOOP_8_modExp_dev_1_while_C_7 = 10'd441,
    COMP_LOOP_8_modExp_dev_1_while_C_8 = 10'd442,
    COMP_LOOP_8_modExp_dev_1_while_C_9 = 10'd443,
    COMP_LOOP_8_modExp_dev_1_while_C_10 = 10'd444,
    COMP_LOOP_8_modExp_dev_1_while_C_11 = 10'd445,
    COMP_LOOP_C_332 = 10'd446,
    COMP_LOOP_C_333 = 10'd447,
    COMP_LOOP_C_334 = 10'd448,
    COMP_LOOP_C_335 = 10'd449,
    COMP_LOOP_C_336 = 10'd450,
    COMP_LOOP_C_337 = 10'd451,
    COMP_LOOP_C_338 = 10'd452,
    COMP_LOOP_C_339 = 10'd453,
    COMP_LOOP_C_340 = 10'd454,
    COMP_LOOP_C_341 = 10'd455,
    COMP_LOOP_C_342 = 10'd456,
    COMP_LOOP_C_343 = 10'd457,
    COMP_LOOP_C_344 = 10'd458,
    COMP_LOOP_C_345 = 10'd459,
    COMP_LOOP_C_346 = 10'd460,
    COMP_LOOP_C_347 = 10'd461,
    COMP_LOOP_C_348 = 10'd462,
    COMP_LOOP_C_349 = 10'd463,
    COMP_LOOP_C_350 = 10'd464,
    COMP_LOOP_C_351 = 10'd465,
    COMP_LOOP_C_352 = 10'd466,
    COMP_LOOP_C_353 = 10'd467,
    COMP_LOOP_C_354 = 10'd468,
    COMP_LOOP_C_355 = 10'd469,
    COMP_LOOP_C_356 = 10'd470,
    COMP_LOOP_C_357 = 10'd471,
    COMP_LOOP_C_358 = 10'd472,
    COMP_LOOP_C_359 = 10'd473,
    COMP_LOOP_C_360 = 10'd474,
    COMP_LOOP_C_361 = 10'd475,
    COMP_LOOP_C_362 = 10'd476,
    COMP_LOOP_C_363 = 10'd477,
    COMP_LOOP_C_364 = 10'd478,
    COMP_LOOP_C_365 = 10'd479,
    COMP_LOOP_C_366 = 10'd480,
    COMP_LOOP_C_367 = 10'd481,
    COMP_LOOP_C_368 = 10'd482,
    COMP_LOOP_C_369 = 10'd483,
    COMP_LOOP_C_370 = 10'd484,
    COMP_LOOP_C_371 = 10'd485,
    COMP_LOOP_C_372 = 10'd486,
    COMP_LOOP_C_373 = 10'd487,
    COMP_LOOP_C_374 = 10'd488,
    COMP_LOOP_C_375 = 10'd489,
    COMP_LOOP_C_376 = 10'd490,
    COMP_LOOP_9_modExp_dev_1_while_C_0 = 10'd491,
    COMP_LOOP_9_modExp_dev_1_while_C_1 = 10'd492,
    COMP_LOOP_9_modExp_dev_1_while_C_2 = 10'd493,
    COMP_LOOP_9_modExp_dev_1_while_C_3 = 10'd494,
    COMP_LOOP_9_modExp_dev_1_while_C_4 = 10'd495,
    COMP_LOOP_9_modExp_dev_1_while_C_5 = 10'd496,
    COMP_LOOP_9_modExp_dev_1_while_C_6 = 10'd497,
    COMP_LOOP_9_modExp_dev_1_while_C_7 = 10'd498,
    COMP_LOOP_9_modExp_dev_1_while_C_8 = 10'd499,
    COMP_LOOP_9_modExp_dev_1_while_C_9 = 10'd500,
    COMP_LOOP_9_modExp_dev_1_while_C_10 = 10'd501,
    COMP_LOOP_9_modExp_dev_1_while_C_11 = 10'd502,
    COMP_LOOP_C_377 = 10'd503,
    COMP_LOOP_C_378 = 10'd504,
    COMP_LOOP_C_379 = 10'd505,
    COMP_LOOP_C_380 = 10'd506,
    COMP_LOOP_C_381 = 10'd507,
    COMP_LOOP_C_382 = 10'd508,
    COMP_LOOP_C_383 = 10'd509,
    COMP_LOOP_C_384 = 10'd510,
    COMP_LOOP_C_385 = 10'd511,
    COMP_LOOP_C_386 = 10'd512,
    COMP_LOOP_C_387 = 10'd513,
    COMP_LOOP_C_388 = 10'd514,
    COMP_LOOP_C_389 = 10'd515,
    COMP_LOOP_C_390 = 10'd516,
    COMP_LOOP_C_391 = 10'd517,
    COMP_LOOP_C_392 = 10'd518,
    COMP_LOOP_C_393 = 10'd519,
    COMP_LOOP_C_394 = 10'd520,
    COMP_LOOP_C_395 = 10'd521,
    COMP_LOOP_C_396 = 10'd522,
    COMP_LOOP_C_397 = 10'd523,
    COMP_LOOP_C_398 = 10'd524,
    COMP_LOOP_C_399 = 10'd525,
    COMP_LOOP_C_400 = 10'd526,
    COMP_LOOP_C_401 = 10'd527,
    COMP_LOOP_C_402 = 10'd528,
    COMP_LOOP_C_403 = 10'd529,
    COMP_LOOP_C_404 = 10'd530,
    COMP_LOOP_C_405 = 10'd531,
    COMP_LOOP_C_406 = 10'd532,
    COMP_LOOP_C_407 = 10'd533,
    COMP_LOOP_C_408 = 10'd534,
    COMP_LOOP_C_409 = 10'd535,
    COMP_LOOP_C_410 = 10'd536,
    COMP_LOOP_C_411 = 10'd537,
    COMP_LOOP_C_412 = 10'd538,
    COMP_LOOP_C_413 = 10'd539,
    COMP_LOOP_C_414 = 10'd540,
    COMP_LOOP_C_415 = 10'd541,
    COMP_LOOP_C_416 = 10'd542,
    COMP_LOOP_C_417 = 10'd543,
    COMP_LOOP_C_418 = 10'd544,
    COMP_LOOP_C_419 = 10'd545,
    COMP_LOOP_C_420 = 10'd546,
    COMP_LOOP_C_421 = 10'd547,
    COMP_LOOP_10_modExp_dev_1_while_C_0 = 10'd548,
    COMP_LOOP_10_modExp_dev_1_while_C_1 = 10'd549,
    COMP_LOOP_10_modExp_dev_1_while_C_2 = 10'd550,
    COMP_LOOP_10_modExp_dev_1_while_C_3 = 10'd551,
    COMP_LOOP_10_modExp_dev_1_while_C_4 = 10'd552,
    COMP_LOOP_10_modExp_dev_1_while_C_5 = 10'd553,
    COMP_LOOP_10_modExp_dev_1_while_C_6 = 10'd554,
    COMP_LOOP_10_modExp_dev_1_while_C_7 = 10'd555,
    COMP_LOOP_10_modExp_dev_1_while_C_8 = 10'd556,
    COMP_LOOP_10_modExp_dev_1_while_C_9 = 10'd557,
    COMP_LOOP_10_modExp_dev_1_while_C_10 = 10'd558,
    COMP_LOOP_10_modExp_dev_1_while_C_11 = 10'd559,
    COMP_LOOP_C_422 = 10'd560,
    COMP_LOOP_C_423 = 10'd561,
    COMP_LOOP_C_424 = 10'd562,
    COMP_LOOP_C_425 = 10'd563,
    COMP_LOOP_C_426 = 10'd564,
    COMP_LOOP_C_427 = 10'd565,
    COMP_LOOP_C_428 = 10'd566,
    COMP_LOOP_C_429 = 10'd567,
    COMP_LOOP_C_430 = 10'd568,
    COMP_LOOP_C_431 = 10'd569,
    COMP_LOOP_C_432 = 10'd570,
    COMP_LOOP_C_433 = 10'd571,
    COMP_LOOP_C_434 = 10'd572,
    COMP_LOOP_C_435 = 10'd573,
    COMP_LOOP_C_436 = 10'd574,
    COMP_LOOP_C_437 = 10'd575,
    COMP_LOOP_C_438 = 10'd576,
    COMP_LOOP_C_439 = 10'd577,
    COMP_LOOP_C_440 = 10'd578,
    COMP_LOOP_C_441 = 10'd579,
    COMP_LOOP_C_442 = 10'd580,
    COMP_LOOP_C_443 = 10'd581,
    COMP_LOOP_C_444 = 10'd582,
    COMP_LOOP_C_445 = 10'd583,
    COMP_LOOP_C_446 = 10'd584,
    COMP_LOOP_C_447 = 10'd585,
    COMP_LOOP_C_448 = 10'd586,
    COMP_LOOP_C_449 = 10'd587,
    COMP_LOOP_C_450 = 10'd588,
    COMP_LOOP_C_451 = 10'd589,
    COMP_LOOP_C_452 = 10'd590,
    COMP_LOOP_C_453 = 10'd591,
    COMP_LOOP_C_454 = 10'd592,
    COMP_LOOP_C_455 = 10'd593,
    COMP_LOOP_C_456 = 10'd594,
    COMP_LOOP_C_457 = 10'd595,
    COMP_LOOP_C_458 = 10'd596,
    COMP_LOOP_C_459 = 10'd597,
    COMP_LOOP_C_460 = 10'd598,
    COMP_LOOP_C_461 = 10'd599,
    COMP_LOOP_C_462 = 10'd600,
    COMP_LOOP_C_463 = 10'd601,
    COMP_LOOP_C_464 = 10'd602,
    COMP_LOOP_C_465 = 10'd603,
    COMP_LOOP_C_466 = 10'd604,
    COMP_LOOP_11_modExp_dev_1_while_C_0 = 10'd605,
    COMP_LOOP_11_modExp_dev_1_while_C_1 = 10'd606,
    COMP_LOOP_11_modExp_dev_1_while_C_2 = 10'd607,
    COMP_LOOP_11_modExp_dev_1_while_C_3 = 10'd608,
    COMP_LOOP_11_modExp_dev_1_while_C_4 = 10'd609,
    COMP_LOOP_11_modExp_dev_1_while_C_5 = 10'd610,
    COMP_LOOP_11_modExp_dev_1_while_C_6 = 10'd611,
    COMP_LOOP_11_modExp_dev_1_while_C_7 = 10'd612,
    COMP_LOOP_11_modExp_dev_1_while_C_8 = 10'd613,
    COMP_LOOP_11_modExp_dev_1_while_C_9 = 10'd614,
    COMP_LOOP_11_modExp_dev_1_while_C_10 = 10'd615,
    COMP_LOOP_11_modExp_dev_1_while_C_11 = 10'd616,
    COMP_LOOP_C_467 = 10'd617,
    COMP_LOOP_C_468 = 10'd618,
    COMP_LOOP_C_469 = 10'd619,
    COMP_LOOP_C_470 = 10'd620,
    COMP_LOOP_C_471 = 10'd621,
    COMP_LOOP_C_472 = 10'd622,
    COMP_LOOP_C_473 = 10'd623,
    COMP_LOOP_C_474 = 10'd624,
    COMP_LOOP_C_475 = 10'd625,
    COMP_LOOP_C_476 = 10'd626,
    COMP_LOOP_C_477 = 10'd627,
    COMP_LOOP_C_478 = 10'd628,
    COMP_LOOP_C_479 = 10'd629,
    COMP_LOOP_C_480 = 10'd630,
    COMP_LOOP_C_481 = 10'd631,
    COMP_LOOP_C_482 = 10'd632,
    COMP_LOOP_C_483 = 10'd633,
    COMP_LOOP_C_484 = 10'd634,
    COMP_LOOP_C_485 = 10'd635,
    COMP_LOOP_C_486 = 10'd636,
    COMP_LOOP_C_487 = 10'd637,
    COMP_LOOP_C_488 = 10'd638,
    COMP_LOOP_C_489 = 10'd639,
    COMP_LOOP_C_490 = 10'd640,
    COMP_LOOP_C_491 = 10'd641,
    COMP_LOOP_C_492 = 10'd642,
    COMP_LOOP_C_493 = 10'd643,
    COMP_LOOP_C_494 = 10'd644,
    COMP_LOOP_C_495 = 10'd645,
    COMP_LOOP_C_496 = 10'd646,
    COMP_LOOP_C_497 = 10'd647,
    COMP_LOOP_C_498 = 10'd648,
    COMP_LOOP_C_499 = 10'd649,
    COMP_LOOP_C_500 = 10'd650,
    COMP_LOOP_C_501 = 10'd651,
    COMP_LOOP_C_502 = 10'd652,
    COMP_LOOP_C_503 = 10'd653,
    COMP_LOOP_C_504 = 10'd654,
    COMP_LOOP_C_505 = 10'd655,
    COMP_LOOP_C_506 = 10'd656,
    COMP_LOOP_C_507 = 10'd657,
    COMP_LOOP_C_508 = 10'd658,
    COMP_LOOP_C_509 = 10'd659,
    COMP_LOOP_C_510 = 10'd660,
    COMP_LOOP_C_511 = 10'd661,
    COMP_LOOP_12_modExp_dev_1_while_C_0 = 10'd662,
    COMP_LOOP_12_modExp_dev_1_while_C_1 = 10'd663,
    COMP_LOOP_12_modExp_dev_1_while_C_2 = 10'd664,
    COMP_LOOP_12_modExp_dev_1_while_C_3 = 10'd665,
    COMP_LOOP_12_modExp_dev_1_while_C_4 = 10'd666,
    COMP_LOOP_12_modExp_dev_1_while_C_5 = 10'd667,
    COMP_LOOP_12_modExp_dev_1_while_C_6 = 10'd668,
    COMP_LOOP_12_modExp_dev_1_while_C_7 = 10'd669,
    COMP_LOOP_12_modExp_dev_1_while_C_8 = 10'd670,
    COMP_LOOP_12_modExp_dev_1_while_C_9 = 10'd671,
    COMP_LOOP_12_modExp_dev_1_while_C_10 = 10'd672,
    COMP_LOOP_12_modExp_dev_1_while_C_11 = 10'd673,
    COMP_LOOP_C_512 = 10'd674,
    COMP_LOOP_C_513 = 10'd675,
    COMP_LOOP_C_514 = 10'd676,
    COMP_LOOP_C_515 = 10'd677,
    COMP_LOOP_C_516 = 10'd678,
    COMP_LOOP_C_517 = 10'd679,
    COMP_LOOP_C_518 = 10'd680,
    COMP_LOOP_C_519 = 10'd681,
    COMP_LOOP_C_520 = 10'd682,
    COMP_LOOP_C_521 = 10'd683,
    COMP_LOOP_C_522 = 10'd684,
    COMP_LOOP_C_523 = 10'd685,
    COMP_LOOP_C_524 = 10'd686,
    COMP_LOOP_C_525 = 10'd687,
    COMP_LOOP_C_526 = 10'd688,
    COMP_LOOP_C_527 = 10'd689,
    COMP_LOOP_C_528 = 10'd690,
    COMP_LOOP_C_529 = 10'd691,
    COMP_LOOP_C_530 = 10'd692,
    COMP_LOOP_C_531 = 10'd693,
    COMP_LOOP_C_532 = 10'd694,
    COMP_LOOP_C_533 = 10'd695,
    COMP_LOOP_C_534 = 10'd696,
    COMP_LOOP_C_535 = 10'd697,
    COMP_LOOP_C_536 = 10'd698,
    COMP_LOOP_C_537 = 10'd699,
    COMP_LOOP_C_538 = 10'd700,
    COMP_LOOP_C_539 = 10'd701,
    COMP_LOOP_C_540 = 10'd702,
    COMP_LOOP_C_541 = 10'd703,
    COMP_LOOP_C_542 = 10'd704,
    COMP_LOOP_C_543 = 10'd705,
    COMP_LOOP_C_544 = 10'd706,
    COMP_LOOP_C_545 = 10'd707,
    COMP_LOOP_C_546 = 10'd708,
    COMP_LOOP_C_547 = 10'd709,
    COMP_LOOP_C_548 = 10'd710,
    COMP_LOOP_C_549 = 10'd711,
    COMP_LOOP_C_550 = 10'd712,
    COMP_LOOP_C_551 = 10'd713,
    COMP_LOOP_C_552 = 10'd714,
    COMP_LOOP_C_553 = 10'd715,
    COMP_LOOP_C_554 = 10'd716,
    COMP_LOOP_C_555 = 10'd717,
    COMP_LOOP_C_556 = 10'd718,
    COMP_LOOP_13_modExp_dev_1_while_C_0 = 10'd719,
    COMP_LOOP_13_modExp_dev_1_while_C_1 = 10'd720,
    COMP_LOOP_13_modExp_dev_1_while_C_2 = 10'd721,
    COMP_LOOP_13_modExp_dev_1_while_C_3 = 10'd722,
    COMP_LOOP_13_modExp_dev_1_while_C_4 = 10'd723,
    COMP_LOOP_13_modExp_dev_1_while_C_5 = 10'd724,
    COMP_LOOP_13_modExp_dev_1_while_C_6 = 10'd725,
    COMP_LOOP_13_modExp_dev_1_while_C_7 = 10'd726,
    COMP_LOOP_13_modExp_dev_1_while_C_8 = 10'd727,
    COMP_LOOP_13_modExp_dev_1_while_C_9 = 10'd728,
    COMP_LOOP_13_modExp_dev_1_while_C_10 = 10'd729,
    COMP_LOOP_13_modExp_dev_1_while_C_11 = 10'd730,
    COMP_LOOP_C_557 = 10'd731,
    COMP_LOOP_C_558 = 10'd732,
    COMP_LOOP_C_559 = 10'd733,
    COMP_LOOP_C_560 = 10'd734,
    COMP_LOOP_C_561 = 10'd735,
    COMP_LOOP_C_562 = 10'd736,
    COMP_LOOP_C_563 = 10'd737,
    COMP_LOOP_C_564 = 10'd738,
    COMP_LOOP_C_565 = 10'd739,
    COMP_LOOP_C_566 = 10'd740,
    COMP_LOOP_C_567 = 10'd741,
    COMP_LOOP_C_568 = 10'd742,
    COMP_LOOP_C_569 = 10'd743,
    COMP_LOOP_C_570 = 10'd744,
    COMP_LOOP_C_571 = 10'd745,
    COMP_LOOP_C_572 = 10'd746,
    COMP_LOOP_C_573 = 10'd747,
    COMP_LOOP_C_574 = 10'd748,
    COMP_LOOP_C_575 = 10'd749,
    COMP_LOOP_C_576 = 10'd750,
    COMP_LOOP_C_577 = 10'd751,
    COMP_LOOP_C_578 = 10'd752,
    COMP_LOOP_C_579 = 10'd753,
    COMP_LOOP_C_580 = 10'd754,
    COMP_LOOP_C_581 = 10'd755,
    COMP_LOOP_C_582 = 10'd756,
    COMP_LOOP_C_583 = 10'd757,
    COMP_LOOP_C_584 = 10'd758,
    COMP_LOOP_C_585 = 10'd759,
    COMP_LOOP_C_586 = 10'd760,
    COMP_LOOP_C_587 = 10'd761,
    COMP_LOOP_C_588 = 10'd762,
    COMP_LOOP_C_589 = 10'd763,
    COMP_LOOP_C_590 = 10'd764,
    COMP_LOOP_C_591 = 10'd765,
    COMP_LOOP_C_592 = 10'd766,
    COMP_LOOP_C_593 = 10'd767,
    COMP_LOOP_C_594 = 10'd768,
    COMP_LOOP_C_595 = 10'd769,
    COMP_LOOP_C_596 = 10'd770,
    COMP_LOOP_C_597 = 10'd771,
    COMP_LOOP_C_598 = 10'd772,
    COMP_LOOP_C_599 = 10'd773,
    COMP_LOOP_C_600 = 10'd774,
    COMP_LOOP_C_601 = 10'd775,
    COMP_LOOP_14_modExp_dev_1_while_C_0 = 10'd776,
    COMP_LOOP_14_modExp_dev_1_while_C_1 = 10'd777,
    COMP_LOOP_14_modExp_dev_1_while_C_2 = 10'd778,
    COMP_LOOP_14_modExp_dev_1_while_C_3 = 10'd779,
    COMP_LOOP_14_modExp_dev_1_while_C_4 = 10'd780,
    COMP_LOOP_14_modExp_dev_1_while_C_5 = 10'd781,
    COMP_LOOP_14_modExp_dev_1_while_C_6 = 10'd782,
    COMP_LOOP_14_modExp_dev_1_while_C_7 = 10'd783,
    COMP_LOOP_14_modExp_dev_1_while_C_8 = 10'd784,
    COMP_LOOP_14_modExp_dev_1_while_C_9 = 10'd785,
    COMP_LOOP_14_modExp_dev_1_while_C_10 = 10'd786,
    COMP_LOOP_14_modExp_dev_1_while_C_11 = 10'd787,
    COMP_LOOP_C_602 = 10'd788,
    COMP_LOOP_C_603 = 10'd789,
    COMP_LOOP_C_604 = 10'd790,
    COMP_LOOP_C_605 = 10'd791,
    COMP_LOOP_C_606 = 10'd792,
    COMP_LOOP_C_607 = 10'd793,
    COMP_LOOP_C_608 = 10'd794,
    COMP_LOOP_C_609 = 10'd795,
    COMP_LOOP_C_610 = 10'd796,
    COMP_LOOP_C_611 = 10'd797,
    COMP_LOOP_C_612 = 10'd798,
    COMP_LOOP_C_613 = 10'd799,
    COMP_LOOP_C_614 = 10'd800,
    COMP_LOOP_C_615 = 10'd801,
    COMP_LOOP_C_616 = 10'd802,
    COMP_LOOP_C_617 = 10'd803,
    COMP_LOOP_C_618 = 10'd804,
    COMP_LOOP_C_619 = 10'd805,
    COMP_LOOP_C_620 = 10'd806,
    COMP_LOOP_C_621 = 10'd807,
    COMP_LOOP_C_622 = 10'd808,
    COMP_LOOP_C_623 = 10'd809,
    COMP_LOOP_C_624 = 10'd810,
    COMP_LOOP_C_625 = 10'd811,
    COMP_LOOP_C_626 = 10'd812,
    COMP_LOOP_C_627 = 10'd813,
    COMP_LOOP_C_628 = 10'd814,
    COMP_LOOP_C_629 = 10'd815,
    COMP_LOOP_C_630 = 10'd816,
    COMP_LOOP_C_631 = 10'd817,
    COMP_LOOP_C_632 = 10'd818,
    COMP_LOOP_C_633 = 10'd819,
    COMP_LOOP_C_634 = 10'd820,
    COMP_LOOP_C_635 = 10'd821,
    COMP_LOOP_C_636 = 10'd822,
    COMP_LOOP_C_637 = 10'd823,
    COMP_LOOP_C_638 = 10'd824,
    COMP_LOOP_C_639 = 10'd825,
    COMP_LOOP_C_640 = 10'd826,
    COMP_LOOP_C_641 = 10'd827,
    COMP_LOOP_C_642 = 10'd828,
    COMP_LOOP_C_643 = 10'd829,
    COMP_LOOP_C_644 = 10'd830,
    COMP_LOOP_C_645 = 10'd831,
    COMP_LOOP_C_646 = 10'd832,
    COMP_LOOP_15_modExp_dev_1_while_C_0 = 10'd833,
    COMP_LOOP_15_modExp_dev_1_while_C_1 = 10'd834,
    COMP_LOOP_15_modExp_dev_1_while_C_2 = 10'd835,
    COMP_LOOP_15_modExp_dev_1_while_C_3 = 10'd836,
    COMP_LOOP_15_modExp_dev_1_while_C_4 = 10'd837,
    COMP_LOOP_15_modExp_dev_1_while_C_5 = 10'd838,
    COMP_LOOP_15_modExp_dev_1_while_C_6 = 10'd839,
    COMP_LOOP_15_modExp_dev_1_while_C_7 = 10'd840,
    COMP_LOOP_15_modExp_dev_1_while_C_8 = 10'd841,
    COMP_LOOP_15_modExp_dev_1_while_C_9 = 10'd842,
    COMP_LOOP_15_modExp_dev_1_while_C_10 = 10'd843,
    COMP_LOOP_15_modExp_dev_1_while_C_11 = 10'd844,
    COMP_LOOP_C_647 = 10'd845,
    COMP_LOOP_C_648 = 10'd846,
    COMP_LOOP_C_649 = 10'd847,
    COMP_LOOP_C_650 = 10'd848,
    COMP_LOOP_C_651 = 10'd849,
    COMP_LOOP_C_652 = 10'd850,
    COMP_LOOP_C_653 = 10'd851,
    COMP_LOOP_C_654 = 10'd852,
    COMP_LOOP_C_655 = 10'd853,
    COMP_LOOP_C_656 = 10'd854,
    COMP_LOOP_C_657 = 10'd855,
    COMP_LOOP_C_658 = 10'd856,
    COMP_LOOP_C_659 = 10'd857,
    COMP_LOOP_C_660 = 10'd858,
    COMP_LOOP_C_661 = 10'd859,
    COMP_LOOP_C_662 = 10'd860,
    COMP_LOOP_C_663 = 10'd861,
    COMP_LOOP_C_664 = 10'd862,
    COMP_LOOP_C_665 = 10'd863,
    COMP_LOOP_C_666 = 10'd864,
    COMP_LOOP_C_667 = 10'd865,
    COMP_LOOP_C_668 = 10'd866,
    COMP_LOOP_C_669 = 10'd867,
    COMP_LOOP_C_670 = 10'd868,
    COMP_LOOP_C_671 = 10'd869,
    COMP_LOOP_C_672 = 10'd870,
    COMP_LOOP_C_673 = 10'd871,
    COMP_LOOP_C_674 = 10'd872,
    COMP_LOOP_C_675 = 10'd873,
    COMP_LOOP_C_676 = 10'd874,
    COMP_LOOP_C_677 = 10'd875,
    COMP_LOOP_C_678 = 10'd876,
    COMP_LOOP_C_679 = 10'd877,
    COMP_LOOP_C_680 = 10'd878,
    COMP_LOOP_C_681 = 10'd879,
    COMP_LOOP_C_682 = 10'd880,
    COMP_LOOP_C_683 = 10'd881,
    COMP_LOOP_C_684 = 10'd882,
    COMP_LOOP_C_685 = 10'd883,
    COMP_LOOP_C_686 = 10'd884,
    COMP_LOOP_C_687 = 10'd885,
    COMP_LOOP_C_688 = 10'd886,
    COMP_LOOP_C_689 = 10'd887,
    COMP_LOOP_C_690 = 10'd888,
    COMP_LOOP_C_691 = 10'd889,
    COMP_LOOP_16_modExp_dev_1_while_C_0 = 10'd890,
    COMP_LOOP_16_modExp_dev_1_while_C_1 = 10'd891,
    COMP_LOOP_16_modExp_dev_1_while_C_2 = 10'd892,
    COMP_LOOP_16_modExp_dev_1_while_C_3 = 10'd893,
    COMP_LOOP_16_modExp_dev_1_while_C_4 = 10'd894,
    COMP_LOOP_16_modExp_dev_1_while_C_5 = 10'd895,
    COMP_LOOP_16_modExp_dev_1_while_C_6 = 10'd896,
    COMP_LOOP_16_modExp_dev_1_while_C_7 = 10'd897,
    COMP_LOOP_16_modExp_dev_1_while_C_8 = 10'd898,
    COMP_LOOP_16_modExp_dev_1_while_C_9 = 10'd899,
    COMP_LOOP_16_modExp_dev_1_while_C_10 = 10'd900,
    COMP_LOOP_16_modExp_dev_1_while_C_11 = 10'd901,
    COMP_LOOP_C_692 = 10'd902,
    COMP_LOOP_C_693 = 10'd903,
    COMP_LOOP_C_694 = 10'd904,
    COMP_LOOP_C_695 = 10'd905,
    COMP_LOOP_C_696 = 10'd906,
    COMP_LOOP_C_697 = 10'd907,
    COMP_LOOP_C_698 = 10'd908,
    COMP_LOOP_C_699 = 10'd909,
    COMP_LOOP_C_700 = 10'd910,
    COMP_LOOP_C_701 = 10'd911,
    COMP_LOOP_C_702 = 10'd912,
    COMP_LOOP_C_703 = 10'd913,
    COMP_LOOP_C_704 = 10'd914,
    COMP_LOOP_C_705 = 10'd915,
    COMP_LOOP_C_706 = 10'd916,
    COMP_LOOP_C_707 = 10'd917,
    COMP_LOOP_C_708 = 10'd918,
    COMP_LOOP_C_709 = 10'd919,
    COMP_LOOP_C_710 = 10'd920,
    COMP_LOOP_C_711 = 10'd921,
    COMP_LOOP_C_712 = 10'd922,
    COMP_LOOP_C_713 = 10'd923,
    COMP_LOOP_C_714 = 10'd924,
    COMP_LOOP_C_715 = 10'd925,
    COMP_LOOP_C_716 = 10'd926,
    COMP_LOOP_C_717 = 10'd927,
    COMP_LOOP_C_718 = 10'd928,
    COMP_LOOP_C_719 = 10'd929,
    COMP_LOOP_C_720 = 10'd930,
    STAGE_VEC_LOOP_C_1 = 10'd931,
    STAGE_MAIN_LOOP_C_4 = 10'd932,
    main_C_1 = 10'd933;

  reg [9:0] state_var;
  reg [9:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : inPlaceNTT_DIF_core_core_fsm_1
    case (state_var)
      STAGE_MAIN_LOOP_C_0 : begin
        fsm_output = 10'b0000000001;
        state_var_NS = STAGE_MAIN_LOOP_C_1;
      end
      STAGE_MAIN_LOOP_C_1 : begin
        fsm_output = 10'b0000000010;
        state_var_NS = STAGE_MAIN_LOOP_C_2;
      end
      STAGE_MAIN_LOOP_C_2 : begin
        fsm_output = 10'b0000000011;
        state_var_NS = STAGE_MAIN_LOOP_C_3;
      end
      STAGE_MAIN_LOOP_C_3 : begin
        fsm_output = 10'b0000000100;
        if ( STAGE_MAIN_LOOP_C_3_tr0 ) begin
          state_var_NS = STAGE_VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = modExp_dev_while_C_0;
        end
      end
      modExp_dev_while_C_0 : begin
        fsm_output = 10'b0000000101;
        state_var_NS = modExp_dev_while_C_1;
      end
      modExp_dev_while_C_1 : begin
        fsm_output = 10'b0000000110;
        state_var_NS = modExp_dev_while_C_2;
      end
      modExp_dev_while_C_2 : begin
        fsm_output = 10'b0000000111;
        state_var_NS = modExp_dev_while_C_3;
      end
      modExp_dev_while_C_3 : begin
        fsm_output = 10'b0000001000;
        state_var_NS = modExp_dev_while_C_4;
      end
      modExp_dev_while_C_4 : begin
        fsm_output = 10'b0000001001;
        state_var_NS = modExp_dev_while_C_5;
      end
      modExp_dev_while_C_5 : begin
        fsm_output = 10'b0000001010;
        state_var_NS = modExp_dev_while_C_6;
      end
      modExp_dev_while_C_6 : begin
        fsm_output = 10'b0000001011;
        state_var_NS = modExp_dev_while_C_7;
      end
      modExp_dev_while_C_7 : begin
        fsm_output = 10'b0000001100;
        state_var_NS = modExp_dev_while_C_8;
      end
      modExp_dev_while_C_8 : begin
        fsm_output = 10'b0000001101;
        state_var_NS = modExp_dev_while_C_9;
      end
      modExp_dev_while_C_9 : begin
        fsm_output = 10'b0000001110;
        state_var_NS = modExp_dev_while_C_10;
      end
      modExp_dev_while_C_10 : begin
        fsm_output = 10'b0000001111;
        state_var_NS = modExp_dev_while_C_11;
      end
      modExp_dev_while_C_11 : begin
        fsm_output = 10'b0000010000;
        if ( modExp_dev_while_C_11_tr0 ) begin
          state_var_NS = STAGE_VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = modExp_dev_while_C_0;
        end
      end
      STAGE_VEC_LOOP_C_0 : begin
        fsm_output = 10'b0000010001;
        if ( STAGE_VEC_LOOP_C_0_tr0 ) begin
          state_var_NS = STAGE_VEC_LOOP_C_1;
        end
        else begin
          state_var_NS = COMP_LOOP_C_0;
        end
      end
      COMP_LOOP_C_0 : begin
        fsm_output = 10'b0000010010;
        state_var_NS = COMP_LOOP_C_1;
      end
      COMP_LOOP_C_1 : begin
        fsm_output = 10'b0000010011;
        state_var_NS = COMP_LOOP_C_2;
      end
      COMP_LOOP_C_2 : begin
        fsm_output = 10'b0000010100;
        state_var_NS = COMP_LOOP_C_3;
      end
      COMP_LOOP_C_3 : begin
        fsm_output = 10'b0000010101;
        state_var_NS = COMP_LOOP_C_4;
      end
      COMP_LOOP_C_4 : begin
        fsm_output = 10'b0000010110;
        state_var_NS = COMP_LOOP_C_5;
      end
      COMP_LOOP_C_5 : begin
        fsm_output = 10'b0000010111;
        state_var_NS = COMP_LOOP_C_6;
      end
      COMP_LOOP_C_6 : begin
        fsm_output = 10'b0000011000;
        state_var_NS = COMP_LOOP_C_7;
      end
      COMP_LOOP_C_7 : begin
        fsm_output = 10'b0000011001;
        state_var_NS = COMP_LOOP_C_8;
      end
      COMP_LOOP_C_8 : begin
        fsm_output = 10'b0000011010;
        state_var_NS = COMP_LOOP_C_9;
      end
      COMP_LOOP_C_9 : begin
        fsm_output = 10'b0000011011;
        state_var_NS = COMP_LOOP_C_10;
      end
      COMP_LOOP_C_10 : begin
        fsm_output = 10'b0000011100;
        state_var_NS = COMP_LOOP_C_11;
      end
      COMP_LOOP_C_11 : begin
        fsm_output = 10'b0000011101;
        state_var_NS = COMP_LOOP_C_12;
      end
      COMP_LOOP_C_12 : begin
        fsm_output = 10'b0000011110;
        state_var_NS = COMP_LOOP_C_13;
      end
      COMP_LOOP_C_13 : begin
        fsm_output = 10'b0000011111;
        state_var_NS = COMP_LOOP_C_14;
      end
      COMP_LOOP_C_14 : begin
        fsm_output = 10'b0000100000;
        state_var_NS = COMP_LOOP_C_15;
      end
      COMP_LOOP_C_15 : begin
        fsm_output = 10'b0000100001;
        state_var_NS = COMP_LOOP_C_16;
      end
      COMP_LOOP_C_16 : begin
        fsm_output = 10'b0000100010;
        if ( COMP_LOOP_C_16_tr0 ) begin
          state_var_NS = COMP_LOOP_C_17;
        end
        else begin
          state_var_NS = COMP_LOOP_1_modExp_dev_1_while_C_0;
        end
      end
      COMP_LOOP_1_modExp_dev_1_while_C_0 : begin
        fsm_output = 10'b0000100011;
        state_var_NS = COMP_LOOP_1_modExp_dev_1_while_C_1;
      end
      COMP_LOOP_1_modExp_dev_1_while_C_1 : begin
        fsm_output = 10'b0000100100;
        state_var_NS = COMP_LOOP_1_modExp_dev_1_while_C_2;
      end
      COMP_LOOP_1_modExp_dev_1_while_C_2 : begin
        fsm_output = 10'b0000100101;
        state_var_NS = COMP_LOOP_1_modExp_dev_1_while_C_3;
      end
      COMP_LOOP_1_modExp_dev_1_while_C_3 : begin
        fsm_output = 10'b0000100110;
        state_var_NS = COMP_LOOP_1_modExp_dev_1_while_C_4;
      end
      COMP_LOOP_1_modExp_dev_1_while_C_4 : begin
        fsm_output = 10'b0000100111;
        state_var_NS = COMP_LOOP_1_modExp_dev_1_while_C_5;
      end
      COMP_LOOP_1_modExp_dev_1_while_C_5 : begin
        fsm_output = 10'b0000101000;
        state_var_NS = COMP_LOOP_1_modExp_dev_1_while_C_6;
      end
      COMP_LOOP_1_modExp_dev_1_while_C_6 : begin
        fsm_output = 10'b0000101001;
        state_var_NS = COMP_LOOP_1_modExp_dev_1_while_C_7;
      end
      COMP_LOOP_1_modExp_dev_1_while_C_7 : begin
        fsm_output = 10'b0000101010;
        state_var_NS = COMP_LOOP_1_modExp_dev_1_while_C_8;
      end
      COMP_LOOP_1_modExp_dev_1_while_C_8 : begin
        fsm_output = 10'b0000101011;
        state_var_NS = COMP_LOOP_1_modExp_dev_1_while_C_9;
      end
      COMP_LOOP_1_modExp_dev_1_while_C_9 : begin
        fsm_output = 10'b0000101100;
        state_var_NS = COMP_LOOP_1_modExp_dev_1_while_C_10;
      end
      COMP_LOOP_1_modExp_dev_1_while_C_10 : begin
        fsm_output = 10'b0000101101;
        state_var_NS = COMP_LOOP_1_modExp_dev_1_while_C_11;
      end
      COMP_LOOP_1_modExp_dev_1_while_C_11 : begin
        fsm_output = 10'b0000101110;
        if ( COMP_LOOP_1_modExp_dev_1_while_C_11_tr0 ) begin
          state_var_NS = COMP_LOOP_C_17;
        end
        else begin
          state_var_NS = COMP_LOOP_1_modExp_dev_1_while_C_0;
        end
      end
      COMP_LOOP_C_17 : begin
        fsm_output = 10'b0000101111;
        state_var_NS = COMP_LOOP_C_18;
      end
      COMP_LOOP_C_18 : begin
        fsm_output = 10'b0000110000;
        state_var_NS = COMP_LOOP_C_19;
      end
      COMP_LOOP_C_19 : begin
        fsm_output = 10'b0000110001;
        state_var_NS = COMP_LOOP_C_20;
      end
      COMP_LOOP_C_20 : begin
        fsm_output = 10'b0000110010;
        state_var_NS = COMP_LOOP_C_21;
      end
      COMP_LOOP_C_21 : begin
        fsm_output = 10'b0000110011;
        state_var_NS = COMP_LOOP_C_22;
      end
      COMP_LOOP_C_22 : begin
        fsm_output = 10'b0000110100;
        state_var_NS = COMP_LOOP_C_23;
      end
      COMP_LOOP_C_23 : begin
        fsm_output = 10'b0000110101;
        state_var_NS = COMP_LOOP_C_24;
      end
      COMP_LOOP_C_24 : begin
        fsm_output = 10'b0000110110;
        state_var_NS = COMP_LOOP_C_25;
      end
      COMP_LOOP_C_25 : begin
        fsm_output = 10'b0000110111;
        state_var_NS = COMP_LOOP_C_26;
      end
      COMP_LOOP_C_26 : begin
        fsm_output = 10'b0000111000;
        state_var_NS = COMP_LOOP_C_27;
      end
      COMP_LOOP_C_27 : begin
        fsm_output = 10'b0000111001;
        state_var_NS = COMP_LOOP_C_28;
      end
      COMP_LOOP_C_28 : begin
        fsm_output = 10'b0000111010;
        state_var_NS = COMP_LOOP_C_29;
      end
      COMP_LOOP_C_29 : begin
        fsm_output = 10'b0000111011;
        state_var_NS = COMP_LOOP_C_30;
      end
      COMP_LOOP_C_30 : begin
        fsm_output = 10'b0000111100;
        state_var_NS = COMP_LOOP_C_31;
      end
      COMP_LOOP_C_31 : begin
        fsm_output = 10'b0000111101;
        state_var_NS = COMP_LOOP_C_32;
      end
      COMP_LOOP_C_32 : begin
        fsm_output = 10'b0000111110;
        state_var_NS = COMP_LOOP_C_33;
      end
      COMP_LOOP_C_33 : begin
        fsm_output = 10'b0000111111;
        state_var_NS = COMP_LOOP_C_34;
      end
      COMP_LOOP_C_34 : begin
        fsm_output = 10'b0001000000;
        state_var_NS = COMP_LOOP_C_35;
      end
      COMP_LOOP_C_35 : begin
        fsm_output = 10'b0001000001;
        state_var_NS = COMP_LOOP_C_36;
      end
      COMP_LOOP_C_36 : begin
        fsm_output = 10'b0001000010;
        state_var_NS = COMP_LOOP_C_37;
      end
      COMP_LOOP_C_37 : begin
        fsm_output = 10'b0001000011;
        state_var_NS = COMP_LOOP_C_38;
      end
      COMP_LOOP_C_38 : begin
        fsm_output = 10'b0001000100;
        state_var_NS = COMP_LOOP_C_39;
      end
      COMP_LOOP_C_39 : begin
        fsm_output = 10'b0001000101;
        state_var_NS = COMP_LOOP_C_40;
      end
      COMP_LOOP_C_40 : begin
        fsm_output = 10'b0001000110;
        state_var_NS = COMP_LOOP_C_41;
      end
      COMP_LOOP_C_41 : begin
        fsm_output = 10'b0001000111;
        state_var_NS = COMP_LOOP_C_42;
      end
      COMP_LOOP_C_42 : begin
        fsm_output = 10'b0001001000;
        state_var_NS = COMP_LOOP_C_43;
      end
      COMP_LOOP_C_43 : begin
        fsm_output = 10'b0001001001;
        state_var_NS = COMP_LOOP_C_44;
      end
      COMP_LOOP_C_44 : begin
        fsm_output = 10'b0001001010;
        state_var_NS = COMP_LOOP_C_45;
      end
      COMP_LOOP_C_45 : begin
        fsm_output = 10'b0001001011;
        if ( COMP_LOOP_C_45_tr0 ) begin
          state_var_NS = STAGE_VEC_LOOP_C_1;
        end
        else begin
          state_var_NS = COMP_LOOP_C_46;
        end
      end
      COMP_LOOP_C_46 : begin
        fsm_output = 10'b0001001100;
        state_var_NS = COMP_LOOP_C_47;
      end
      COMP_LOOP_C_47 : begin
        fsm_output = 10'b0001001101;
        state_var_NS = COMP_LOOP_C_48;
      end
      COMP_LOOP_C_48 : begin
        fsm_output = 10'b0001001110;
        state_var_NS = COMP_LOOP_C_49;
      end
      COMP_LOOP_C_49 : begin
        fsm_output = 10'b0001001111;
        state_var_NS = COMP_LOOP_C_50;
      end
      COMP_LOOP_C_50 : begin
        fsm_output = 10'b0001010000;
        state_var_NS = COMP_LOOP_C_51;
      end
      COMP_LOOP_C_51 : begin
        fsm_output = 10'b0001010001;
        state_var_NS = COMP_LOOP_C_52;
      end
      COMP_LOOP_C_52 : begin
        fsm_output = 10'b0001010010;
        state_var_NS = COMP_LOOP_C_53;
      end
      COMP_LOOP_C_53 : begin
        fsm_output = 10'b0001010011;
        state_var_NS = COMP_LOOP_C_54;
      end
      COMP_LOOP_C_54 : begin
        fsm_output = 10'b0001010100;
        state_var_NS = COMP_LOOP_C_55;
      end
      COMP_LOOP_C_55 : begin
        fsm_output = 10'b0001010101;
        state_var_NS = COMP_LOOP_C_56;
      end
      COMP_LOOP_C_56 : begin
        fsm_output = 10'b0001010110;
        state_var_NS = COMP_LOOP_C_57;
      end
      COMP_LOOP_C_57 : begin
        fsm_output = 10'b0001010111;
        state_var_NS = COMP_LOOP_C_58;
      end
      COMP_LOOP_C_58 : begin
        fsm_output = 10'b0001011000;
        state_var_NS = COMP_LOOP_C_59;
      end
      COMP_LOOP_C_59 : begin
        fsm_output = 10'b0001011001;
        state_var_NS = COMP_LOOP_C_60;
      end
      COMP_LOOP_C_60 : begin
        fsm_output = 10'b0001011010;
        state_var_NS = COMP_LOOP_C_61;
      end
      COMP_LOOP_C_61 : begin
        fsm_output = 10'b0001011011;
        state_var_NS = COMP_LOOP_2_modExp_dev_1_while_C_0;
      end
      COMP_LOOP_2_modExp_dev_1_while_C_0 : begin
        fsm_output = 10'b0001011100;
        state_var_NS = COMP_LOOP_2_modExp_dev_1_while_C_1;
      end
      COMP_LOOP_2_modExp_dev_1_while_C_1 : begin
        fsm_output = 10'b0001011101;
        state_var_NS = COMP_LOOP_2_modExp_dev_1_while_C_2;
      end
      COMP_LOOP_2_modExp_dev_1_while_C_2 : begin
        fsm_output = 10'b0001011110;
        state_var_NS = COMP_LOOP_2_modExp_dev_1_while_C_3;
      end
      COMP_LOOP_2_modExp_dev_1_while_C_3 : begin
        fsm_output = 10'b0001011111;
        state_var_NS = COMP_LOOP_2_modExp_dev_1_while_C_4;
      end
      COMP_LOOP_2_modExp_dev_1_while_C_4 : begin
        fsm_output = 10'b0001100000;
        state_var_NS = COMP_LOOP_2_modExp_dev_1_while_C_5;
      end
      COMP_LOOP_2_modExp_dev_1_while_C_5 : begin
        fsm_output = 10'b0001100001;
        state_var_NS = COMP_LOOP_2_modExp_dev_1_while_C_6;
      end
      COMP_LOOP_2_modExp_dev_1_while_C_6 : begin
        fsm_output = 10'b0001100010;
        state_var_NS = COMP_LOOP_2_modExp_dev_1_while_C_7;
      end
      COMP_LOOP_2_modExp_dev_1_while_C_7 : begin
        fsm_output = 10'b0001100011;
        state_var_NS = COMP_LOOP_2_modExp_dev_1_while_C_8;
      end
      COMP_LOOP_2_modExp_dev_1_while_C_8 : begin
        fsm_output = 10'b0001100100;
        state_var_NS = COMP_LOOP_2_modExp_dev_1_while_C_9;
      end
      COMP_LOOP_2_modExp_dev_1_while_C_9 : begin
        fsm_output = 10'b0001100101;
        state_var_NS = COMP_LOOP_2_modExp_dev_1_while_C_10;
      end
      COMP_LOOP_2_modExp_dev_1_while_C_10 : begin
        fsm_output = 10'b0001100110;
        state_var_NS = COMP_LOOP_2_modExp_dev_1_while_C_11;
      end
      COMP_LOOP_2_modExp_dev_1_while_C_11 : begin
        fsm_output = 10'b0001100111;
        if ( COMP_LOOP_2_modExp_dev_1_while_C_11_tr0 ) begin
          state_var_NS = COMP_LOOP_C_62;
        end
        else begin
          state_var_NS = COMP_LOOP_2_modExp_dev_1_while_C_0;
        end
      end
      COMP_LOOP_C_62 : begin
        fsm_output = 10'b0001101000;
        state_var_NS = COMP_LOOP_C_63;
      end
      COMP_LOOP_C_63 : begin
        fsm_output = 10'b0001101001;
        state_var_NS = COMP_LOOP_C_64;
      end
      COMP_LOOP_C_64 : begin
        fsm_output = 10'b0001101010;
        state_var_NS = COMP_LOOP_C_65;
      end
      COMP_LOOP_C_65 : begin
        fsm_output = 10'b0001101011;
        state_var_NS = COMP_LOOP_C_66;
      end
      COMP_LOOP_C_66 : begin
        fsm_output = 10'b0001101100;
        state_var_NS = COMP_LOOP_C_67;
      end
      COMP_LOOP_C_67 : begin
        fsm_output = 10'b0001101101;
        state_var_NS = COMP_LOOP_C_68;
      end
      COMP_LOOP_C_68 : begin
        fsm_output = 10'b0001101110;
        state_var_NS = COMP_LOOP_C_69;
      end
      COMP_LOOP_C_69 : begin
        fsm_output = 10'b0001101111;
        state_var_NS = COMP_LOOP_C_70;
      end
      COMP_LOOP_C_70 : begin
        fsm_output = 10'b0001110000;
        state_var_NS = COMP_LOOP_C_71;
      end
      COMP_LOOP_C_71 : begin
        fsm_output = 10'b0001110001;
        state_var_NS = COMP_LOOP_C_72;
      end
      COMP_LOOP_C_72 : begin
        fsm_output = 10'b0001110010;
        state_var_NS = COMP_LOOP_C_73;
      end
      COMP_LOOP_C_73 : begin
        fsm_output = 10'b0001110011;
        state_var_NS = COMP_LOOP_C_74;
      end
      COMP_LOOP_C_74 : begin
        fsm_output = 10'b0001110100;
        state_var_NS = COMP_LOOP_C_75;
      end
      COMP_LOOP_C_75 : begin
        fsm_output = 10'b0001110101;
        state_var_NS = COMP_LOOP_C_76;
      end
      COMP_LOOP_C_76 : begin
        fsm_output = 10'b0001110110;
        state_var_NS = COMP_LOOP_C_77;
      end
      COMP_LOOP_C_77 : begin
        fsm_output = 10'b0001110111;
        state_var_NS = COMP_LOOP_C_78;
      end
      COMP_LOOP_C_78 : begin
        fsm_output = 10'b0001111000;
        state_var_NS = COMP_LOOP_C_79;
      end
      COMP_LOOP_C_79 : begin
        fsm_output = 10'b0001111001;
        state_var_NS = COMP_LOOP_C_80;
      end
      COMP_LOOP_C_80 : begin
        fsm_output = 10'b0001111010;
        state_var_NS = COMP_LOOP_C_81;
      end
      COMP_LOOP_C_81 : begin
        fsm_output = 10'b0001111011;
        state_var_NS = COMP_LOOP_C_82;
      end
      COMP_LOOP_C_82 : begin
        fsm_output = 10'b0001111100;
        state_var_NS = COMP_LOOP_C_83;
      end
      COMP_LOOP_C_83 : begin
        fsm_output = 10'b0001111101;
        state_var_NS = COMP_LOOP_C_84;
      end
      COMP_LOOP_C_84 : begin
        fsm_output = 10'b0001111110;
        state_var_NS = COMP_LOOP_C_85;
      end
      COMP_LOOP_C_85 : begin
        fsm_output = 10'b0001111111;
        state_var_NS = COMP_LOOP_C_86;
      end
      COMP_LOOP_C_86 : begin
        fsm_output = 10'b0010000000;
        state_var_NS = COMP_LOOP_C_87;
      end
      COMP_LOOP_C_87 : begin
        fsm_output = 10'b0010000001;
        state_var_NS = COMP_LOOP_C_88;
      end
      COMP_LOOP_C_88 : begin
        fsm_output = 10'b0010000010;
        state_var_NS = COMP_LOOP_C_89;
      end
      COMP_LOOP_C_89 : begin
        fsm_output = 10'b0010000011;
        state_var_NS = COMP_LOOP_C_90;
      end
      COMP_LOOP_C_90 : begin
        fsm_output = 10'b0010000100;
        if ( COMP_LOOP_C_90_tr0 ) begin
          state_var_NS = STAGE_VEC_LOOP_C_1;
        end
        else begin
          state_var_NS = COMP_LOOP_C_91;
        end
      end
      COMP_LOOP_C_91 : begin
        fsm_output = 10'b0010000101;
        state_var_NS = COMP_LOOP_C_92;
      end
      COMP_LOOP_C_92 : begin
        fsm_output = 10'b0010000110;
        state_var_NS = COMP_LOOP_C_93;
      end
      COMP_LOOP_C_93 : begin
        fsm_output = 10'b0010000111;
        state_var_NS = COMP_LOOP_C_94;
      end
      COMP_LOOP_C_94 : begin
        fsm_output = 10'b0010001000;
        state_var_NS = COMP_LOOP_C_95;
      end
      COMP_LOOP_C_95 : begin
        fsm_output = 10'b0010001001;
        state_var_NS = COMP_LOOP_C_96;
      end
      COMP_LOOP_C_96 : begin
        fsm_output = 10'b0010001010;
        state_var_NS = COMP_LOOP_C_97;
      end
      COMP_LOOP_C_97 : begin
        fsm_output = 10'b0010001011;
        state_var_NS = COMP_LOOP_C_98;
      end
      COMP_LOOP_C_98 : begin
        fsm_output = 10'b0010001100;
        state_var_NS = COMP_LOOP_C_99;
      end
      COMP_LOOP_C_99 : begin
        fsm_output = 10'b0010001101;
        state_var_NS = COMP_LOOP_C_100;
      end
      COMP_LOOP_C_100 : begin
        fsm_output = 10'b0010001110;
        state_var_NS = COMP_LOOP_C_101;
      end
      COMP_LOOP_C_101 : begin
        fsm_output = 10'b0010001111;
        state_var_NS = COMP_LOOP_C_102;
      end
      COMP_LOOP_C_102 : begin
        fsm_output = 10'b0010010000;
        state_var_NS = COMP_LOOP_C_103;
      end
      COMP_LOOP_C_103 : begin
        fsm_output = 10'b0010010001;
        state_var_NS = COMP_LOOP_C_104;
      end
      COMP_LOOP_C_104 : begin
        fsm_output = 10'b0010010010;
        state_var_NS = COMP_LOOP_C_105;
      end
      COMP_LOOP_C_105 : begin
        fsm_output = 10'b0010010011;
        state_var_NS = COMP_LOOP_C_106;
      end
      COMP_LOOP_C_106 : begin
        fsm_output = 10'b0010010100;
        state_var_NS = COMP_LOOP_3_modExp_dev_1_while_C_0;
      end
      COMP_LOOP_3_modExp_dev_1_while_C_0 : begin
        fsm_output = 10'b0010010101;
        state_var_NS = COMP_LOOP_3_modExp_dev_1_while_C_1;
      end
      COMP_LOOP_3_modExp_dev_1_while_C_1 : begin
        fsm_output = 10'b0010010110;
        state_var_NS = COMP_LOOP_3_modExp_dev_1_while_C_2;
      end
      COMP_LOOP_3_modExp_dev_1_while_C_2 : begin
        fsm_output = 10'b0010010111;
        state_var_NS = COMP_LOOP_3_modExp_dev_1_while_C_3;
      end
      COMP_LOOP_3_modExp_dev_1_while_C_3 : begin
        fsm_output = 10'b0010011000;
        state_var_NS = COMP_LOOP_3_modExp_dev_1_while_C_4;
      end
      COMP_LOOP_3_modExp_dev_1_while_C_4 : begin
        fsm_output = 10'b0010011001;
        state_var_NS = COMP_LOOP_3_modExp_dev_1_while_C_5;
      end
      COMP_LOOP_3_modExp_dev_1_while_C_5 : begin
        fsm_output = 10'b0010011010;
        state_var_NS = COMP_LOOP_3_modExp_dev_1_while_C_6;
      end
      COMP_LOOP_3_modExp_dev_1_while_C_6 : begin
        fsm_output = 10'b0010011011;
        state_var_NS = COMP_LOOP_3_modExp_dev_1_while_C_7;
      end
      COMP_LOOP_3_modExp_dev_1_while_C_7 : begin
        fsm_output = 10'b0010011100;
        state_var_NS = COMP_LOOP_3_modExp_dev_1_while_C_8;
      end
      COMP_LOOP_3_modExp_dev_1_while_C_8 : begin
        fsm_output = 10'b0010011101;
        state_var_NS = COMP_LOOP_3_modExp_dev_1_while_C_9;
      end
      COMP_LOOP_3_modExp_dev_1_while_C_9 : begin
        fsm_output = 10'b0010011110;
        state_var_NS = COMP_LOOP_3_modExp_dev_1_while_C_10;
      end
      COMP_LOOP_3_modExp_dev_1_while_C_10 : begin
        fsm_output = 10'b0010011111;
        state_var_NS = COMP_LOOP_3_modExp_dev_1_while_C_11;
      end
      COMP_LOOP_3_modExp_dev_1_while_C_11 : begin
        fsm_output = 10'b0010100000;
        if ( COMP_LOOP_3_modExp_dev_1_while_C_11_tr0 ) begin
          state_var_NS = COMP_LOOP_C_107;
        end
        else begin
          state_var_NS = COMP_LOOP_3_modExp_dev_1_while_C_0;
        end
      end
      COMP_LOOP_C_107 : begin
        fsm_output = 10'b0010100001;
        state_var_NS = COMP_LOOP_C_108;
      end
      COMP_LOOP_C_108 : begin
        fsm_output = 10'b0010100010;
        state_var_NS = COMP_LOOP_C_109;
      end
      COMP_LOOP_C_109 : begin
        fsm_output = 10'b0010100011;
        state_var_NS = COMP_LOOP_C_110;
      end
      COMP_LOOP_C_110 : begin
        fsm_output = 10'b0010100100;
        state_var_NS = COMP_LOOP_C_111;
      end
      COMP_LOOP_C_111 : begin
        fsm_output = 10'b0010100101;
        state_var_NS = COMP_LOOP_C_112;
      end
      COMP_LOOP_C_112 : begin
        fsm_output = 10'b0010100110;
        state_var_NS = COMP_LOOP_C_113;
      end
      COMP_LOOP_C_113 : begin
        fsm_output = 10'b0010100111;
        state_var_NS = COMP_LOOP_C_114;
      end
      COMP_LOOP_C_114 : begin
        fsm_output = 10'b0010101000;
        state_var_NS = COMP_LOOP_C_115;
      end
      COMP_LOOP_C_115 : begin
        fsm_output = 10'b0010101001;
        state_var_NS = COMP_LOOP_C_116;
      end
      COMP_LOOP_C_116 : begin
        fsm_output = 10'b0010101010;
        state_var_NS = COMP_LOOP_C_117;
      end
      COMP_LOOP_C_117 : begin
        fsm_output = 10'b0010101011;
        state_var_NS = COMP_LOOP_C_118;
      end
      COMP_LOOP_C_118 : begin
        fsm_output = 10'b0010101100;
        state_var_NS = COMP_LOOP_C_119;
      end
      COMP_LOOP_C_119 : begin
        fsm_output = 10'b0010101101;
        state_var_NS = COMP_LOOP_C_120;
      end
      COMP_LOOP_C_120 : begin
        fsm_output = 10'b0010101110;
        state_var_NS = COMP_LOOP_C_121;
      end
      COMP_LOOP_C_121 : begin
        fsm_output = 10'b0010101111;
        state_var_NS = COMP_LOOP_C_122;
      end
      COMP_LOOP_C_122 : begin
        fsm_output = 10'b0010110000;
        state_var_NS = COMP_LOOP_C_123;
      end
      COMP_LOOP_C_123 : begin
        fsm_output = 10'b0010110001;
        state_var_NS = COMP_LOOP_C_124;
      end
      COMP_LOOP_C_124 : begin
        fsm_output = 10'b0010110010;
        state_var_NS = COMP_LOOP_C_125;
      end
      COMP_LOOP_C_125 : begin
        fsm_output = 10'b0010110011;
        state_var_NS = COMP_LOOP_C_126;
      end
      COMP_LOOP_C_126 : begin
        fsm_output = 10'b0010110100;
        state_var_NS = COMP_LOOP_C_127;
      end
      COMP_LOOP_C_127 : begin
        fsm_output = 10'b0010110101;
        state_var_NS = COMP_LOOP_C_128;
      end
      COMP_LOOP_C_128 : begin
        fsm_output = 10'b0010110110;
        state_var_NS = COMP_LOOP_C_129;
      end
      COMP_LOOP_C_129 : begin
        fsm_output = 10'b0010110111;
        state_var_NS = COMP_LOOP_C_130;
      end
      COMP_LOOP_C_130 : begin
        fsm_output = 10'b0010111000;
        state_var_NS = COMP_LOOP_C_131;
      end
      COMP_LOOP_C_131 : begin
        fsm_output = 10'b0010111001;
        state_var_NS = COMP_LOOP_C_132;
      end
      COMP_LOOP_C_132 : begin
        fsm_output = 10'b0010111010;
        state_var_NS = COMP_LOOP_C_133;
      end
      COMP_LOOP_C_133 : begin
        fsm_output = 10'b0010111011;
        state_var_NS = COMP_LOOP_C_134;
      end
      COMP_LOOP_C_134 : begin
        fsm_output = 10'b0010111100;
        state_var_NS = COMP_LOOP_C_135;
      end
      COMP_LOOP_C_135 : begin
        fsm_output = 10'b0010111101;
        if ( COMP_LOOP_C_135_tr0 ) begin
          state_var_NS = STAGE_VEC_LOOP_C_1;
        end
        else begin
          state_var_NS = COMP_LOOP_C_136;
        end
      end
      COMP_LOOP_C_136 : begin
        fsm_output = 10'b0010111110;
        state_var_NS = COMP_LOOP_C_137;
      end
      COMP_LOOP_C_137 : begin
        fsm_output = 10'b0010111111;
        state_var_NS = COMP_LOOP_C_138;
      end
      COMP_LOOP_C_138 : begin
        fsm_output = 10'b0011000000;
        state_var_NS = COMP_LOOP_C_139;
      end
      COMP_LOOP_C_139 : begin
        fsm_output = 10'b0011000001;
        state_var_NS = COMP_LOOP_C_140;
      end
      COMP_LOOP_C_140 : begin
        fsm_output = 10'b0011000010;
        state_var_NS = COMP_LOOP_C_141;
      end
      COMP_LOOP_C_141 : begin
        fsm_output = 10'b0011000011;
        state_var_NS = COMP_LOOP_C_142;
      end
      COMP_LOOP_C_142 : begin
        fsm_output = 10'b0011000100;
        state_var_NS = COMP_LOOP_C_143;
      end
      COMP_LOOP_C_143 : begin
        fsm_output = 10'b0011000101;
        state_var_NS = COMP_LOOP_C_144;
      end
      COMP_LOOP_C_144 : begin
        fsm_output = 10'b0011000110;
        state_var_NS = COMP_LOOP_C_145;
      end
      COMP_LOOP_C_145 : begin
        fsm_output = 10'b0011000111;
        state_var_NS = COMP_LOOP_C_146;
      end
      COMP_LOOP_C_146 : begin
        fsm_output = 10'b0011001000;
        state_var_NS = COMP_LOOP_C_147;
      end
      COMP_LOOP_C_147 : begin
        fsm_output = 10'b0011001001;
        state_var_NS = COMP_LOOP_C_148;
      end
      COMP_LOOP_C_148 : begin
        fsm_output = 10'b0011001010;
        state_var_NS = COMP_LOOP_C_149;
      end
      COMP_LOOP_C_149 : begin
        fsm_output = 10'b0011001011;
        state_var_NS = COMP_LOOP_C_150;
      end
      COMP_LOOP_C_150 : begin
        fsm_output = 10'b0011001100;
        state_var_NS = COMP_LOOP_C_151;
      end
      COMP_LOOP_C_151 : begin
        fsm_output = 10'b0011001101;
        state_var_NS = COMP_LOOP_4_modExp_dev_1_while_C_0;
      end
      COMP_LOOP_4_modExp_dev_1_while_C_0 : begin
        fsm_output = 10'b0011001110;
        state_var_NS = COMP_LOOP_4_modExp_dev_1_while_C_1;
      end
      COMP_LOOP_4_modExp_dev_1_while_C_1 : begin
        fsm_output = 10'b0011001111;
        state_var_NS = COMP_LOOP_4_modExp_dev_1_while_C_2;
      end
      COMP_LOOP_4_modExp_dev_1_while_C_2 : begin
        fsm_output = 10'b0011010000;
        state_var_NS = COMP_LOOP_4_modExp_dev_1_while_C_3;
      end
      COMP_LOOP_4_modExp_dev_1_while_C_3 : begin
        fsm_output = 10'b0011010001;
        state_var_NS = COMP_LOOP_4_modExp_dev_1_while_C_4;
      end
      COMP_LOOP_4_modExp_dev_1_while_C_4 : begin
        fsm_output = 10'b0011010010;
        state_var_NS = COMP_LOOP_4_modExp_dev_1_while_C_5;
      end
      COMP_LOOP_4_modExp_dev_1_while_C_5 : begin
        fsm_output = 10'b0011010011;
        state_var_NS = COMP_LOOP_4_modExp_dev_1_while_C_6;
      end
      COMP_LOOP_4_modExp_dev_1_while_C_6 : begin
        fsm_output = 10'b0011010100;
        state_var_NS = COMP_LOOP_4_modExp_dev_1_while_C_7;
      end
      COMP_LOOP_4_modExp_dev_1_while_C_7 : begin
        fsm_output = 10'b0011010101;
        state_var_NS = COMP_LOOP_4_modExp_dev_1_while_C_8;
      end
      COMP_LOOP_4_modExp_dev_1_while_C_8 : begin
        fsm_output = 10'b0011010110;
        state_var_NS = COMP_LOOP_4_modExp_dev_1_while_C_9;
      end
      COMP_LOOP_4_modExp_dev_1_while_C_9 : begin
        fsm_output = 10'b0011010111;
        state_var_NS = COMP_LOOP_4_modExp_dev_1_while_C_10;
      end
      COMP_LOOP_4_modExp_dev_1_while_C_10 : begin
        fsm_output = 10'b0011011000;
        state_var_NS = COMP_LOOP_4_modExp_dev_1_while_C_11;
      end
      COMP_LOOP_4_modExp_dev_1_while_C_11 : begin
        fsm_output = 10'b0011011001;
        if ( COMP_LOOP_4_modExp_dev_1_while_C_11_tr0 ) begin
          state_var_NS = COMP_LOOP_C_152;
        end
        else begin
          state_var_NS = COMP_LOOP_4_modExp_dev_1_while_C_0;
        end
      end
      COMP_LOOP_C_152 : begin
        fsm_output = 10'b0011011010;
        state_var_NS = COMP_LOOP_C_153;
      end
      COMP_LOOP_C_153 : begin
        fsm_output = 10'b0011011011;
        state_var_NS = COMP_LOOP_C_154;
      end
      COMP_LOOP_C_154 : begin
        fsm_output = 10'b0011011100;
        state_var_NS = COMP_LOOP_C_155;
      end
      COMP_LOOP_C_155 : begin
        fsm_output = 10'b0011011101;
        state_var_NS = COMP_LOOP_C_156;
      end
      COMP_LOOP_C_156 : begin
        fsm_output = 10'b0011011110;
        state_var_NS = COMP_LOOP_C_157;
      end
      COMP_LOOP_C_157 : begin
        fsm_output = 10'b0011011111;
        state_var_NS = COMP_LOOP_C_158;
      end
      COMP_LOOP_C_158 : begin
        fsm_output = 10'b0011100000;
        state_var_NS = COMP_LOOP_C_159;
      end
      COMP_LOOP_C_159 : begin
        fsm_output = 10'b0011100001;
        state_var_NS = COMP_LOOP_C_160;
      end
      COMP_LOOP_C_160 : begin
        fsm_output = 10'b0011100010;
        state_var_NS = COMP_LOOP_C_161;
      end
      COMP_LOOP_C_161 : begin
        fsm_output = 10'b0011100011;
        state_var_NS = COMP_LOOP_C_162;
      end
      COMP_LOOP_C_162 : begin
        fsm_output = 10'b0011100100;
        state_var_NS = COMP_LOOP_C_163;
      end
      COMP_LOOP_C_163 : begin
        fsm_output = 10'b0011100101;
        state_var_NS = COMP_LOOP_C_164;
      end
      COMP_LOOP_C_164 : begin
        fsm_output = 10'b0011100110;
        state_var_NS = COMP_LOOP_C_165;
      end
      COMP_LOOP_C_165 : begin
        fsm_output = 10'b0011100111;
        state_var_NS = COMP_LOOP_C_166;
      end
      COMP_LOOP_C_166 : begin
        fsm_output = 10'b0011101000;
        state_var_NS = COMP_LOOP_C_167;
      end
      COMP_LOOP_C_167 : begin
        fsm_output = 10'b0011101001;
        state_var_NS = COMP_LOOP_C_168;
      end
      COMP_LOOP_C_168 : begin
        fsm_output = 10'b0011101010;
        state_var_NS = COMP_LOOP_C_169;
      end
      COMP_LOOP_C_169 : begin
        fsm_output = 10'b0011101011;
        state_var_NS = COMP_LOOP_C_170;
      end
      COMP_LOOP_C_170 : begin
        fsm_output = 10'b0011101100;
        state_var_NS = COMP_LOOP_C_171;
      end
      COMP_LOOP_C_171 : begin
        fsm_output = 10'b0011101101;
        state_var_NS = COMP_LOOP_C_172;
      end
      COMP_LOOP_C_172 : begin
        fsm_output = 10'b0011101110;
        state_var_NS = COMP_LOOP_C_173;
      end
      COMP_LOOP_C_173 : begin
        fsm_output = 10'b0011101111;
        state_var_NS = COMP_LOOP_C_174;
      end
      COMP_LOOP_C_174 : begin
        fsm_output = 10'b0011110000;
        state_var_NS = COMP_LOOP_C_175;
      end
      COMP_LOOP_C_175 : begin
        fsm_output = 10'b0011110001;
        state_var_NS = COMP_LOOP_C_176;
      end
      COMP_LOOP_C_176 : begin
        fsm_output = 10'b0011110010;
        state_var_NS = COMP_LOOP_C_177;
      end
      COMP_LOOP_C_177 : begin
        fsm_output = 10'b0011110011;
        state_var_NS = COMP_LOOP_C_178;
      end
      COMP_LOOP_C_178 : begin
        fsm_output = 10'b0011110100;
        state_var_NS = COMP_LOOP_C_179;
      end
      COMP_LOOP_C_179 : begin
        fsm_output = 10'b0011110101;
        state_var_NS = COMP_LOOP_C_180;
      end
      COMP_LOOP_C_180 : begin
        fsm_output = 10'b0011110110;
        if ( COMP_LOOP_C_180_tr0 ) begin
          state_var_NS = STAGE_VEC_LOOP_C_1;
        end
        else begin
          state_var_NS = COMP_LOOP_C_181;
        end
      end
      COMP_LOOP_C_181 : begin
        fsm_output = 10'b0011110111;
        state_var_NS = COMP_LOOP_C_182;
      end
      COMP_LOOP_C_182 : begin
        fsm_output = 10'b0011111000;
        state_var_NS = COMP_LOOP_C_183;
      end
      COMP_LOOP_C_183 : begin
        fsm_output = 10'b0011111001;
        state_var_NS = COMP_LOOP_C_184;
      end
      COMP_LOOP_C_184 : begin
        fsm_output = 10'b0011111010;
        state_var_NS = COMP_LOOP_C_185;
      end
      COMP_LOOP_C_185 : begin
        fsm_output = 10'b0011111011;
        state_var_NS = COMP_LOOP_C_186;
      end
      COMP_LOOP_C_186 : begin
        fsm_output = 10'b0011111100;
        state_var_NS = COMP_LOOP_C_187;
      end
      COMP_LOOP_C_187 : begin
        fsm_output = 10'b0011111101;
        state_var_NS = COMP_LOOP_C_188;
      end
      COMP_LOOP_C_188 : begin
        fsm_output = 10'b0011111110;
        state_var_NS = COMP_LOOP_C_189;
      end
      COMP_LOOP_C_189 : begin
        fsm_output = 10'b0011111111;
        state_var_NS = COMP_LOOP_C_190;
      end
      COMP_LOOP_C_190 : begin
        fsm_output = 10'b0100000000;
        state_var_NS = COMP_LOOP_C_191;
      end
      COMP_LOOP_C_191 : begin
        fsm_output = 10'b0100000001;
        state_var_NS = COMP_LOOP_C_192;
      end
      COMP_LOOP_C_192 : begin
        fsm_output = 10'b0100000010;
        state_var_NS = COMP_LOOP_C_193;
      end
      COMP_LOOP_C_193 : begin
        fsm_output = 10'b0100000011;
        state_var_NS = COMP_LOOP_C_194;
      end
      COMP_LOOP_C_194 : begin
        fsm_output = 10'b0100000100;
        state_var_NS = COMP_LOOP_C_195;
      end
      COMP_LOOP_C_195 : begin
        fsm_output = 10'b0100000101;
        state_var_NS = COMP_LOOP_C_196;
      end
      COMP_LOOP_C_196 : begin
        fsm_output = 10'b0100000110;
        state_var_NS = COMP_LOOP_5_modExp_dev_1_while_C_0;
      end
      COMP_LOOP_5_modExp_dev_1_while_C_0 : begin
        fsm_output = 10'b0100000111;
        state_var_NS = COMP_LOOP_5_modExp_dev_1_while_C_1;
      end
      COMP_LOOP_5_modExp_dev_1_while_C_1 : begin
        fsm_output = 10'b0100001000;
        state_var_NS = COMP_LOOP_5_modExp_dev_1_while_C_2;
      end
      COMP_LOOP_5_modExp_dev_1_while_C_2 : begin
        fsm_output = 10'b0100001001;
        state_var_NS = COMP_LOOP_5_modExp_dev_1_while_C_3;
      end
      COMP_LOOP_5_modExp_dev_1_while_C_3 : begin
        fsm_output = 10'b0100001010;
        state_var_NS = COMP_LOOP_5_modExp_dev_1_while_C_4;
      end
      COMP_LOOP_5_modExp_dev_1_while_C_4 : begin
        fsm_output = 10'b0100001011;
        state_var_NS = COMP_LOOP_5_modExp_dev_1_while_C_5;
      end
      COMP_LOOP_5_modExp_dev_1_while_C_5 : begin
        fsm_output = 10'b0100001100;
        state_var_NS = COMP_LOOP_5_modExp_dev_1_while_C_6;
      end
      COMP_LOOP_5_modExp_dev_1_while_C_6 : begin
        fsm_output = 10'b0100001101;
        state_var_NS = COMP_LOOP_5_modExp_dev_1_while_C_7;
      end
      COMP_LOOP_5_modExp_dev_1_while_C_7 : begin
        fsm_output = 10'b0100001110;
        state_var_NS = COMP_LOOP_5_modExp_dev_1_while_C_8;
      end
      COMP_LOOP_5_modExp_dev_1_while_C_8 : begin
        fsm_output = 10'b0100001111;
        state_var_NS = COMP_LOOP_5_modExp_dev_1_while_C_9;
      end
      COMP_LOOP_5_modExp_dev_1_while_C_9 : begin
        fsm_output = 10'b0100010000;
        state_var_NS = COMP_LOOP_5_modExp_dev_1_while_C_10;
      end
      COMP_LOOP_5_modExp_dev_1_while_C_10 : begin
        fsm_output = 10'b0100010001;
        state_var_NS = COMP_LOOP_5_modExp_dev_1_while_C_11;
      end
      COMP_LOOP_5_modExp_dev_1_while_C_11 : begin
        fsm_output = 10'b0100010010;
        if ( COMP_LOOP_5_modExp_dev_1_while_C_11_tr0 ) begin
          state_var_NS = COMP_LOOP_C_197;
        end
        else begin
          state_var_NS = COMP_LOOP_5_modExp_dev_1_while_C_0;
        end
      end
      COMP_LOOP_C_197 : begin
        fsm_output = 10'b0100010011;
        state_var_NS = COMP_LOOP_C_198;
      end
      COMP_LOOP_C_198 : begin
        fsm_output = 10'b0100010100;
        state_var_NS = COMP_LOOP_C_199;
      end
      COMP_LOOP_C_199 : begin
        fsm_output = 10'b0100010101;
        state_var_NS = COMP_LOOP_C_200;
      end
      COMP_LOOP_C_200 : begin
        fsm_output = 10'b0100010110;
        state_var_NS = COMP_LOOP_C_201;
      end
      COMP_LOOP_C_201 : begin
        fsm_output = 10'b0100010111;
        state_var_NS = COMP_LOOP_C_202;
      end
      COMP_LOOP_C_202 : begin
        fsm_output = 10'b0100011000;
        state_var_NS = COMP_LOOP_C_203;
      end
      COMP_LOOP_C_203 : begin
        fsm_output = 10'b0100011001;
        state_var_NS = COMP_LOOP_C_204;
      end
      COMP_LOOP_C_204 : begin
        fsm_output = 10'b0100011010;
        state_var_NS = COMP_LOOP_C_205;
      end
      COMP_LOOP_C_205 : begin
        fsm_output = 10'b0100011011;
        state_var_NS = COMP_LOOP_C_206;
      end
      COMP_LOOP_C_206 : begin
        fsm_output = 10'b0100011100;
        state_var_NS = COMP_LOOP_C_207;
      end
      COMP_LOOP_C_207 : begin
        fsm_output = 10'b0100011101;
        state_var_NS = COMP_LOOP_C_208;
      end
      COMP_LOOP_C_208 : begin
        fsm_output = 10'b0100011110;
        state_var_NS = COMP_LOOP_C_209;
      end
      COMP_LOOP_C_209 : begin
        fsm_output = 10'b0100011111;
        state_var_NS = COMP_LOOP_C_210;
      end
      COMP_LOOP_C_210 : begin
        fsm_output = 10'b0100100000;
        state_var_NS = COMP_LOOP_C_211;
      end
      COMP_LOOP_C_211 : begin
        fsm_output = 10'b0100100001;
        state_var_NS = COMP_LOOP_C_212;
      end
      COMP_LOOP_C_212 : begin
        fsm_output = 10'b0100100010;
        state_var_NS = COMP_LOOP_C_213;
      end
      COMP_LOOP_C_213 : begin
        fsm_output = 10'b0100100011;
        state_var_NS = COMP_LOOP_C_214;
      end
      COMP_LOOP_C_214 : begin
        fsm_output = 10'b0100100100;
        state_var_NS = COMP_LOOP_C_215;
      end
      COMP_LOOP_C_215 : begin
        fsm_output = 10'b0100100101;
        state_var_NS = COMP_LOOP_C_216;
      end
      COMP_LOOP_C_216 : begin
        fsm_output = 10'b0100100110;
        state_var_NS = COMP_LOOP_C_217;
      end
      COMP_LOOP_C_217 : begin
        fsm_output = 10'b0100100111;
        state_var_NS = COMP_LOOP_C_218;
      end
      COMP_LOOP_C_218 : begin
        fsm_output = 10'b0100101000;
        state_var_NS = COMP_LOOP_C_219;
      end
      COMP_LOOP_C_219 : begin
        fsm_output = 10'b0100101001;
        state_var_NS = COMP_LOOP_C_220;
      end
      COMP_LOOP_C_220 : begin
        fsm_output = 10'b0100101010;
        state_var_NS = COMP_LOOP_C_221;
      end
      COMP_LOOP_C_221 : begin
        fsm_output = 10'b0100101011;
        state_var_NS = COMP_LOOP_C_222;
      end
      COMP_LOOP_C_222 : begin
        fsm_output = 10'b0100101100;
        state_var_NS = COMP_LOOP_C_223;
      end
      COMP_LOOP_C_223 : begin
        fsm_output = 10'b0100101101;
        state_var_NS = COMP_LOOP_C_224;
      end
      COMP_LOOP_C_224 : begin
        fsm_output = 10'b0100101110;
        state_var_NS = COMP_LOOP_C_225;
      end
      COMP_LOOP_C_225 : begin
        fsm_output = 10'b0100101111;
        if ( COMP_LOOP_C_225_tr0 ) begin
          state_var_NS = STAGE_VEC_LOOP_C_1;
        end
        else begin
          state_var_NS = COMP_LOOP_C_226;
        end
      end
      COMP_LOOP_C_226 : begin
        fsm_output = 10'b0100110000;
        state_var_NS = COMP_LOOP_C_227;
      end
      COMP_LOOP_C_227 : begin
        fsm_output = 10'b0100110001;
        state_var_NS = COMP_LOOP_C_228;
      end
      COMP_LOOP_C_228 : begin
        fsm_output = 10'b0100110010;
        state_var_NS = COMP_LOOP_C_229;
      end
      COMP_LOOP_C_229 : begin
        fsm_output = 10'b0100110011;
        state_var_NS = COMP_LOOP_C_230;
      end
      COMP_LOOP_C_230 : begin
        fsm_output = 10'b0100110100;
        state_var_NS = COMP_LOOP_C_231;
      end
      COMP_LOOP_C_231 : begin
        fsm_output = 10'b0100110101;
        state_var_NS = COMP_LOOP_C_232;
      end
      COMP_LOOP_C_232 : begin
        fsm_output = 10'b0100110110;
        state_var_NS = COMP_LOOP_C_233;
      end
      COMP_LOOP_C_233 : begin
        fsm_output = 10'b0100110111;
        state_var_NS = COMP_LOOP_C_234;
      end
      COMP_LOOP_C_234 : begin
        fsm_output = 10'b0100111000;
        state_var_NS = COMP_LOOP_C_235;
      end
      COMP_LOOP_C_235 : begin
        fsm_output = 10'b0100111001;
        state_var_NS = COMP_LOOP_C_236;
      end
      COMP_LOOP_C_236 : begin
        fsm_output = 10'b0100111010;
        state_var_NS = COMP_LOOP_C_237;
      end
      COMP_LOOP_C_237 : begin
        fsm_output = 10'b0100111011;
        state_var_NS = COMP_LOOP_C_238;
      end
      COMP_LOOP_C_238 : begin
        fsm_output = 10'b0100111100;
        state_var_NS = COMP_LOOP_C_239;
      end
      COMP_LOOP_C_239 : begin
        fsm_output = 10'b0100111101;
        state_var_NS = COMP_LOOP_C_240;
      end
      COMP_LOOP_C_240 : begin
        fsm_output = 10'b0100111110;
        state_var_NS = COMP_LOOP_C_241;
      end
      COMP_LOOP_C_241 : begin
        fsm_output = 10'b0100111111;
        state_var_NS = COMP_LOOP_6_modExp_dev_1_while_C_0;
      end
      COMP_LOOP_6_modExp_dev_1_while_C_0 : begin
        fsm_output = 10'b0101000000;
        state_var_NS = COMP_LOOP_6_modExp_dev_1_while_C_1;
      end
      COMP_LOOP_6_modExp_dev_1_while_C_1 : begin
        fsm_output = 10'b0101000001;
        state_var_NS = COMP_LOOP_6_modExp_dev_1_while_C_2;
      end
      COMP_LOOP_6_modExp_dev_1_while_C_2 : begin
        fsm_output = 10'b0101000010;
        state_var_NS = COMP_LOOP_6_modExp_dev_1_while_C_3;
      end
      COMP_LOOP_6_modExp_dev_1_while_C_3 : begin
        fsm_output = 10'b0101000011;
        state_var_NS = COMP_LOOP_6_modExp_dev_1_while_C_4;
      end
      COMP_LOOP_6_modExp_dev_1_while_C_4 : begin
        fsm_output = 10'b0101000100;
        state_var_NS = COMP_LOOP_6_modExp_dev_1_while_C_5;
      end
      COMP_LOOP_6_modExp_dev_1_while_C_5 : begin
        fsm_output = 10'b0101000101;
        state_var_NS = COMP_LOOP_6_modExp_dev_1_while_C_6;
      end
      COMP_LOOP_6_modExp_dev_1_while_C_6 : begin
        fsm_output = 10'b0101000110;
        state_var_NS = COMP_LOOP_6_modExp_dev_1_while_C_7;
      end
      COMP_LOOP_6_modExp_dev_1_while_C_7 : begin
        fsm_output = 10'b0101000111;
        state_var_NS = COMP_LOOP_6_modExp_dev_1_while_C_8;
      end
      COMP_LOOP_6_modExp_dev_1_while_C_8 : begin
        fsm_output = 10'b0101001000;
        state_var_NS = COMP_LOOP_6_modExp_dev_1_while_C_9;
      end
      COMP_LOOP_6_modExp_dev_1_while_C_9 : begin
        fsm_output = 10'b0101001001;
        state_var_NS = COMP_LOOP_6_modExp_dev_1_while_C_10;
      end
      COMP_LOOP_6_modExp_dev_1_while_C_10 : begin
        fsm_output = 10'b0101001010;
        state_var_NS = COMP_LOOP_6_modExp_dev_1_while_C_11;
      end
      COMP_LOOP_6_modExp_dev_1_while_C_11 : begin
        fsm_output = 10'b0101001011;
        if ( COMP_LOOP_6_modExp_dev_1_while_C_11_tr0 ) begin
          state_var_NS = COMP_LOOP_C_242;
        end
        else begin
          state_var_NS = COMP_LOOP_6_modExp_dev_1_while_C_0;
        end
      end
      COMP_LOOP_C_242 : begin
        fsm_output = 10'b0101001100;
        state_var_NS = COMP_LOOP_C_243;
      end
      COMP_LOOP_C_243 : begin
        fsm_output = 10'b0101001101;
        state_var_NS = COMP_LOOP_C_244;
      end
      COMP_LOOP_C_244 : begin
        fsm_output = 10'b0101001110;
        state_var_NS = COMP_LOOP_C_245;
      end
      COMP_LOOP_C_245 : begin
        fsm_output = 10'b0101001111;
        state_var_NS = COMP_LOOP_C_246;
      end
      COMP_LOOP_C_246 : begin
        fsm_output = 10'b0101010000;
        state_var_NS = COMP_LOOP_C_247;
      end
      COMP_LOOP_C_247 : begin
        fsm_output = 10'b0101010001;
        state_var_NS = COMP_LOOP_C_248;
      end
      COMP_LOOP_C_248 : begin
        fsm_output = 10'b0101010010;
        state_var_NS = COMP_LOOP_C_249;
      end
      COMP_LOOP_C_249 : begin
        fsm_output = 10'b0101010011;
        state_var_NS = COMP_LOOP_C_250;
      end
      COMP_LOOP_C_250 : begin
        fsm_output = 10'b0101010100;
        state_var_NS = COMP_LOOP_C_251;
      end
      COMP_LOOP_C_251 : begin
        fsm_output = 10'b0101010101;
        state_var_NS = COMP_LOOP_C_252;
      end
      COMP_LOOP_C_252 : begin
        fsm_output = 10'b0101010110;
        state_var_NS = COMP_LOOP_C_253;
      end
      COMP_LOOP_C_253 : begin
        fsm_output = 10'b0101010111;
        state_var_NS = COMP_LOOP_C_254;
      end
      COMP_LOOP_C_254 : begin
        fsm_output = 10'b0101011000;
        state_var_NS = COMP_LOOP_C_255;
      end
      COMP_LOOP_C_255 : begin
        fsm_output = 10'b0101011001;
        state_var_NS = COMP_LOOP_C_256;
      end
      COMP_LOOP_C_256 : begin
        fsm_output = 10'b0101011010;
        state_var_NS = COMP_LOOP_C_257;
      end
      COMP_LOOP_C_257 : begin
        fsm_output = 10'b0101011011;
        state_var_NS = COMP_LOOP_C_258;
      end
      COMP_LOOP_C_258 : begin
        fsm_output = 10'b0101011100;
        state_var_NS = COMP_LOOP_C_259;
      end
      COMP_LOOP_C_259 : begin
        fsm_output = 10'b0101011101;
        state_var_NS = COMP_LOOP_C_260;
      end
      COMP_LOOP_C_260 : begin
        fsm_output = 10'b0101011110;
        state_var_NS = COMP_LOOP_C_261;
      end
      COMP_LOOP_C_261 : begin
        fsm_output = 10'b0101011111;
        state_var_NS = COMP_LOOP_C_262;
      end
      COMP_LOOP_C_262 : begin
        fsm_output = 10'b0101100000;
        state_var_NS = COMP_LOOP_C_263;
      end
      COMP_LOOP_C_263 : begin
        fsm_output = 10'b0101100001;
        state_var_NS = COMP_LOOP_C_264;
      end
      COMP_LOOP_C_264 : begin
        fsm_output = 10'b0101100010;
        state_var_NS = COMP_LOOP_C_265;
      end
      COMP_LOOP_C_265 : begin
        fsm_output = 10'b0101100011;
        state_var_NS = COMP_LOOP_C_266;
      end
      COMP_LOOP_C_266 : begin
        fsm_output = 10'b0101100100;
        state_var_NS = COMP_LOOP_C_267;
      end
      COMP_LOOP_C_267 : begin
        fsm_output = 10'b0101100101;
        state_var_NS = COMP_LOOP_C_268;
      end
      COMP_LOOP_C_268 : begin
        fsm_output = 10'b0101100110;
        state_var_NS = COMP_LOOP_C_269;
      end
      COMP_LOOP_C_269 : begin
        fsm_output = 10'b0101100111;
        state_var_NS = COMP_LOOP_C_270;
      end
      COMP_LOOP_C_270 : begin
        fsm_output = 10'b0101101000;
        if ( COMP_LOOP_C_270_tr0 ) begin
          state_var_NS = STAGE_VEC_LOOP_C_1;
        end
        else begin
          state_var_NS = COMP_LOOP_C_271;
        end
      end
      COMP_LOOP_C_271 : begin
        fsm_output = 10'b0101101001;
        state_var_NS = COMP_LOOP_C_272;
      end
      COMP_LOOP_C_272 : begin
        fsm_output = 10'b0101101010;
        state_var_NS = COMP_LOOP_C_273;
      end
      COMP_LOOP_C_273 : begin
        fsm_output = 10'b0101101011;
        state_var_NS = COMP_LOOP_C_274;
      end
      COMP_LOOP_C_274 : begin
        fsm_output = 10'b0101101100;
        state_var_NS = COMP_LOOP_C_275;
      end
      COMP_LOOP_C_275 : begin
        fsm_output = 10'b0101101101;
        state_var_NS = COMP_LOOP_C_276;
      end
      COMP_LOOP_C_276 : begin
        fsm_output = 10'b0101101110;
        state_var_NS = COMP_LOOP_C_277;
      end
      COMP_LOOP_C_277 : begin
        fsm_output = 10'b0101101111;
        state_var_NS = COMP_LOOP_C_278;
      end
      COMP_LOOP_C_278 : begin
        fsm_output = 10'b0101110000;
        state_var_NS = COMP_LOOP_C_279;
      end
      COMP_LOOP_C_279 : begin
        fsm_output = 10'b0101110001;
        state_var_NS = COMP_LOOP_C_280;
      end
      COMP_LOOP_C_280 : begin
        fsm_output = 10'b0101110010;
        state_var_NS = COMP_LOOP_C_281;
      end
      COMP_LOOP_C_281 : begin
        fsm_output = 10'b0101110011;
        state_var_NS = COMP_LOOP_C_282;
      end
      COMP_LOOP_C_282 : begin
        fsm_output = 10'b0101110100;
        state_var_NS = COMP_LOOP_C_283;
      end
      COMP_LOOP_C_283 : begin
        fsm_output = 10'b0101110101;
        state_var_NS = COMP_LOOP_C_284;
      end
      COMP_LOOP_C_284 : begin
        fsm_output = 10'b0101110110;
        state_var_NS = COMP_LOOP_C_285;
      end
      COMP_LOOP_C_285 : begin
        fsm_output = 10'b0101110111;
        state_var_NS = COMP_LOOP_C_286;
      end
      COMP_LOOP_C_286 : begin
        fsm_output = 10'b0101111000;
        state_var_NS = COMP_LOOP_7_modExp_dev_1_while_C_0;
      end
      COMP_LOOP_7_modExp_dev_1_while_C_0 : begin
        fsm_output = 10'b0101111001;
        state_var_NS = COMP_LOOP_7_modExp_dev_1_while_C_1;
      end
      COMP_LOOP_7_modExp_dev_1_while_C_1 : begin
        fsm_output = 10'b0101111010;
        state_var_NS = COMP_LOOP_7_modExp_dev_1_while_C_2;
      end
      COMP_LOOP_7_modExp_dev_1_while_C_2 : begin
        fsm_output = 10'b0101111011;
        state_var_NS = COMP_LOOP_7_modExp_dev_1_while_C_3;
      end
      COMP_LOOP_7_modExp_dev_1_while_C_3 : begin
        fsm_output = 10'b0101111100;
        state_var_NS = COMP_LOOP_7_modExp_dev_1_while_C_4;
      end
      COMP_LOOP_7_modExp_dev_1_while_C_4 : begin
        fsm_output = 10'b0101111101;
        state_var_NS = COMP_LOOP_7_modExp_dev_1_while_C_5;
      end
      COMP_LOOP_7_modExp_dev_1_while_C_5 : begin
        fsm_output = 10'b0101111110;
        state_var_NS = COMP_LOOP_7_modExp_dev_1_while_C_6;
      end
      COMP_LOOP_7_modExp_dev_1_while_C_6 : begin
        fsm_output = 10'b0101111111;
        state_var_NS = COMP_LOOP_7_modExp_dev_1_while_C_7;
      end
      COMP_LOOP_7_modExp_dev_1_while_C_7 : begin
        fsm_output = 10'b0110000000;
        state_var_NS = COMP_LOOP_7_modExp_dev_1_while_C_8;
      end
      COMP_LOOP_7_modExp_dev_1_while_C_8 : begin
        fsm_output = 10'b0110000001;
        state_var_NS = COMP_LOOP_7_modExp_dev_1_while_C_9;
      end
      COMP_LOOP_7_modExp_dev_1_while_C_9 : begin
        fsm_output = 10'b0110000010;
        state_var_NS = COMP_LOOP_7_modExp_dev_1_while_C_10;
      end
      COMP_LOOP_7_modExp_dev_1_while_C_10 : begin
        fsm_output = 10'b0110000011;
        state_var_NS = COMP_LOOP_7_modExp_dev_1_while_C_11;
      end
      COMP_LOOP_7_modExp_dev_1_while_C_11 : begin
        fsm_output = 10'b0110000100;
        if ( COMP_LOOP_7_modExp_dev_1_while_C_11_tr0 ) begin
          state_var_NS = COMP_LOOP_C_287;
        end
        else begin
          state_var_NS = COMP_LOOP_7_modExp_dev_1_while_C_0;
        end
      end
      COMP_LOOP_C_287 : begin
        fsm_output = 10'b0110000101;
        state_var_NS = COMP_LOOP_C_288;
      end
      COMP_LOOP_C_288 : begin
        fsm_output = 10'b0110000110;
        state_var_NS = COMP_LOOP_C_289;
      end
      COMP_LOOP_C_289 : begin
        fsm_output = 10'b0110000111;
        state_var_NS = COMP_LOOP_C_290;
      end
      COMP_LOOP_C_290 : begin
        fsm_output = 10'b0110001000;
        state_var_NS = COMP_LOOP_C_291;
      end
      COMP_LOOP_C_291 : begin
        fsm_output = 10'b0110001001;
        state_var_NS = COMP_LOOP_C_292;
      end
      COMP_LOOP_C_292 : begin
        fsm_output = 10'b0110001010;
        state_var_NS = COMP_LOOP_C_293;
      end
      COMP_LOOP_C_293 : begin
        fsm_output = 10'b0110001011;
        state_var_NS = COMP_LOOP_C_294;
      end
      COMP_LOOP_C_294 : begin
        fsm_output = 10'b0110001100;
        state_var_NS = COMP_LOOP_C_295;
      end
      COMP_LOOP_C_295 : begin
        fsm_output = 10'b0110001101;
        state_var_NS = COMP_LOOP_C_296;
      end
      COMP_LOOP_C_296 : begin
        fsm_output = 10'b0110001110;
        state_var_NS = COMP_LOOP_C_297;
      end
      COMP_LOOP_C_297 : begin
        fsm_output = 10'b0110001111;
        state_var_NS = COMP_LOOP_C_298;
      end
      COMP_LOOP_C_298 : begin
        fsm_output = 10'b0110010000;
        state_var_NS = COMP_LOOP_C_299;
      end
      COMP_LOOP_C_299 : begin
        fsm_output = 10'b0110010001;
        state_var_NS = COMP_LOOP_C_300;
      end
      COMP_LOOP_C_300 : begin
        fsm_output = 10'b0110010010;
        state_var_NS = COMP_LOOP_C_301;
      end
      COMP_LOOP_C_301 : begin
        fsm_output = 10'b0110010011;
        state_var_NS = COMP_LOOP_C_302;
      end
      COMP_LOOP_C_302 : begin
        fsm_output = 10'b0110010100;
        state_var_NS = COMP_LOOP_C_303;
      end
      COMP_LOOP_C_303 : begin
        fsm_output = 10'b0110010101;
        state_var_NS = COMP_LOOP_C_304;
      end
      COMP_LOOP_C_304 : begin
        fsm_output = 10'b0110010110;
        state_var_NS = COMP_LOOP_C_305;
      end
      COMP_LOOP_C_305 : begin
        fsm_output = 10'b0110010111;
        state_var_NS = COMP_LOOP_C_306;
      end
      COMP_LOOP_C_306 : begin
        fsm_output = 10'b0110011000;
        state_var_NS = COMP_LOOP_C_307;
      end
      COMP_LOOP_C_307 : begin
        fsm_output = 10'b0110011001;
        state_var_NS = COMP_LOOP_C_308;
      end
      COMP_LOOP_C_308 : begin
        fsm_output = 10'b0110011010;
        state_var_NS = COMP_LOOP_C_309;
      end
      COMP_LOOP_C_309 : begin
        fsm_output = 10'b0110011011;
        state_var_NS = COMP_LOOP_C_310;
      end
      COMP_LOOP_C_310 : begin
        fsm_output = 10'b0110011100;
        state_var_NS = COMP_LOOP_C_311;
      end
      COMP_LOOP_C_311 : begin
        fsm_output = 10'b0110011101;
        state_var_NS = COMP_LOOP_C_312;
      end
      COMP_LOOP_C_312 : begin
        fsm_output = 10'b0110011110;
        state_var_NS = COMP_LOOP_C_313;
      end
      COMP_LOOP_C_313 : begin
        fsm_output = 10'b0110011111;
        state_var_NS = COMP_LOOP_C_314;
      end
      COMP_LOOP_C_314 : begin
        fsm_output = 10'b0110100000;
        state_var_NS = COMP_LOOP_C_315;
      end
      COMP_LOOP_C_315 : begin
        fsm_output = 10'b0110100001;
        if ( COMP_LOOP_C_315_tr0 ) begin
          state_var_NS = STAGE_VEC_LOOP_C_1;
        end
        else begin
          state_var_NS = COMP_LOOP_C_316;
        end
      end
      COMP_LOOP_C_316 : begin
        fsm_output = 10'b0110100010;
        state_var_NS = COMP_LOOP_C_317;
      end
      COMP_LOOP_C_317 : begin
        fsm_output = 10'b0110100011;
        state_var_NS = COMP_LOOP_C_318;
      end
      COMP_LOOP_C_318 : begin
        fsm_output = 10'b0110100100;
        state_var_NS = COMP_LOOP_C_319;
      end
      COMP_LOOP_C_319 : begin
        fsm_output = 10'b0110100101;
        state_var_NS = COMP_LOOP_C_320;
      end
      COMP_LOOP_C_320 : begin
        fsm_output = 10'b0110100110;
        state_var_NS = COMP_LOOP_C_321;
      end
      COMP_LOOP_C_321 : begin
        fsm_output = 10'b0110100111;
        state_var_NS = COMP_LOOP_C_322;
      end
      COMP_LOOP_C_322 : begin
        fsm_output = 10'b0110101000;
        state_var_NS = COMP_LOOP_C_323;
      end
      COMP_LOOP_C_323 : begin
        fsm_output = 10'b0110101001;
        state_var_NS = COMP_LOOP_C_324;
      end
      COMP_LOOP_C_324 : begin
        fsm_output = 10'b0110101010;
        state_var_NS = COMP_LOOP_C_325;
      end
      COMP_LOOP_C_325 : begin
        fsm_output = 10'b0110101011;
        state_var_NS = COMP_LOOP_C_326;
      end
      COMP_LOOP_C_326 : begin
        fsm_output = 10'b0110101100;
        state_var_NS = COMP_LOOP_C_327;
      end
      COMP_LOOP_C_327 : begin
        fsm_output = 10'b0110101101;
        state_var_NS = COMP_LOOP_C_328;
      end
      COMP_LOOP_C_328 : begin
        fsm_output = 10'b0110101110;
        state_var_NS = COMP_LOOP_C_329;
      end
      COMP_LOOP_C_329 : begin
        fsm_output = 10'b0110101111;
        state_var_NS = COMP_LOOP_C_330;
      end
      COMP_LOOP_C_330 : begin
        fsm_output = 10'b0110110000;
        state_var_NS = COMP_LOOP_C_331;
      end
      COMP_LOOP_C_331 : begin
        fsm_output = 10'b0110110001;
        state_var_NS = COMP_LOOP_8_modExp_dev_1_while_C_0;
      end
      COMP_LOOP_8_modExp_dev_1_while_C_0 : begin
        fsm_output = 10'b0110110010;
        state_var_NS = COMP_LOOP_8_modExp_dev_1_while_C_1;
      end
      COMP_LOOP_8_modExp_dev_1_while_C_1 : begin
        fsm_output = 10'b0110110011;
        state_var_NS = COMP_LOOP_8_modExp_dev_1_while_C_2;
      end
      COMP_LOOP_8_modExp_dev_1_while_C_2 : begin
        fsm_output = 10'b0110110100;
        state_var_NS = COMP_LOOP_8_modExp_dev_1_while_C_3;
      end
      COMP_LOOP_8_modExp_dev_1_while_C_3 : begin
        fsm_output = 10'b0110110101;
        state_var_NS = COMP_LOOP_8_modExp_dev_1_while_C_4;
      end
      COMP_LOOP_8_modExp_dev_1_while_C_4 : begin
        fsm_output = 10'b0110110110;
        state_var_NS = COMP_LOOP_8_modExp_dev_1_while_C_5;
      end
      COMP_LOOP_8_modExp_dev_1_while_C_5 : begin
        fsm_output = 10'b0110110111;
        state_var_NS = COMP_LOOP_8_modExp_dev_1_while_C_6;
      end
      COMP_LOOP_8_modExp_dev_1_while_C_6 : begin
        fsm_output = 10'b0110111000;
        state_var_NS = COMP_LOOP_8_modExp_dev_1_while_C_7;
      end
      COMP_LOOP_8_modExp_dev_1_while_C_7 : begin
        fsm_output = 10'b0110111001;
        state_var_NS = COMP_LOOP_8_modExp_dev_1_while_C_8;
      end
      COMP_LOOP_8_modExp_dev_1_while_C_8 : begin
        fsm_output = 10'b0110111010;
        state_var_NS = COMP_LOOP_8_modExp_dev_1_while_C_9;
      end
      COMP_LOOP_8_modExp_dev_1_while_C_9 : begin
        fsm_output = 10'b0110111011;
        state_var_NS = COMP_LOOP_8_modExp_dev_1_while_C_10;
      end
      COMP_LOOP_8_modExp_dev_1_while_C_10 : begin
        fsm_output = 10'b0110111100;
        state_var_NS = COMP_LOOP_8_modExp_dev_1_while_C_11;
      end
      COMP_LOOP_8_modExp_dev_1_while_C_11 : begin
        fsm_output = 10'b0110111101;
        if ( COMP_LOOP_8_modExp_dev_1_while_C_11_tr0 ) begin
          state_var_NS = COMP_LOOP_C_332;
        end
        else begin
          state_var_NS = COMP_LOOP_8_modExp_dev_1_while_C_0;
        end
      end
      COMP_LOOP_C_332 : begin
        fsm_output = 10'b0110111110;
        state_var_NS = COMP_LOOP_C_333;
      end
      COMP_LOOP_C_333 : begin
        fsm_output = 10'b0110111111;
        state_var_NS = COMP_LOOP_C_334;
      end
      COMP_LOOP_C_334 : begin
        fsm_output = 10'b0111000000;
        state_var_NS = COMP_LOOP_C_335;
      end
      COMP_LOOP_C_335 : begin
        fsm_output = 10'b0111000001;
        state_var_NS = COMP_LOOP_C_336;
      end
      COMP_LOOP_C_336 : begin
        fsm_output = 10'b0111000010;
        state_var_NS = COMP_LOOP_C_337;
      end
      COMP_LOOP_C_337 : begin
        fsm_output = 10'b0111000011;
        state_var_NS = COMP_LOOP_C_338;
      end
      COMP_LOOP_C_338 : begin
        fsm_output = 10'b0111000100;
        state_var_NS = COMP_LOOP_C_339;
      end
      COMP_LOOP_C_339 : begin
        fsm_output = 10'b0111000101;
        state_var_NS = COMP_LOOP_C_340;
      end
      COMP_LOOP_C_340 : begin
        fsm_output = 10'b0111000110;
        state_var_NS = COMP_LOOP_C_341;
      end
      COMP_LOOP_C_341 : begin
        fsm_output = 10'b0111000111;
        state_var_NS = COMP_LOOP_C_342;
      end
      COMP_LOOP_C_342 : begin
        fsm_output = 10'b0111001000;
        state_var_NS = COMP_LOOP_C_343;
      end
      COMP_LOOP_C_343 : begin
        fsm_output = 10'b0111001001;
        state_var_NS = COMP_LOOP_C_344;
      end
      COMP_LOOP_C_344 : begin
        fsm_output = 10'b0111001010;
        state_var_NS = COMP_LOOP_C_345;
      end
      COMP_LOOP_C_345 : begin
        fsm_output = 10'b0111001011;
        state_var_NS = COMP_LOOP_C_346;
      end
      COMP_LOOP_C_346 : begin
        fsm_output = 10'b0111001100;
        state_var_NS = COMP_LOOP_C_347;
      end
      COMP_LOOP_C_347 : begin
        fsm_output = 10'b0111001101;
        state_var_NS = COMP_LOOP_C_348;
      end
      COMP_LOOP_C_348 : begin
        fsm_output = 10'b0111001110;
        state_var_NS = COMP_LOOP_C_349;
      end
      COMP_LOOP_C_349 : begin
        fsm_output = 10'b0111001111;
        state_var_NS = COMP_LOOP_C_350;
      end
      COMP_LOOP_C_350 : begin
        fsm_output = 10'b0111010000;
        state_var_NS = COMP_LOOP_C_351;
      end
      COMP_LOOP_C_351 : begin
        fsm_output = 10'b0111010001;
        state_var_NS = COMP_LOOP_C_352;
      end
      COMP_LOOP_C_352 : begin
        fsm_output = 10'b0111010010;
        state_var_NS = COMP_LOOP_C_353;
      end
      COMP_LOOP_C_353 : begin
        fsm_output = 10'b0111010011;
        state_var_NS = COMP_LOOP_C_354;
      end
      COMP_LOOP_C_354 : begin
        fsm_output = 10'b0111010100;
        state_var_NS = COMP_LOOP_C_355;
      end
      COMP_LOOP_C_355 : begin
        fsm_output = 10'b0111010101;
        state_var_NS = COMP_LOOP_C_356;
      end
      COMP_LOOP_C_356 : begin
        fsm_output = 10'b0111010110;
        state_var_NS = COMP_LOOP_C_357;
      end
      COMP_LOOP_C_357 : begin
        fsm_output = 10'b0111010111;
        state_var_NS = COMP_LOOP_C_358;
      end
      COMP_LOOP_C_358 : begin
        fsm_output = 10'b0111011000;
        state_var_NS = COMP_LOOP_C_359;
      end
      COMP_LOOP_C_359 : begin
        fsm_output = 10'b0111011001;
        state_var_NS = COMP_LOOP_C_360;
      end
      COMP_LOOP_C_360 : begin
        fsm_output = 10'b0111011010;
        if ( COMP_LOOP_C_360_tr0 ) begin
          state_var_NS = STAGE_VEC_LOOP_C_1;
        end
        else begin
          state_var_NS = COMP_LOOP_C_361;
        end
      end
      COMP_LOOP_C_361 : begin
        fsm_output = 10'b0111011011;
        state_var_NS = COMP_LOOP_C_362;
      end
      COMP_LOOP_C_362 : begin
        fsm_output = 10'b0111011100;
        state_var_NS = COMP_LOOP_C_363;
      end
      COMP_LOOP_C_363 : begin
        fsm_output = 10'b0111011101;
        state_var_NS = COMP_LOOP_C_364;
      end
      COMP_LOOP_C_364 : begin
        fsm_output = 10'b0111011110;
        state_var_NS = COMP_LOOP_C_365;
      end
      COMP_LOOP_C_365 : begin
        fsm_output = 10'b0111011111;
        state_var_NS = COMP_LOOP_C_366;
      end
      COMP_LOOP_C_366 : begin
        fsm_output = 10'b0111100000;
        state_var_NS = COMP_LOOP_C_367;
      end
      COMP_LOOP_C_367 : begin
        fsm_output = 10'b0111100001;
        state_var_NS = COMP_LOOP_C_368;
      end
      COMP_LOOP_C_368 : begin
        fsm_output = 10'b0111100010;
        state_var_NS = COMP_LOOP_C_369;
      end
      COMP_LOOP_C_369 : begin
        fsm_output = 10'b0111100011;
        state_var_NS = COMP_LOOP_C_370;
      end
      COMP_LOOP_C_370 : begin
        fsm_output = 10'b0111100100;
        state_var_NS = COMP_LOOP_C_371;
      end
      COMP_LOOP_C_371 : begin
        fsm_output = 10'b0111100101;
        state_var_NS = COMP_LOOP_C_372;
      end
      COMP_LOOP_C_372 : begin
        fsm_output = 10'b0111100110;
        state_var_NS = COMP_LOOP_C_373;
      end
      COMP_LOOP_C_373 : begin
        fsm_output = 10'b0111100111;
        state_var_NS = COMP_LOOP_C_374;
      end
      COMP_LOOP_C_374 : begin
        fsm_output = 10'b0111101000;
        state_var_NS = COMP_LOOP_C_375;
      end
      COMP_LOOP_C_375 : begin
        fsm_output = 10'b0111101001;
        state_var_NS = COMP_LOOP_C_376;
      end
      COMP_LOOP_C_376 : begin
        fsm_output = 10'b0111101010;
        state_var_NS = COMP_LOOP_9_modExp_dev_1_while_C_0;
      end
      COMP_LOOP_9_modExp_dev_1_while_C_0 : begin
        fsm_output = 10'b0111101011;
        state_var_NS = COMP_LOOP_9_modExp_dev_1_while_C_1;
      end
      COMP_LOOP_9_modExp_dev_1_while_C_1 : begin
        fsm_output = 10'b0111101100;
        state_var_NS = COMP_LOOP_9_modExp_dev_1_while_C_2;
      end
      COMP_LOOP_9_modExp_dev_1_while_C_2 : begin
        fsm_output = 10'b0111101101;
        state_var_NS = COMP_LOOP_9_modExp_dev_1_while_C_3;
      end
      COMP_LOOP_9_modExp_dev_1_while_C_3 : begin
        fsm_output = 10'b0111101110;
        state_var_NS = COMP_LOOP_9_modExp_dev_1_while_C_4;
      end
      COMP_LOOP_9_modExp_dev_1_while_C_4 : begin
        fsm_output = 10'b0111101111;
        state_var_NS = COMP_LOOP_9_modExp_dev_1_while_C_5;
      end
      COMP_LOOP_9_modExp_dev_1_while_C_5 : begin
        fsm_output = 10'b0111110000;
        state_var_NS = COMP_LOOP_9_modExp_dev_1_while_C_6;
      end
      COMP_LOOP_9_modExp_dev_1_while_C_6 : begin
        fsm_output = 10'b0111110001;
        state_var_NS = COMP_LOOP_9_modExp_dev_1_while_C_7;
      end
      COMP_LOOP_9_modExp_dev_1_while_C_7 : begin
        fsm_output = 10'b0111110010;
        state_var_NS = COMP_LOOP_9_modExp_dev_1_while_C_8;
      end
      COMP_LOOP_9_modExp_dev_1_while_C_8 : begin
        fsm_output = 10'b0111110011;
        state_var_NS = COMP_LOOP_9_modExp_dev_1_while_C_9;
      end
      COMP_LOOP_9_modExp_dev_1_while_C_9 : begin
        fsm_output = 10'b0111110100;
        state_var_NS = COMP_LOOP_9_modExp_dev_1_while_C_10;
      end
      COMP_LOOP_9_modExp_dev_1_while_C_10 : begin
        fsm_output = 10'b0111110101;
        state_var_NS = COMP_LOOP_9_modExp_dev_1_while_C_11;
      end
      COMP_LOOP_9_modExp_dev_1_while_C_11 : begin
        fsm_output = 10'b0111110110;
        if ( COMP_LOOP_9_modExp_dev_1_while_C_11_tr0 ) begin
          state_var_NS = COMP_LOOP_C_377;
        end
        else begin
          state_var_NS = COMP_LOOP_9_modExp_dev_1_while_C_0;
        end
      end
      COMP_LOOP_C_377 : begin
        fsm_output = 10'b0111110111;
        state_var_NS = COMP_LOOP_C_378;
      end
      COMP_LOOP_C_378 : begin
        fsm_output = 10'b0111111000;
        state_var_NS = COMP_LOOP_C_379;
      end
      COMP_LOOP_C_379 : begin
        fsm_output = 10'b0111111001;
        state_var_NS = COMP_LOOP_C_380;
      end
      COMP_LOOP_C_380 : begin
        fsm_output = 10'b0111111010;
        state_var_NS = COMP_LOOP_C_381;
      end
      COMP_LOOP_C_381 : begin
        fsm_output = 10'b0111111011;
        state_var_NS = COMP_LOOP_C_382;
      end
      COMP_LOOP_C_382 : begin
        fsm_output = 10'b0111111100;
        state_var_NS = COMP_LOOP_C_383;
      end
      COMP_LOOP_C_383 : begin
        fsm_output = 10'b0111111101;
        state_var_NS = COMP_LOOP_C_384;
      end
      COMP_LOOP_C_384 : begin
        fsm_output = 10'b0111111110;
        state_var_NS = COMP_LOOP_C_385;
      end
      COMP_LOOP_C_385 : begin
        fsm_output = 10'b0111111111;
        state_var_NS = COMP_LOOP_C_386;
      end
      COMP_LOOP_C_386 : begin
        fsm_output = 10'b1000000000;
        state_var_NS = COMP_LOOP_C_387;
      end
      COMP_LOOP_C_387 : begin
        fsm_output = 10'b1000000001;
        state_var_NS = COMP_LOOP_C_388;
      end
      COMP_LOOP_C_388 : begin
        fsm_output = 10'b1000000010;
        state_var_NS = COMP_LOOP_C_389;
      end
      COMP_LOOP_C_389 : begin
        fsm_output = 10'b1000000011;
        state_var_NS = COMP_LOOP_C_390;
      end
      COMP_LOOP_C_390 : begin
        fsm_output = 10'b1000000100;
        state_var_NS = COMP_LOOP_C_391;
      end
      COMP_LOOP_C_391 : begin
        fsm_output = 10'b1000000101;
        state_var_NS = COMP_LOOP_C_392;
      end
      COMP_LOOP_C_392 : begin
        fsm_output = 10'b1000000110;
        state_var_NS = COMP_LOOP_C_393;
      end
      COMP_LOOP_C_393 : begin
        fsm_output = 10'b1000000111;
        state_var_NS = COMP_LOOP_C_394;
      end
      COMP_LOOP_C_394 : begin
        fsm_output = 10'b1000001000;
        state_var_NS = COMP_LOOP_C_395;
      end
      COMP_LOOP_C_395 : begin
        fsm_output = 10'b1000001001;
        state_var_NS = COMP_LOOP_C_396;
      end
      COMP_LOOP_C_396 : begin
        fsm_output = 10'b1000001010;
        state_var_NS = COMP_LOOP_C_397;
      end
      COMP_LOOP_C_397 : begin
        fsm_output = 10'b1000001011;
        state_var_NS = COMP_LOOP_C_398;
      end
      COMP_LOOP_C_398 : begin
        fsm_output = 10'b1000001100;
        state_var_NS = COMP_LOOP_C_399;
      end
      COMP_LOOP_C_399 : begin
        fsm_output = 10'b1000001101;
        state_var_NS = COMP_LOOP_C_400;
      end
      COMP_LOOP_C_400 : begin
        fsm_output = 10'b1000001110;
        state_var_NS = COMP_LOOP_C_401;
      end
      COMP_LOOP_C_401 : begin
        fsm_output = 10'b1000001111;
        state_var_NS = COMP_LOOP_C_402;
      end
      COMP_LOOP_C_402 : begin
        fsm_output = 10'b1000010000;
        state_var_NS = COMP_LOOP_C_403;
      end
      COMP_LOOP_C_403 : begin
        fsm_output = 10'b1000010001;
        state_var_NS = COMP_LOOP_C_404;
      end
      COMP_LOOP_C_404 : begin
        fsm_output = 10'b1000010010;
        state_var_NS = COMP_LOOP_C_405;
      end
      COMP_LOOP_C_405 : begin
        fsm_output = 10'b1000010011;
        if ( COMP_LOOP_C_405_tr0 ) begin
          state_var_NS = STAGE_VEC_LOOP_C_1;
        end
        else begin
          state_var_NS = COMP_LOOP_C_406;
        end
      end
      COMP_LOOP_C_406 : begin
        fsm_output = 10'b1000010100;
        state_var_NS = COMP_LOOP_C_407;
      end
      COMP_LOOP_C_407 : begin
        fsm_output = 10'b1000010101;
        state_var_NS = COMP_LOOP_C_408;
      end
      COMP_LOOP_C_408 : begin
        fsm_output = 10'b1000010110;
        state_var_NS = COMP_LOOP_C_409;
      end
      COMP_LOOP_C_409 : begin
        fsm_output = 10'b1000010111;
        state_var_NS = COMP_LOOP_C_410;
      end
      COMP_LOOP_C_410 : begin
        fsm_output = 10'b1000011000;
        state_var_NS = COMP_LOOP_C_411;
      end
      COMP_LOOP_C_411 : begin
        fsm_output = 10'b1000011001;
        state_var_NS = COMP_LOOP_C_412;
      end
      COMP_LOOP_C_412 : begin
        fsm_output = 10'b1000011010;
        state_var_NS = COMP_LOOP_C_413;
      end
      COMP_LOOP_C_413 : begin
        fsm_output = 10'b1000011011;
        state_var_NS = COMP_LOOP_C_414;
      end
      COMP_LOOP_C_414 : begin
        fsm_output = 10'b1000011100;
        state_var_NS = COMP_LOOP_C_415;
      end
      COMP_LOOP_C_415 : begin
        fsm_output = 10'b1000011101;
        state_var_NS = COMP_LOOP_C_416;
      end
      COMP_LOOP_C_416 : begin
        fsm_output = 10'b1000011110;
        state_var_NS = COMP_LOOP_C_417;
      end
      COMP_LOOP_C_417 : begin
        fsm_output = 10'b1000011111;
        state_var_NS = COMP_LOOP_C_418;
      end
      COMP_LOOP_C_418 : begin
        fsm_output = 10'b1000100000;
        state_var_NS = COMP_LOOP_C_419;
      end
      COMP_LOOP_C_419 : begin
        fsm_output = 10'b1000100001;
        state_var_NS = COMP_LOOP_C_420;
      end
      COMP_LOOP_C_420 : begin
        fsm_output = 10'b1000100010;
        state_var_NS = COMP_LOOP_C_421;
      end
      COMP_LOOP_C_421 : begin
        fsm_output = 10'b1000100011;
        state_var_NS = COMP_LOOP_10_modExp_dev_1_while_C_0;
      end
      COMP_LOOP_10_modExp_dev_1_while_C_0 : begin
        fsm_output = 10'b1000100100;
        state_var_NS = COMP_LOOP_10_modExp_dev_1_while_C_1;
      end
      COMP_LOOP_10_modExp_dev_1_while_C_1 : begin
        fsm_output = 10'b1000100101;
        state_var_NS = COMP_LOOP_10_modExp_dev_1_while_C_2;
      end
      COMP_LOOP_10_modExp_dev_1_while_C_2 : begin
        fsm_output = 10'b1000100110;
        state_var_NS = COMP_LOOP_10_modExp_dev_1_while_C_3;
      end
      COMP_LOOP_10_modExp_dev_1_while_C_3 : begin
        fsm_output = 10'b1000100111;
        state_var_NS = COMP_LOOP_10_modExp_dev_1_while_C_4;
      end
      COMP_LOOP_10_modExp_dev_1_while_C_4 : begin
        fsm_output = 10'b1000101000;
        state_var_NS = COMP_LOOP_10_modExp_dev_1_while_C_5;
      end
      COMP_LOOP_10_modExp_dev_1_while_C_5 : begin
        fsm_output = 10'b1000101001;
        state_var_NS = COMP_LOOP_10_modExp_dev_1_while_C_6;
      end
      COMP_LOOP_10_modExp_dev_1_while_C_6 : begin
        fsm_output = 10'b1000101010;
        state_var_NS = COMP_LOOP_10_modExp_dev_1_while_C_7;
      end
      COMP_LOOP_10_modExp_dev_1_while_C_7 : begin
        fsm_output = 10'b1000101011;
        state_var_NS = COMP_LOOP_10_modExp_dev_1_while_C_8;
      end
      COMP_LOOP_10_modExp_dev_1_while_C_8 : begin
        fsm_output = 10'b1000101100;
        state_var_NS = COMP_LOOP_10_modExp_dev_1_while_C_9;
      end
      COMP_LOOP_10_modExp_dev_1_while_C_9 : begin
        fsm_output = 10'b1000101101;
        state_var_NS = COMP_LOOP_10_modExp_dev_1_while_C_10;
      end
      COMP_LOOP_10_modExp_dev_1_while_C_10 : begin
        fsm_output = 10'b1000101110;
        state_var_NS = COMP_LOOP_10_modExp_dev_1_while_C_11;
      end
      COMP_LOOP_10_modExp_dev_1_while_C_11 : begin
        fsm_output = 10'b1000101111;
        if ( COMP_LOOP_10_modExp_dev_1_while_C_11_tr0 ) begin
          state_var_NS = COMP_LOOP_C_422;
        end
        else begin
          state_var_NS = COMP_LOOP_10_modExp_dev_1_while_C_0;
        end
      end
      COMP_LOOP_C_422 : begin
        fsm_output = 10'b1000110000;
        state_var_NS = COMP_LOOP_C_423;
      end
      COMP_LOOP_C_423 : begin
        fsm_output = 10'b1000110001;
        state_var_NS = COMP_LOOP_C_424;
      end
      COMP_LOOP_C_424 : begin
        fsm_output = 10'b1000110010;
        state_var_NS = COMP_LOOP_C_425;
      end
      COMP_LOOP_C_425 : begin
        fsm_output = 10'b1000110011;
        state_var_NS = COMP_LOOP_C_426;
      end
      COMP_LOOP_C_426 : begin
        fsm_output = 10'b1000110100;
        state_var_NS = COMP_LOOP_C_427;
      end
      COMP_LOOP_C_427 : begin
        fsm_output = 10'b1000110101;
        state_var_NS = COMP_LOOP_C_428;
      end
      COMP_LOOP_C_428 : begin
        fsm_output = 10'b1000110110;
        state_var_NS = COMP_LOOP_C_429;
      end
      COMP_LOOP_C_429 : begin
        fsm_output = 10'b1000110111;
        state_var_NS = COMP_LOOP_C_430;
      end
      COMP_LOOP_C_430 : begin
        fsm_output = 10'b1000111000;
        state_var_NS = COMP_LOOP_C_431;
      end
      COMP_LOOP_C_431 : begin
        fsm_output = 10'b1000111001;
        state_var_NS = COMP_LOOP_C_432;
      end
      COMP_LOOP_C_432 : begin
        fsm_output = 10'b1000111010;
        state_var_NS = COMP_LOOP_C_433;
      end
      COMP_LOOP_C_433 : begin
        fsm_output = 10'b1000111011;
        state_var_NS = COMP_LOOP_C_434;
      end
      COMP_LOOP_C_434 : begin
        fsm_output = 10'b1000111100;
        state_var_NS = COMP_LOOP_C_435;
      end
      COMP_LOOP_C_435 : begin
        fsm_output = 10'b1000111101;
        state_var_NS = COMP_LOOP_C_436;
      end
      COMP_LOOP_C_436 : begin
        fsm_output = 10'b1000111110;
        state_var_NS = COMP_LOOP_C_437;
      end
      COMP_LOOP_C_437 : begin
        fsm_output = 10'b1000111111;
        state_var_NS = COMP_LOOP_C_438;
      end
      COMP_LOOP_C_438 : begin
        fsm_output = 10'b1001000000;
        state_var_NS = COMP_LOOP_C_439;
      end
      COMP_LOOP_C_439 : begin
        fsm_output = 10'b1001000001;
        state_var_NS = COMP_LOOP_C_440;
      end
      COMP_LOOP_C_440 : begin
        fsm_output = 10'b1001000010;
        state_var_NS = COMP_LOOP_C_441;
      end
      COMP_LOOP_C_441 : begin
        fsm_output = 10'b1001000011;
        state_var_NS = COMP_LOOP_C_442;
      end
      COMP_LOOP_C_442 : begin
        fsm_output = 10'b1001000100;
        state_var_NS = COMP_LOOP_C_443;
      end
      COMP_LOOP_C_443 : begin
        fsm_output = 10'b1001000101;
        state_var_NS = COMP_LOOP_C_444;
      end
      COMP_LOOP_C_444 : begin
        fsm_output = 10'b1001000110;
        state_var_NS = COMP_LOOP_C_445;
      end
      COMP_LOOP_C_445 : begin
        fsm_output = 10'b1001000111;
        state_var_NS = COMP_LOOP_C_446;
      end
      COMP_LOOP_C_446 : begin
        fsm_output = 10'b1001001000;
        state_var_NS = COMP_LOOP_C_447;
      end
      COMP_LOOP_C_447 : begin
        fsm_output = 10'b1001001001;
        state_var_NS = COMP_LOOP_C_448;
      end
      COMP_LOOP_C_448 : begin
        fsm_output = 10'b1001001010;
        state_var_NS = COMP_LOOP_C_449;
      end
      COMP_LOOP_C_449 : begin
        fsm_output = 10'b1001001011;
        state_var_NS = COMP_LOOP_C_450;
      end
      COMP_LOOP_C_450 : begin
        fsm_output = 10'b1001001100;
        if ( COMP_LOOP_C_450_tr0 ) begin
          state_var_NS = STAGE_VEC_LOOP_C_1;
        end
        else begin
          state_var_NS = COMP_LOOP_C_451;
        end
      end
      COMP_LOOP_C_451 : begin
        fsm_output = 10'b1001001101;
        state_var_NS = COMP_LOOP_C_452;
      end
      COMP_LOOP_C_452 : begin
        fsm_output = 10'b1001001110;
        state_var_NS = COMP_LOOP_C_453;
      end
      COMP_LOOP_C_453 : begin
        fsm_output = 10'b1001001111;
        state_var_NS = COMP_LOOP_C_454;
      end
      COMP_LOOP_C_454 : begin
        fsm_output = 10'b1001010000;
        state_var_NS = COMP_LOOP_C_455;
      end
      COMP_LOOP_C_455 : begin
        fsm_output = 10'b1001010001;
        state_var_NS = COMP_LOOP_C_456;
      end
      COMP_LOOP_C_456 : begin
        fsm_output = 10'b1001010010;
        state_var_NS = COMP_LOOP_C_457;
      end
      COMP_LOOP_C_457 : begin
        fsm_output = 10'b1001010011;
        state_var_NS = COMP_LOOP_C_458;
      end
      COMP_LOOP_C_458 : begin
        fsm_output = 10'b1001010100;
        state_var_NS = COMP_LOOP_C_459;
      end
      COMP_LOOP_C_459 : begin
        fsm_output = 10'b1001010101;
        state_var_NS = COMP_LOOP_C_460;
      end
      COMP_LOOP_C_460 : begin
        fsm_output = 10'b1001010110;
        state_var_NS = COMP_LOOP_C_461;
      end
      COMP_LOOP_C_461 : begin
        fsm_output = 10'b1001010111;
        state_var_NS = COMP_LOOP_C_462;
      end
      COMP_LOOP_C_462 : begin
        fsm_output = 10'b1001011000;
        state_var_NS = COMP_LOOP_C_463;
      end
      COMP_LOOP_C_463 : begin
        fsm_output = 10'b1001011001;
        state_var_NS = COMP_LOOP_C_464;
      end
      COMP_LOOP_C_464 : begin
        fsm_output = 10'b1001011010;
        state_var_NS = COMP_LOOP_C_465;
      end
      COMP_LOOP_C_465 : begin
        fsm_output = 10'b1001011011;
        state_var_NS = COMP_LOOP_C_466;
      end
      COMP_LOOP_C_466 : begin
        fsm_output = 10'b1001011100;
        state_var_NS = COMP_LOOP_11_modExp_dev_1_while_C_0;
      end
      COMP_LOOP_11_modExp_dev_1_while_C_0 : begin
        fsm_output = 10'b1001011101;
        state_var_NS = COMP_LOOP_11_modExp_dev_1_while_C_1;
      end
      COMP_LOOP_11_modExp_dev_1_while_C_1 : begin
        fsm_output = 10'b1001011110;
        state_var_NS = COMP_LOOP_11_modExp_dev_1_while_C_2;
      end
      COMP_LOOP_11_modExp_dev_1_while_C_2 : begin
        fsm_output = 10'b1001011111;
        state_var_NS = COMP_LOOP_11_modExp_dev_1_while_C_3;
      end
      COMP_LOOP_11_modExp_dev_1_while_C_3 : begin
        fsm_output = 10'b1001100000;
        state_var_NS = COMP_LOOP_11_modExp_dev_1_while_C_4;
      end
      COMP_LOOP_11_modExp_dev_1_while_C_4 : begin
        fsm_output = 10'b1001100001;
        state_var_NS = COMP_LOOP_11_modExp_dev_1_while_C_5;
      end
      COMP_LOOP_11_modExp_dev_1_while_C_5 : begin
        fsm_output = 10'b1001100010;
        state_var_NS = COMP_LOOP_11_modExp_dev_1_while_C_6;
      end
      COMP_LOOP_11_modExp_dev_1_while_C_6 : begin
        fsm_output = 10'b1001100011;
        state_var_NS = COMP_LOOP_11_modExp_dev_1_while_C_7;
      end
      COMP_LOOP_11_modExp_dev_1_while_C_7 : begin
        fsm_output = 10'b1001100100;
        state_var_NS = COMP_LOOP_11_modExp_dev_1_while_C_8;
      end
      COMP_LOOP_11_modExp_dev_1_while_C_8 : begin
        fsm_output = 10'b1001100101;
        state_var_NS = COMP_LOOP_11_modExp_dev_1_while_C_9;
      end
      COMP_LOOP_11_modExp_dev_1_while_C_9 : begin
        fsm_output = 10'b1001100110;
        state_var_NS = COMP_LOOP_11_modExp_dev_1_while_C_10;
      end
      COMP_LOOP_11_modExp_dev_1_while_C_10 : begin
        fsm_output = 10'b1001100111;
        state_var_NS = COMP_LOOP_11_modExp_dev_1_while_C_11;
      end
      COMP_LOOP_11_modExp_dev_1_while_C_11 : begin
        fsm_output = 10'b1001101000;
        if ( COMP_LOOP_11_modExp_dev_1_while_C_11_tr0 ) begin
          state_var_NS = COMP_LOOP_C_467;
        end
        else begin
          state_var_NS = COMP_LOOP_11_modExp_dev_1_while_C_0;
        end
      end
      COMP_LOOP_C_467 : begin
        fsm_output = 10'b1001101001;
        state_var_NS = COMP_LOOP_C_468;
      end
      COMP_LOOP_C_468 : begin
        fsm_output = 10'b1001101010;
        state_var_NS = COMP_LOOP_C_469;
      end
      COMP_LOOP_C_469 : begin
        fsm_output = 10'b1001101011;
        state_var_NS = COMP_LOOP_C_470;
      end
      COMP_LOOP_C_470 : begin
        fsm_output = 10'b1001101100;
        state_var_NS = COMP_LOOP_C_471;
      end
      COMP_LOOP_C_471 : begin
        fsm_output = 10'b1001101101;
        state_var_NS = COMP_LOOP_C_472;
      end
      COMP_LOOP_C_472 : begin
        fsm_output = 10'b1001101110;
        state_var_NS = COMP_LOOP_C_473;
      end
      COMP_LOOP_C_473 : begin
        fsm_output = 10'b1001101111;
        state_var_NS = COMP_LOOP_C_474;
      end
      COMP_LOOP_C_474 : begin
        fsm_output = 10'b1001110000;
        state_var_NS = COMP_LOOP_C_475;
      end
      COMP_LOOP_C_475 : begin
        fsm_output = 10'b1001110001;
        state_var_NS = COMP_LOOP_C_476;
      end
      COMP_LOOP_C_476 : begin
        fsm_output = 10'b1001110010;
        state_var_NS = COMP_LOOP_C_477;
      end
      COMP_LOOP_C_477 : begin
        fsm_output = 10'b1001110011;
        state_var_NS = COMP_LOOP_C_478;
      end
      COMP_LOOP_C_478 : begin
        fsm_output = 10'b1001110100;
        state_var_NS = COMP_LOOP_C_479;
      end
      COMP_LOOP_C_479 : begin
        fsm_output = 10'b1001110101;
        state_var_NS = COMP_LOOP_C_480;
      end
      COMP_LOOP_C_480 : begin
        fsm_output = 10'b1001110110;
        state_var_NS = COMP_LOOP_C_481;
      end
      COMP_LOOP_C_481 : begin
        fsm_output = 10'b1001110111;
        state_var_NS = COMP_LOOP_C_482;
      end
      COMP_LOOP_C_482 : begin
        fsm_output = 10'b1001111000;
        state_var_NS = COMP_LOOP_C_483;
      end
      COMP_LOOP_C_483 : begin
        fsm_output = 10'b1001111001;
        state_var_NS = COMP_LOOP_C_484;
      end
      COMP_LOOP_C_484 : begin
        fsm_output = 10'b1001111010;
        state_var_NS = COMP_LOOP_C_485;
      end
      COMP_LOOP_C_485 : begin
        fsm_output = 10'b1001111011;
        state_var_NS = COMP_LOOP_C_486;
      end
      COMP_LOOP_C_486 : begin
        fsm_output = 10'b1001111100;
        state_var_NS = COMP_LOOP_C_487;
      end
      COMP_LOOP_C_487 : begin
        fsm_output = 10'b1001111101;
        state_var_NS = COMP_LOOP_C_488;
      end
      COMP_LOOP_C_488 : begin
        fsm_output = 10'b1001111110;
        state_var_NS = COMP_LOOP_C_489;
      end
      COMP_LOOP_C_489 : begin
        fsm_output = 10'b1001111111;
        state_var_NS = COMP_LOOP_C_490;
      end
      COMP_LOOP_C_490 : begin
        fsm_output = 10'b1010000000;
        state_var_NS = COMP_LOOP_C_491;
      end
      COMP_LOOP_C_491 : begin
        fsm_output = 10'b1010000001;
        state_var_NS = COMP_LOOP_C_492;
      end
      COMP_LOOP_C_492 : begin
        fsm_output = 10'b1010000010;
        state_var_NS = COMP_LOOP_C_493;
      end
      COMP_LOOP_C_493 : begin
        fsm_output = 10'b1010000011;
        state_var_NS = COMP_LOOP_C_494;
      end
      COMP_LOOP_C_494 : begin
        fsm_output = 10'b1010000100;
        state_var_NS = COMP_LOOP_C_495;
      end
      COMP_LOOP_C_495 : begin
        fsm_output = 10'b1010000101;
        if ( COMP_LOOP_C_495_tr0 ) begin
          state_var_NS = STAGE_VEC_LOOP_C_1;
        end
        else begin
          state_var_NS = COMP_LOOP_C_496;
        end
      end
      COMP_LOOP_C_496 : begin
        fsm_output = 10'b1010000110;
        state_var_NS = COMP_LOOP_C_497;
      end
      COMP_LOOP_C_497 : begin
        fsm_output = 10'b1010000111;
        state_var_NS = COMP_LOOP_C_498;
      end
      COMP_LOOP_C_498 : begin
        fsm_output = 10'b1010001000;
        state_var_NS = COMP_LOOP_C_499;
      end
      COMP_LOOP_C_499 : begin
        fsm_output = 10'b1010001001;
        state_var_NS = COMP_LOOP_C_500;
      end
      COMP_LOOP_C_500 : begin
        fsm_output = 10'b1010001010;
        state_var_NS = COMP_LOOP_C_501;
      end
      COMP_LOOP_C_501 : begin
        fsm_output = 10'b1010001011;
        state_var_NS = COMP_LOOP_C_502;
      end
      COMP_LOOP_C_502 : begin
        fsm_output = 10'b1010001100;
        state_var_NS = COMP_LOOP_C_503;
      end
      COMP_LOOP_C_503 : begin
        fsm_output = 10'b1010001101;
        state_var_NS = COMP_LOOP_C_504;
      end
      COMP_LOOP_C_504 : begin
        fsm_output = 10'b1010001110;
        state_var_NS = COMP_LOOP_C_505;
      end
      COMP_LOOP_C_505 : begin
        fsm_output = 10'b1010001111;
        state_var_NS = COMP_LOOP_C_506;
      end
      COMP_LOOP_C_506 : begin
        fsm_output = 10'b1010010000;
        state_var_NS = COMP_LOOP_C_507;
      end
      COMP_LOOP_C_507 : begin
        fsm_output = 10'b1010010001;
        state_var_NS = COMP_LOOP_C_508;
      end
      COMP_LOOP_C_508 : begin
        fsm_output = 10'b1010010010;
        state_var_NS = COMP_LOOP_C_509;
      end
      COMP_LOOP_C_509 : begin
        fsm_output = 10'b1010010011;
        state_var_NS = COMP_LOOP_C_510;
      end
      COMP_LOOP_C_510 : begin
        fsm_output = 10'b1010010100;
        state_var_NS = COMP_LOOP_C_511;
      end
      COMP_LOOP_C_511 : begin
        fsm_output = 10'b1010010101;
        state_var_NS = COMP_LOOP_12_modExp_dev_1_while_C_0;
      end
      COMP_LOOP_12_modExp_dev_1_while_C_0 : begin
        fsm_output = 10'b1010010110;
        state_var_NS = COMP_LOOP_12_modExp_dev_1_while_C_1;
      end
      COMP_LOOP_12_modExp_dev_1_while_C_1 : begin
        fsm_output = 10'b1010010111;
        state_var_NS = COMP_LOOP_12_modExp_dev_1_while_C_2;
      end
      COMP_LOOP_12_modExp_dev_1_while_C_2 : begin
        fsm_output = 10'b1010011000;
        state_var_NS = COMP_LOOP_12_modExp_dev_1_while_C_3;
      end
      COMP_LOOP_12_modExp_dev_1_while_C_3 : begin
        fsm_output = 10'b1010011001;
        state_var_NS = COMP_LOOP_12_modExp_dev_1_while_C_4;
      end
      COMP_LOOP_12_modExp_dev_1_while_C_4 : begin
        fsm_output = 10'b1010011010;
        state_var_NS = COMP_LOOP_12_modExp_dev_1_while_C_5;
      end
      COMP_LOOP_12_modExp_dev_1_while_C_5 : begin
        fsm_output = 10'b1010011011;
        state_var_NS = COMP_LOOP_12_modExp_dev_1_while_C_6;
      end
      COMP_LOOP_12_modExp_dev_1_while_C_6 : begin
        fsm_output = 10'b1010011100;
        state_var_NS = COMP_LOOP_12_modExp_dev_1_while_C_7;
      end
      COMP_LOOP_12_modExp_dev_1_while_C_7 : begin
        fsm_output = 10'b1010011101;
        state_var_NS = COMP_LOOP_12_modExp_dev_1_while_C_8;
      end
      COMP_LOOP_12_modExp_dev_1_while_C_8 : begin
        fsm_output = 10'b1010011110;
        state_var_NS = COMP_LOOP_12_modExp_dev_1_while_C_9;
      end
      COMP_LOOP_12_modExp_dev_1_while_C_9 : begin
        fsm_output = 10'b1010011111;
        state_var_NS = COMP_LOOP_12_modExp_dev_1_while_C_10;
      end
      COMP_LOOP_12_modExp_dev_1_while_C_10 : begin
        fsm_output = 10'b1010100000;
        state_var_NS = COMP_LOOP_12_modExp_dev_1_while_C_11;
      end
      COMP_LOOP_12_modExp_dev_1_while_C_11 : begin
        fsm_output = 10'b1010100001;
        if ( COMP_LOOP_12_modExp_dev_1_while_C_11_tr0 ) begin
          state_var_NS = COMP_LOOP_C_512;
        end
        else begin
          state_var_NS = COMP_LOOP_12_modExp_dev_1_while_C_0;
        end
      end
      COMP_LOOP_C_512 : begin
        fsm_output = 10'b1010100010;
        state_var_NS = COMP_LOOP_C_513;
      end
      COMP_LOOP_C_513 : begin
        fsm_output = 10'b1010100011;
        state_var_NS = COMP_LOOP_C_514;
      end
      COMP_LOOP_C_514 : begin
        fsm_output = 10'b1010100100;
        state_var_NS = COMP_LOOP_C_515;
      end
      COMP_LOOP_C_515 : begin
        fsm_output = 10'b1010100101;
        state_var_NS = COMP_LOOP_C_516;
      end
      COMP_LOOP_C_516 : begin
        fsm_output = 10'b1010100110;
        state_var_NS = COMP_LOOP_C_517;
      end
      COMP_LOOP_C_517 : begin
        fsm_output = 10'b1010100111;
        state_var_NS = COMP_LOOP_C_518;
      end
      COMP_LOOP_C_518 : begin
        fsm_output = 10'b1010101000;
        state_var_NS = COMP_LOOP_C_519;
      end
      COMP_LOOP_C_519 : begin
        fsm_output = 10'b1010101001;
        state_var_NS = COMP_LOOP_C_520;
      end
      COMP_LOOP_C_520 : begin
        fsm_output = 10'b1010101010;
        state_var_NS = COMP_LOOP_C_521;
      end
      COMP_LOOP_C_521 : begin
        fsm_output = 10'b1010101011;
        state_var_NS = COMP_LOOP_C_522;
      end
      COMP_LOOP_C_522 : begin
        fsm_output = 10'b1010101100;
        state_var_NS = COMP_LOOP_C_523;
      end
      COMP_LOOP_C_523 : begin
        fsm_output = 10'b1010101101;
        state_var_NS = COMP_LOOP_C_524;
      end
      COMP_LOOP_C_524 : begin
        fsm_output = 10'b1010101110;
        state_var_NS = COMP_LOOP_C_525;
      end
      COMP_LOOP_C_525 : begin
        fsm_output = 10'b1010101111;
        state_var_NS = COMP_LOOP_C_526;
      end
      COMP_LOOP_C_526 : begin
        fsm_output = 10'b1010110000;
        state_var_NS = COMP_LOOP_C_527;
      end
      COMP_LOOP_C_527 : begin
        fsm_output = 10'b1010110001;
        state_var_NS = COMP_LOOP_C_528;
      end
      COMP_LOOP_C_528 : begin
        fsm_output = 10'b1010110010;
        state_var_NS = COMP_LOOP_C_529;
      end
      COMP_LOOP_C_529 : begin
        fsm_output = 10'b1010110011;
        state_var_NS = COMP_LOOP_C_530;
      end
      COMP_LOOP_C_530 : begin
        fsm_output = 10'b1010110100;
        state_var_NS = COMP_LOOP_C_531;
      end
      COMP_LOOP_C_531 : begin
        fsm_output = 10'b1010110101;
        state_var_NS = COMP_LOOP_C_532;
      end
      COMP_LOOP_C_532 : begin
        fsm_output = 10'b1010110110;
        state_var_NS = COMP_LOOP_C_533;
      end
      COMP_LOOP_C_533 : begin
        fsm_output = 10'b1010110111;
        state_var_NS = COMP_LOOP_C_534;
      end
      COMP_LOOP_C_534 : begin
        fsm_output = 10'b1010111000;
        state_var_NS = COMP_LOOP_C_535;
      end
      COMP_LOOP_C_535 : begin
        fsm_output = 10'b1010111001;
        state_var_NS = COMP_LOOP_C_536;
      end
      COMP_LOOP_C_536 : begin
        fsm_output = 10'b1010111010;
        state_var_NS = COMP_LOOP_C_537;
      end
      COMP_LOOP_C_537 : begin
        fsm_output = 10'b1010111011;
        state_var_NS = COMP_LOOP_C_538;
      end
      COMP_LOOP_C_538 : begin
        fsm_output = 10'b1010111100;
        state_var_NS = COMP_LOOP_C_539;
      end
      COMP_LOOP_C_539 : begin
        fsm_output = 10'b1010111101;
        state_var_NS = COMP_LOOP_C_540;
      end
      COMP_LOOP_C_540 : begin
        fsm_output = 10'b1010111110;
        if ( COMP_LOOP_C_540_tr0 ) begin
          state_var_NS = STAGE_VEC_LOOP_C_1;
        end
        else begin
          state_var_NS = COMP_LOOP_C_541;
        end
      end
      COMP_LOOP_C_541 : begin
        fsm_output = 10'b1010111111;
        state_var_NS = COMP_LOOP_C_542;
      end
      COMP_LOOP_C_542 : begin
        fsm_output = 10'b1011000000;
        state_var_NS = COMP_LOOP_C_543;
      end
      COMP_LOOP_C_543 : begin
        fsm_output = 10'b1011000001;
        state_var_NS = COMP_LOOP_C_544;
      end
      COMP_LOOP_C_544 : begin
        fsm_output = 10'b1011000010;
        state_var_NS = COMP_LOOP_C_545;
      end
      COMP_LOOP_C_545 : begin
        fsm_output = 10'b1011000011;
        state_var_NS = COMP_LOOP_C_546;
      end
      COMP_LOOP_C_546 : begin
        fsm_output = 10'b1011000100;
        state_var_NS = COMP_LOOP_C_547;
      end
      COMP_LOOP_C_547 : begin
        fsm_output = 10'b1011000101;
        state_var_NS = COMP_LOOP_C_548;
      end
      COMP_LOOP_C_548 : begin
        fsm_output = 10'b1011000110;
        state_var_NS = COMP_LOOP_C_549;
      end
      COMP_LOOP_C_549 : begin
        fsm_output = 10'b1011000111;
        state_var_NS = COMP_LOOP_C_550;
      end
      COMP_LOOP_C_550 : begin
        fsm_output = 10'b1011001000;
        state_var_NS = COMP_LOOP_C_551;
      end
      COMP_LOOP_C_551 : begin
        fsm_output = 10'b1011001001;
        state_var_NS = COMP_LOOP_C_552;
      end
      COMP_LOOP_C_552 : begin
        fsm_output = 10'b1011001010;
        state_var_NS = COMP_LOOP_C_553;
      end
      COMP_LOOP_C_553 : begin
        fsm_output = 10'b1011001011;
        state_var_NS = COMP_LOOP_C_554;
      end
      COMP_LOOP_C_554 : begin
        fsm_output = 10'b1011001100;
        state_var_NS = COMP_LOOP_C_555;
      end
      COMP_LOOP_C_555 : begin
        fsm_output = 10'b1011001101;
        state_var_NS = COMP_LOOP_C_556;
      end
      COMP_LOOP_C_556 : begin
        fsm_output = 10'b1011001110;
        state_var_NS = COMP_LOOP_13_modExp_dev_1_while_C_0;
      end
      COMP_LOOP_13_modExp_dev_1_while_C_0 : begin
        fsm_output = 10'b1011001111;
        state_var_NS = COMP_LOOP_13_modExp_dev_1_while_C_1;
      end
      COMP_LOOP_13_modExp_dev_1_while_C_1 : begin
        fsm_output = 10'b1011010000;
        state_var_NS = COMP_LOOP_13_modExp_dev_1_while_C_2;
      end
      COMP_LOOP_13_modExp_dev_1_while_C_2 : begin
        fsm_output = 10'b1011010001;
        state_var_NS = COMP_LOOP_13_modExp_dev_1_while_C_3;
      end
      COMP_LOOP_13_modExp_dev_1_while_C_3 : begin
        fsm_output = 10'b1011010010;
        state_var_NS = COMP_LOOP_13_modExp_dev_1_while_C_4;
      end
      COMP_LOOP_13_modExp_dev_1_while_C_4 : begin
        fsm_output = 10'b1011010011;
        state_var_NS = COMP_LOOP_13_modExp_dev_1_while_C_5;
      end
      COMP_LOOP_13_modExp_dev_1_while_C_5 : begin
        fsm_output = 10'b1011010100;
        state_var_NS = COMP_LOOP_13_modExp_dev_1_while_C_6;
      end
      COMP_LOOP_13_modExp_dev_1_while_C_6 : begin
        fsm_output = 10'b1011010101;
        state_var_NS = COMP_LOOP_13_modExp_dev_1_while_C_7;
      end
      COMP_LOOP_13_modExp_dev_1_while_C_7 : begin
        fsm_output = 10'b1011010110;
        state_var_NS = COMP_LOOP_13_modExp_dev_1_while_C_8;
      end
      COMP_LOOP_13_modExp_dev_1_while_C_8 : begin
        fsm_output = 10'b1011010111;
        state_var_NS = COMP_LOOP_13_modExp_dev_1_while_C_9;
      end
      COMP_LOOP_13_modExp_dev_1_while_C_9 : begin
        fsm_output = 10'b1011011000;
        state_var_NS = COMP_LOOP_13_modExp_dev_1_while_C_10;
      end
      COMP_LOOP_13_modExp_dev_1_while_C_10 : begin
        fsm_output = 10'b1011011001;
        state_var_NS = COMP_LOOP_13_modExp_dev_1_while_C_11;
      end
      COMP_LOOP_13_modExp_dev_1_while_C_11 : begin
        fsm_output = 10'b1011011010;
        if ( COMP_LOOP_13_modExp_dev_1_while_C_11_tr0 ) begin
          state_var_NS = COMP_LOOP_C_557;
        end
        else begin
          state_var_NS = COMP_LOOP_13_modExp_dev_1_while_C_0;
        end
      end
      COMP_LOOP_C_557 : begin
        fsm_output = 10'b1011011011;
        state_var_NS = COMP_LOOP_C_558;
      end
      COMP_LOOP_C_558 : begin
        fsm_output = 10'b1011011100;
        state_var_NS = COMP_LOOP_C_559;
      end
      COMP_LOOP_C_559 : begin
        fsm_output = 10'b1011011101;
        state_var_NS = COMP_LOOP_C_560;
      end
      COMP_LOOP_C_560 : begin
        fsm_output = 10'b1011011110;
        state_var_NS = COMP_LOOP_C_561;
      end
      COMP_LOOP_C_561 : begin
        fsm_output = 10'b1011011111;
        state_var_NS = COMP_LOOP_C_562;
      end
      COMP_LOOP_C_562 : begin
        fsm_output = 10'b1011100000;
        state_var_NS = COMP_LOOP_C_563;
      end
      COMP_LOOP_C_563 : begin
        fsm_output = 10'b1011100001;
        state_var_NS = COMP_LOOP_C_564;
      end
      COMP_LOOP_C_564 : begin
        fsm_output = 10'b1011100010;
        state_var_NS = COMP_LOOP_C_565;
      end
      COMP_LOOP_C_565 : begin
        fsm_output = 10'b1011100011;
        state_var_NS = COMP_LOOP_C_566;
      end
      COMP_LOOP_C_566 : begin
        fsm_output = 10'b1011100100;
        state_var_NS = COMP_LOOP_C_567;
      end
      COMP_LOOP_C_567 : begin
        fsm_output = 10'b1011100101;
        state_var_NS = COMP_LOOP_C_568;
      end
      COMP_LOOP_C_568 : begin
        fsm_output = 10'b1011100110;
        state_var_NS = COMP_LOOP_C_569;
      end
      COMP_LOOP_C_569 : begin
        fsm_output = 10'b1011100111;
        state_var_NS = COMP_LOOP_C_570;
      end
      COMP_LOOP_C_570 : begin
        fsm_output = 10'b1011101000;
        state_var_NS = COMP_LOOP_C_571;
      end
      COMP_LOOP_C_571 : begin
        fsm_output = 10'b1011101001;
        state_var_NS = COMP_LOOP_C_572;
      end
      COMP_LOOP_C_572 : begin
        fsm_output = 10'b1011101010;
        state_var_NS = COMP_LOOP_C_573;
      end
      COMP_LOOP_C_573 : begin
        fsm_output = 10'b1011101011;
        state_var_NS = COMP_LOOP_C_574;
      end
      COMP_LOOP_C_574 : begin
        fsm_output = 10'b1011101100;
        state_var_NS = COMP_LOOP_C_575;
      end
      COMP_LOOP_C_575 : begin
        fsm_output = 10'b1011101101;
        state_var_NS = COMP_LOOP_C_576;
      end
      COMP_LOOP_C_576 : begin
        fsm_output = 10'b1011101110;
        state_var_NS = COMP_LOOP_C_577;
      end
      COMP_LOOP_C_577 : begin
        fsm_output = 10'b1011101111;
        state_var_NS = COMP_LOOP_C_578;
      end
      COMP_LOOP_C_578 : begin
        fsm_output = 10'b1011110000;
        state_var_NS = COMP_LOOP_C_579;
      end
      COMP_LOOP_C_579 : begin
        fsm_output = 10'b1011110001;
        state_var_NS = COMP_LOOP_C_580;
      end
      COMP_LOOP_C_580 : begin
        fsm_output = 10'b1011110010;
        state_var_NS = COMP_LOOP_C_581;
      end
      COMP_LOOP_C_581 : begin
        fsm_output = 10'b1011110011;
        state_var_NS = COMP_LOOP_C_582;
      end
      COMP_LOOP_C_582 : begin
        fsm_output = 10'b1011110100;
        state_var_NS = COMP_LOOP_C_583;
      end
      COMP_LOOP_C_583 : begin
        fsm_output = 10'b1011110101;
        state_var_NS = COMP_LOOP_C_584;
      end
      COMP_LOOP_C_584 : begin
        fsm_output = 10'b1011110110;
        state_var_NS = COMP_LOOP_C_585;
      end
      COMP_LOOP_C_585 : begin
        fsm_output = 10'b1011110111;
        if ( COMP_LOOP_C_585_tr0 ) begin
          state_var_NS = STAGE_VEC_LOOP_C_1;
        end
        else begin
          state_var_NS = COMP_LOOP_C_586;
        end
      end
      COMP_LOOP_C_586 : begin
        fsm_output = 10'b1011111000;
        state_var_NS = COMP_LOOP_C_587;
      end
      COMP_LOOP_C_587 : begin
        fsm_output = 10'b1011111001;
        state_var_NS = COMP_LOOP_C_588;
      end
      COMP_LOOP_C_588 : begin
        fsm_output = 10'b1011111010;
        state_var_NS = COMP_LOOP_C_589;
      end
      COMP_LOOP_C_589 : begin
        fsm_output = 10'b1011111011;
        state_var_NS = COMP_LOOP_C_590;
      end
      COMP_LOOP_C_590 : begin
        fsm_output = 10'b1011111100;
        state_var_NS = COMP_LOOP_C_591;
      end
      COMP_LOOP_C_591 : begin
        fsm_output = 10'b1011111101;
        state_var_NS = COMP_LOOP_C_592;
      end
      COMP_LOOP_C_592 : begin
        fsm_output = 10'b1011111110;
        state_var_NS = COMP_LOOP_C_593;
      end
      COMP_LOOP_C_593 : begin
        fsm_output = 10'b1011111111;
        state_var_NS = COMP_LOOP_C_594;
      end
      COMP_LOOP_C_594 : begin
        fsm_output = 10'b1100000000;
        state_var_NS = COMP_LOOP_C_595;
      end
      COMP_LOOP_C_595 : begin
        fsm_output = 10'b1100000001;
        state_var_NS = COMP_LOOP_C_596;
      end
      COMP_LOOP_C_596 : begin
        fsm_output = 10'b1100000010;
        state_var_NS = COMP_LOOP_C_597;
      end
      COMP_LOOP_C_597 : begin
        fsm_output = 10'b1100000011;
        state_var_NS = COMP_LOOP_C_598;
      end
      COMP_LOOP_C_598 : begin
        fsm_output = 10'b1100000100;
        state_var_NS = COMP_LOOP_C_599;
      end
      COMP_LOOP_C_599 : begin
        fsm_output = 10'b1100000101;
        state_var_NS = COMP_LOOP_C_600;
      end
      COMP_LOOP_C_600 : begin
        fsm_output = 10'b1100000110;
        state_var_NS = COMP_LOOP_C_601;
      end
      COMP_LOOP_C_601 : begin
        fsm_output = 10'b1100000111;
        state_var_NS = COMP_LOOP_14_modExp_dev_1_while_C_0;
      end
      COMP_LOOP_14_modExp_dev_1_while_C_0 : begin
        fsm_output = 10'b1100001000;
        state_var_NS = COMP_LOOP_14_modExp_dev_1_while_C_1;
      end
      COMP_LOOP_14_modExp_dev_1_while_C_1 : begin
        fsm_output = 10'b1100001001;
        state_var_NS = COMP_LOOP_14_modExp_dev_1_while_C_2;
      end
      COMP_LOOP_14_modExp_dev_1_while_C_2 : begin
        fsm_output = 10'b1100001010;
        state_var_NS = COMP_LOOP_14_modExp_dev_1_while_C_3;
      end
      COMP_LOOP_14_modExp_dev_1_while_C_3 : begin
        fsm_output = 10'b1100001011;
        state_var_NS = COMP_LOOP_14_modExp_dev_1_while_C_4;
      end
      COMP_LOOP_14_modExp_dev_1_while_C_4 : begin
        fsm_output = 10'b1100001100;
        state_var_NS = COMP_LOOP_14_modExp_dev_1_while_C_5;
      end
      COMP_LOOP_14_modExp_dev_1_while_C_5 : begin
        fsm_output = 10'b1100001101;
        state_var_NS = COMP_LOOP_14_modExp_dev_1_while_C_6;
      end
      COMP_LOOP_14_modExp_dev_1_while_C_6 : begin
        fsm_output = 10'b1100001110;
        state_var_NS = COMP_LOOP_14_modExp_dev_1_while_C_7;
      end
      COMP_LOOP_14_modExp_dev_1_while_C_7 : begin
        fsm_output = 10'b1100001111;
        state_var_NS = COMP_LOOP_14_modExp_dev_1_while_C_8;
      end
      COMP_LOOP_14_modExp_dev_1_while_C_8 : begin
        fsm_output = 10'b1100010000;
        state_var_NS = COMP_LOOP_14_modExp_dev_1_while_C_9;
      end
      COMP_LOOP_14_modExp_dev_1_while_C_9 : begin
        fsm_output = 10'b1100010001;
        state_var_NS = COMP_LOOP_14_modExp_dev_1_while_C_10;
      end
      COMP_LOOP_14_modExp_dev_1_while_C_10 : begin
        fsm_output = 10'b1100010010;
        state_var_NS = COMP_LOOP_14_modExp_dev_1_while_C_11;
      end
      COMP_LOOP_14_modExp_dev_1_while_C_11 : begin
        fsm_output = 10'b1100010011;
        if ( COMP_LOOP_14_modExp_dev_1_while_C_11_tr0 ) begin
          state_var_NS = COMP_LOOP_C_602;
        end
        else begin
          state_var_NS = COMP_LOOP_14_modExp_dev_1_while_C_0;
        end
      end
      COMP_LOOP_C_602 : begin
        fsm_output = 10'b1100010100;
        state_var_NS = COMP_LOOP_C_603;
      end
      COMP_LOOP_C_603 : begin
        fsm_output = 10'b1100010101;
        state_var_NS = COMP_LOOP_C_604;
      end
      COMP_LOOP_C_604 : begin
        fsm_output = 10'b1100010110;
        state_var_NS = COMP_LOOP_C_605;
      end
      COMP_LOOP_C_605 : begin
        fsm_output = 10'b1100010111;
        state_var_NS = COMP_LOOP_C_606;
      end
      COMP_LOOP_C_606 : begin
        fsm_output = 10'b1100011000;
        state_var_NS = COMP_LOOP_C_607;
      end
      COMP_LOOP_C_607 : begin
        fsm_output = 10'b1100011001;
        state_var_NS = COMP_LOOP_C_608;
      end
      COMP_LOOP_C_608 : begin
        fsm_output = 10'b1100011010;
        state_var_NS = COMP_LOOP_C_609;
      end
      COMP_LOOP_C_609 : begin
        fsm_output = 10'b1100011011;
        state_var_NS = COMP_LOOP_C_610;
      end
      COMP_LOOP_C_610 : begin
        fsm_output = 10'b1100011100;
        state_var_NS = COMP_LOOP_C_611;
      end
      COMP_LOOP_C_611 : begin
        fsm_output = 10'b1100011101;
        state_var_NS = COMP_LOOP_C_612;
      end
      COMP_LOOP_C_612 : begin
        fsm_output = 10'b1100011110;
        state_var_NS = COMP_LOOP_C_613;
      end
      COMP_LOOP_C_613 : begin
        fsm_output = 10'b1100011111;
        state_var_NS = COMP_LOOP_C_614;
      end
      COMP_LOOP_C_614 : begin
        fsm_output = 10'b1100100000;
        state_var_NS = COMP_LOOP_C_615;
      end
      COMP_LOOP_C_615 : begin
        fsm_output = 10'b1100100001;
        state_var_NS = COMP_LOOP_C_616;
      end
      COMP_LOOP_C_616 : begin
        fsm_output = 10'b1100100010;
        state_var_NS = COMP_LOOP_C_617;
      end
      COMP_LOOP_C_617 : begin
        fsm_output = 10'b1100100011;
        state_var_NS = COMP_LOOP_C_618;
      end
      COMP_LOOP_C_618 : begin
        fsm_output = 10'b1100100100;
        state_var_NS = COMP_LOOP_C_619;
      end
      COMP_LOOP_C_619 : begin
        fsm_output = 10'b1100100101;
        state_var_NS = COMP_LOOP_C_620;
      end
      COMP_LOOP_C_620 : begin
        fsm_output = 10'b1100100110;
        state_var_NS = COMP_LOOP_C_621;
      end
      COMP_LOOP_C_621 : begin
        fsm_output = 10'b1100100111;
        state_var_NS = COMP_LOOP_C_622;
      end
      COMP_LOOP_C_622 : begin
        fsm_output = 10'b1100101000;
        state_var_NS = COMP_LOOP_C_623;
      end
      COMP_LOOP_C_623 : begin
        fsm_output = 10'b1100101001;
        state_var_NS = COMP_LOOP_C_624;
      end
      COMP_LOOP_C_624 : begin
        fsm_output = 10'b1100101010;
        state_var_NS = COMP_LOOP_C_625;
      end
      COMP_LOOP_C_625 : begin
        fsm_output = 10'b1100101011;
        state_var_NS = COMP_LOOP_C_626;
      end
      COMP_LOOP_C_626 : begin
        fsm_output = 10'b1100101100;
        state_var_NS = COMP_LOOP_C_627;
      end
      COMP_LOOP_C_627 : begin
        fsm_output = 10'b1100101101;
        state_var_NS = COMP_LOOP_C_628;
      end
      COMP_LOOP_C_628 : begin
        fsm_output = 10'b1100101110;
        state_var_NS = COMP_LOOP_C_629;
      end
      COMP_LOOP_C_629 : begin
        fsm_output = 10'b1100101111;
        state_var_NS = COMP_LOOP_C_630;
      end
      COMP_LOOP_C_630 : begin
        fsm_output = 10'b1100110000;
        if ( COMP_LOOP_C_630_tr0 ) begin
          state_var_NS = STAGE_VEC_LOOP_C_1;
        end
        else begin
          state_var_NS = COMP_LOOP_C_631;
        end
      end
      COMP_LOOP_C_631 : begin
        fsm_output = 10'b1100110001;
        state_var_NS = COMP_LOOP_C_632;
      end
      COMP_LOOP_C_632 : begin
        fsm_output = 10'b1100110010;
        state_var_NS = COMP_LOOP_C_633;
      end
      COMP_LOOP_C_633 : begin
        fsm_output = 10'b1100110011;
        state_var_NS = COMP_LOOP_C_634;
      end
      COMP_LOOP_C_634 : begin
        fsm_output = 10'b1100110100;
        state_var_NS = COMP_LOOP_C_635;
      end
      COMP_LOOP_C_635 : begin
        fsm_output = 10'b1100110101;
        state_var_NS = COMP_LOOP_C_636;
      end
      COMP_LOOP_C_636 : begin
        fsm_output = 10'b1100110110;
        state_var_NS = COMP_LOOP_C_637;
      end
      COMP_LOOP_C_637 : begin
        fsm_output = 10'b1100110111;
        state_var_NS = COMP_LOOP_C_638;
      end
      COMP_LOOP_C_638 : begin
        fsm_output = 10'b1100111000;
        state_var_NS = COMP_LOOP_C_639;
      end
      COMP_LOOP_C_639 : begin
        fsm_output = 10'b1100111001;
        state_var_NS = COMP_LOOP_C_640;
      end
      COMP_LOOP_C_640 : begin
        fsm_output = 10'b1100111010;
        state_var_NS = COMP_LOOP_C_641;
      end
      COMP_LOOP_C_641 : begin
        fsm_output = 10'b1100111011;
        state_var_NS = COMP_LOOP_C_642;
      end
      COMP_LOOP_C_642 : begin
        fsm_output = 10'b1100111100;
        state_var_NS = COMP_LOOP_C_643;
      end
      COMP_LOOP_C_643 : begin
        fsm_output = 10'b1100111101;
        state_var_NS = COMP_LOOP_C_644;
      end
      COMP_LOOP_C_644 : begin
        fsm_output = 10'b1100111110;
        state_var_NS = COMP_LOOP_C_645;
      end
      COMP_LOOP_C_645 : begin
        fsm_output = 10'b1100111111;
        state_var_NS = COMP_LOOP_C_646;
      end
      COMP_LOOP_C_646 : begin
        fsm_output = 10'b1101000000;
        state_var_NS = COMP_LOOP_15_modExp_dev_1_while_C_0;
      end
      COMP_LOOP_15_modExp_dev_1_while_C_0 : begin
        fsm_output = 10'b1101000001;
        state_var_NS = COMP_LOOP_15_modExp_dev_1_while_C_1;
      end
      COMP_LOOP_15_modExp_dev_1_while_C_1 : begin
        fsm_output = 10'b1101000010;
        state_var_NS = COMP_LOOP_15_modExp_dev_1_while_C_2;
      end
      COMP_LOOP_15_modExp_dev_1_while_C_2 : begin
        fsm_output = 10'b1101000011;
        state_var_NS = COMP_LOOP_15_modExp_dev_1_while_C_3;
      end
      COMP_LOOP_15_modExp_dev_1_while_C_3 : begin
        fsm_output = 10'b1101000100;
        state_var_NS = COMP_LOOP_15_modExp_dev_1_while_C_4;
      end
      COMP_LOOP_15_modExp_dev_1_while_C_4 : begin
        fsm_output = 10'b1101000101;
        state_var_NS = COMP_LOOP_15_modExp_dev_1_while_C_5;
      end
      COMP_LOOP_15_modExp_dev_1_while_C_5 : begin
        fsm_output = 10'b1101000110;
        state_var_NS = COMP_LOOP_15_modExp_dev_1_while_C_6;
      end
      COMP_LOOP_15_modExp_dev_1_while_C_6 : begin
        fsm_output = 10'b1101000111;
        state_var_NS = COMP_LOOP_15_modExp_dev_1_while_C_7;
      end
      COMP_LOOP_15_modExp_dev_1_while_C_7 : begin
        fsm_output = 10'b1101001000;
        state_var_NS = COMP_LOOP_15_modExp_dev_1_while_C_8;
      end
      COMP_LOOP_15_modExp_dev_1_while_C_8 : begin
        fsm_output = 10'b1101001001;
        state_var_NS = COMP_LOOP_15_modExp_dev_1_while_C_9;
      end
      COMP_LOOP_15_modExp_dev_1_while_C_9 : begin
        fsm_output = 10'b1101001010;
        state_var_NS = COMP_LOOP_15_modExp_dev_1_while_C_10;
      end
      COMP_LOOP_15_modExp_dev_1_while_C_10 : begin
        fsm_output = 10'b1101001011;
        state_var_NS = COMP_LOOP_15_modExp_dev_1_while_C_11;
      end
      COMP_LOOP_15_modExp_dev_1_while_C_11 : begin
        fsm_output = 10'b1101001100;
        if ( COMP_LOOP_15_modExp_dev_1_while_C_11_tr0 ) begin
          state_var_NS = COMP_LOOP_C_647;
        end
        else begin
          state_var_NS = COMP_LOOP_15_modExp_dev_1_while_C_0;
        end
      end
      COMP_LOOP_C_647 : begin
        fsm_output = 10'b1101001101;
        state_var_NS = COMP_LOOP_C_648;
      end
      COMP_LOOP_C_648 : begin
        fsm_output = 10'b1101001110;
        state_var_NS = COMP_LOOP_C_649;
      end
      COMP_LOOP_C_649 : begin
        fsm_output = 10'b1101001111;
        state_var_NS = COMP_LOOP_C_650;
      end
      COMP_LOOP_C_650 : begin
        fsm_output = 10'b1101010000;
        state_var_NS = COMP_LOOP_C_651;
      end
      COMP_LOOP_C_651 : begin
        fsm_output = 10'b1101010001;
        state_var_NS = COMP_LOOP_C_652;
      end
      COMP_LOOP_C_652 : begin
        fsm_output = 10'b1101010010;
        state_var_NS = COMP_LOOP_C_653;
      end
      COMP_LOOP_C_653 : begin
        fsm_output = 10'b1101010011;
        state_var_NS = COMP_LOOP_C_654;
      end
      COMP_LOOP_C_654 : begin
        fsm_output = 10'b1101010100;
        state_var_NS = COMP_LOOP_C_655;
      end
      COMP_LOOP_C_655 : begin
        fsm_output = 10'b1101010101;
        state_var_NS = COMP_LOOP_C_656;
      end
      COMP_LOOP_C_656 : begin
        fsm_output = 10'b1101010110;
        state_var_NS = COMP_LOOP_C_657;
      end
      COMP_LOOP_C_657 : begin
        fsm_output = 10'b1101010111;
        state_var_NS = COMP_LOOP_C_658;
      end
      COMP_LOOP_C_658 : begin
        fsm_output = 10'b1101011000;
        state_var_NS = COMP_LOOP_C_659;
      end
      COMP_LOOP_C_659 : begin
        fsm_output = 10'b1101011001;
        state_var_NS = COMP_LOOP_C_660;
      end
      COMP_LOOP_C_660 : begin
        fsm_output = 10'b1101011010;
        state_var_NS = COMP_LOOP_C_661;
      end
      COMP_LOOP_C_661 : begin
        fsm_output = 10'b1101011011;
        state_var_NS = COMP_LOOP_C_662;
      end
      COMP_LOOP_C_662 : begin
        fsm_output = 10'b1101011100;
        state_var_NS = COMP_LOOP_C_663;
      end
      COMP_LOOP_C_663 : begin
        fsm_output = 10'b1101011101;
        state_var_NS = COMP_LOOP_C_664;
      end
      COMP_LOOP_C_664 : begin
        fsm_output = 10'b1101011110;
        state_var_NS = COMP_LOOP_C_665;
      end
      COMP_LOOP_C_665 : begin
        fsm_output = 10'b1101011111;
        state_var_NS = COMP_LOOP_C_666;
      end
      COMP_LOOP_C_666 : begin
        fsm_output = 10'b1101100000;
        state_var_NS = COMP_LOOP_C_667;
      end
      COMP_LOOP_C_667 : begin
        fsm_output = 10'b1101100001;
        state_var_NS = COMP_LOOP_C_668;
      end
      COMP_LOOP_C_668 : begin
        fsm_output = 10'b1101100010;
        state_var_NS = COMP_LOOP_C_669;
      end
      COMP_LOOP_C_669 : begin
        fsm_output = 10'b1101100011;
        state_var_NS = COMP_LOOP_C_670;
      end
      COMP_LOOP_C_670 : begin
        fsm_output = 10'b1101100100;
        state_var_NS = COMP_LOOP_C_671;
      end
      COMP_LOOP_C_671 : begin
        fsm_output = 10'b1101100101;
        state_var_NS = COMP_LOOP_C_672;
      end
      COMP_LOOP_C_672 : begin
        fsm_output = 10'b1101100110;
        state_var_NS = COMP_LOOP_C_673;
      end
      COMP_LOOP_C_673 : begin
        fsm_output = 10'b1101100111;
        state_var_NS = COMP_LOOP_C_674;
      end
      COMP_LOOP_C_674 : begin
        fsm_output = 10'b1101101000;
        state_var_NS = COMP_LOOP_C_675;
      end
      COMP_LOOP_C_675 : begin
        fsm_output = 10'b1101101001;
        if ( COMP_LOOP_C_675_tr0 ) begin
          state_var_NS = STAGE_VEC_LOOP_C_1;
        end
        else begin
          state_var_NS = COMP_LOOP_C_676;
        end
      end
      COMP_LOOP_C_676 : begin
        fsm_output = 10'b1101101010;
        state_var_NS = COMP_LOOP_C_677;
      end
      COMP_LOOP_C_677 : begin
        fsm_output = 10'b1101101011;
        state_var_NS = COMP_LOOP_C_678;
      end
      COMP_LOOP_C_678 : begin
        fsm_output = 10'b1101101100;
        state_var_NS = COMP_LOOP_C_679;
      end
      COMP_LOOP_C_679 : begin
        fsm_output = 10'b1101101101;
        state_var_NS = COMP_LOOP_C_680;
      end
      COMP_LOOP_C_680 : begin
        fsm_output = 10'b1101101110;
        state_var_NS = COMP_LOOP_C_681;
      end
      COMP_LOOP_C_681 : begin
        fsm_output = 10'b1101101111;
        state_var_NS = COMP_LOOP_C_682;
      end
      COMP_LOOP_C_682 : begin
        fsm_output = 10'b1101110000;
        state_var_NS = COMP_LOOP_C_683;
      end
      COMP_LOOP_C_683 : begin
        fsm_output = 10'b1101110001;
        state_var_NS = COMP_LOOP_C_684;
      end
      COMP_LOOP_C_684 : begin
        fsm_output = 10'b1101110010;
        state_var_NS = COMP_LOOP_C_685;
      end
      COMP_LOOP_C_685 : begin
        fsm_output = 10'b1101110011;
        state_var_NS = COMP_LOOP_C_686;
      end
      COMP_LOOP_C_686 : begin
        fsm_output = 10'b1101110100;
        state_var_NS = COMP_LOOP_C_687;
      end
      COMP_LOOP_C_687 : begin
        fsm_output = 10'b1101110101;
        state_var_NS = COMP_LOOP_C_688;
      end
      COMP_LOOP_C_688 : begin
        fsm_output = 10'b1101110110;
        state_var_NS = COMP_LOOP_C_689;
      end
      COMP_LOOP_C_689 : begin
        fsm_output = 10'b1101110111;
        state_var_NS = COMP_LOOP_C_690;
      end
      COMP_LOOP_C_690 : begin
        fsm_output = 10'b1101111000;
        state_var_NS = COMP_LOOP_C_691;
      end
      COMP_LOOP_C_691 : begin
        fsm_output = 10'b1101111001;
        state_var_NS = COMP_LOOP_16_modExp_dev_1_while_C_0;
      end
      COMP_LOOP_16_modExp_dev_1_while_C_0 : begin
        fsm_output = 10'b1101111010;
        state_var_NS = COMP_LOOP_16_modExp_dev_1_while_C_1;
      end
      COMP_LOOP_16_modExp_dev_1_while_C_1 : begin
        fsm_output = 10'b1101111011;
        state_var_NS = COMP_LOOP_16_modExp_dev_1_while_C_2;
      end
      COMP_LOOP_16_modExp_dev_1_while_C_2 : begin
        fsm_output = 10'b1101111100;
        state_var_NS = COMP_LOOP_16_modExp_dev_1_while_C_3;
      end
      COMP_LOOP_16_modExp_dev_1_while_C_3 : begin
        fsm_output = 10'b1101111101;
        state_var_NS = COMP_LOOP_16_modExp_dev_1_while_C_4;
      end
      COMP_LOOP_16_modExp_dev_1_while_C_4 : begin
        fsm_output = 10'b1101111110;
        state_var_NS = COMP_LOOP_16_modExp_dev_1_while_C_5;
      end
      COMP_LOOP_16_modExp_dev_1_while_C_5 : begin
        fsm_output = 10'b1101111111;
        state_var_NS = COMP_LOOP_16_modExp_dev_1_while_C_6;
      end
      COMP_LOOP_16_modExp_dev_1_while_C_6 : begin
        fsm_output = 10'b1110000000;
        state_var_NS = COMP_LOOP_16_modExp_dev_1_while_C_7;
      end
      COMP_LOOP_16_modExp_dev_1_while_C_7 : begin
        fsm_output = 10'b1110000001;
        state_var_NS = COMP_LOOP_16_modExp_dev_1_while_C_8;
      end
      COMP_LOOP_16_modExp_dev_1_while_C_8 : begin
        fsm_output = 10'b1110000010;
        state_var_NS = COMP_LOOP_16_modExp_dev_1_while_C_9;
      end
      COMP_LOOP_16_modExp_dev_1_while_C_9 : begin
        fsm_output = 10'b1110000011;
        state_var_NS = COMP_LOOP_16_modExp_dev_1_while_C_10;
      end
      COMP_LOOP_16_modExp_dev_1_while_C_10 : begin
        fsm_output = 10'b1110000100;
        state_var_NS = COMP_LOOP_16_modExp_dev_1_while_C_11;
      end
      COMP_LOOP_16_modExp_dev_1_while_C_11 : begin
        fsm_output = 10'b1110000101;
        if ( COMP_LOOP_16_modExp_dev_1_while_C_11_tr0 ) begin
          state_var_NS = COMP_LOOP_C_692;
        end
        else begin
          state_var_NS = COMP_LOOP_16_modExp_dev_1_while_C_0;
        end
      end
      COMP_LOOP_C_692 : begin
        fsm_output = 10'b1110000110;
        state_var_NS = COMP_LOOP_C_693;
      end
      COMP_LOOP_C_693 : begin
        fsm_output = 10'b1110000111;
        state_var_NS = COMP_LOOP_C_694;
      end
      COMP_LOOP_C_694 : begin
        fsm_output = 10'b1110001000;
        state_var_NS = COMP_LOOP_C_695;
      end
      COMP_LOOP_C_695 : begin
        fsm_output = 10'b1110001001;
        state_var_NS = COMP_LOOP_C_696;
      end
      COMP_LOOP_C_696 : begin
        fsm_output = 10'b1110001010;
        state_var_NS = COMP_LOOP_C_697;
      end
      COMP_LOOP_C_697 : begin
        fsm_output = 10'b1110001011;
        state_var_NS = COMP_LOOP_C_698;
      end
      COMP_LOOP_C_698 : begin
        fsm_output = 10'b1110001100;
        state_var_NS = COMP_LOOP_C_699;
      end
      COMP_LOOP_C_699 : begin
        fsm_output = 10'b1110001101;
        state_var_NS = COMP_LOOP_C_700;
      end
      COMP_LOOP_C_700 : begin
        fsm_output = 10'b1110001110;
        state_var_NS = COMP_LOOP_C_701;
      end
      COMP_LOOP_C_701 : begin
        fsm_output = 10'b1110001111;
        state_var_NS = COMP_LOOP_C_702;
      end
      COMP_LOOP_C_702 : begin
        fsm_output = 10'b1110010000;
        state_var_NS = COMP_LOOP_C_703;
      end
      COMP_LOOP_C_703 : begin
        fsm_output = 10'b1110010001;
        state_var_NS = COMP_LOOP_C_704;
      end
      COMP_LOOP_C_704 : begin
        fsm_output = 10'b1110010010;
        state_var_NS = COMP_LOOP_C_705;
      end
      COMP_LOOP_C_705 : begin
        fsm_output = 10'b1110010011;
        state_var_NS = COMP_LOOP_C_706;
      end
      COMP_LOOP_C_706 : begin
        fsm_output = 10'b1110010100;
        state_var_NS = COMP_LOOP_C_707;
      end
      COMP_LOOP_C_707 : begin
        fsm_output = 10'b1110010101;
        state_var_NS = COMP_LOOP_C_708;
      end
      COMP_LOOP_C_708 : begin
        fsm_output = 10'b1110010110;
        state_var_NS = COMP_LOOP_C_709;
      end
      COMP_LOOP_C_709 : begin
        fsm_output = 10'b1110010111;
        state_var_NS = COMP_LOOP_C_710;
      end
      COMP_LOOP_C_710 : begin
        fsm_output = 10'b1110011000;
        state_var_NS = COMP_LOOP_C_711;
      end
      COMP_LOOP_C_711 : begin
        fsm_output = 10'b1110011001;
        state_var_NS = COMP_LOOP_C_712;
      end
      COMP_LOOP_C_712 : begin
        fsm_output = 10'b1110011010;
        state_var_NS = COMP_LOOP_C_713;
      end
      COMP_LOOP_C_713 : begin
        fsm_output = 10'b1110011011;
        state_var_NS = COMP_LOOP_C_714;
      end
      COMP_LOOP_C_714 : begin
        fsm_output = 10'b1110011100;
        state_var_NS = COMP_LOOP_C_715;
      end
      COMP_LOOP_C_715 : begin
        fsm_output = 10'b1110011101;
        state_var_NS = COMP_LOOP_C_716;
      end
      COMP_LOOP_C_716 : begin
        fsm_output = 10'b1110011110;
        state_var_NS = COMP_LOOP_C_717;
      end
      COMP_LOOP_C_717 : begin
        fsm_output = 10'b1110011111;
        state_var_NS = COMP_LOOP_C_718;
      end
      COMP_LOOP_C_718 : begin
        fsm_output = 10'b1110100000;
        state_var_NS = COMP_LOOP_C_719;
      end
      COMP_LOOP_C_719 : begin
        fsm_output = 10'b1110100001;
        state_var_NS = COMP_LOOP_C_720;
      end
      COMP_LOOP_C_720 : begin
        fsm_output = 10'b1110100010;
        if ( COMP_LOOP_C_720_tr0 ) begin
          state_var_NS = STAGE_VEC_LOOP_C_1;
        end
        else begin
          state_var_NS = COMP_LOOP_C_0;
        end
      end
      STAGE_VEC_LOOP_C_1 : begin
        fsm_output = 10'b1110100011;
        if ( STAGE_VEC_LOOP_C_1_tr0 ) begin
          state_var_NS = STAGE_MAIN_LOOP_C_4;
        end
        else begin
          state_var_NS = STAGE_VEC_LOOP_C_0;
        end
      end
      STAGE_MAIN_LOOP_C_4 : begin
        fsm_output = 10'b1110100100;
        if ( STAGE_MAIN_LOOP_C_4_tr0 ) begin
          state_var_NS = main_C_1;
        end
        else begin
          state_var_NS = STAGE_MAIN_LOOP_C_0;
        end
      end
      main_C_1 : begin
        fsm_output = 10'b1110100101;
        state_var_NS = main_C_0;
      end
      // main_C_0
      default : begin
        fsm_output = 10'b0000000000;
        state_var_NS = STAGE_MAIN_LOOP_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( rst ) begin
      state_var <= main_C_0;
    end
    else begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_core_wait_dp
// ------------------------------------------------------------------


module inPlaceNTT_DIF_core_wait_dp (
  ensig_cgo_iro, ensig_cgo, COMP_LOOP_1_modulo_dev_cmp_ccs_ccore_en
);
  input ensig_cgo_iro;
  input ensig_cgo;
  output COMP_LOOP_1_modulo_dev_cmp_ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  assign COMP_LOOP_1_modulo_dev_cmp_ccs_ccore_en = ensig_cgo | ensig_cgo_iro;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_core
// ------------------------------------------------------------------


module inPlaceNTT_DIF_core (
  clk, rst, vec_rsc_triosy_0_0_lz, vec_rsc_triosy_0_1_lz, vec_rsc_triosy_0_2_lz,
      vec_rsc_triosy_0_3_lz, vec_rsc_triosy_0_4_lz, vec_rsc_triosy_0_5_lz, vec_rsc_triosy_0_6_lz,
      vec_rsc_triosy_0_7_lz, vec_rsc_triosy_0_8_lz, vec_rsc_triosy_0_9_lz, vec_rsc_triosy_0_10_lz,
      vec_rsc_triosy_0_11_lz, vec_rsc_triosy_0_12_lz, vec_rsc_triosy_0_13_lz, vec_rsc_triosy_0_14_lz,
      vec_rsc_triosy_0_15_lz, p_rsc_dat, p_rsc_triosy_lz, r_rsc_dat, r_rsc_triosy_lz,
      vec_rsc_0_0_i_qa_d, vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d, vec_rsc_0_1_i_qa_d,
      vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d, vec_rsc_0_2_i_qa_d, vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_3_i_qa_d, vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d, vec_rsc_0_4_i_qa_d,
      vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d, vec_rsc_0_5_i_qa_d, vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_6_i_qa_d, vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d, vec_rsc_0_7_i_qa_d,
      vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d, vec_rsc_0_8_i_qa_d, vec_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_9_i_qa_d, vec_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d, vec_rsc_0_10_i_qa_d,
      vec_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d, vec_rsc_0_11_i_qa_d, vec_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_12_i_qa_d, vec_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d, vec_rsc_0_13_i_qa_d,
      vec_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d, vec_rsc_0_14_i_qa_d, vec_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_15_i_qa_d, vec_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d, vec_rsc_0_0_i_adra_d_pff,
      vec_rsc_0_0_i_da_d_pff, vec_rsc_0_0_i_wea_d_pff, vec_rsc_0_1_i_wea_d_pff, vec_rsc_0_2_i_wea_d_pff,
      vec_rsc_0_3_i_wea_d_pff, vec_rsc_0_4_i_wea_d_pff, vec_rsc_0_5_i_wea_d_pff,
      vec_rsc_0_6_i_wea_d_pff, vec_rsc_0_7_i_wea_d_pff, vec_rsc_0_8_i_wea_d_pff,
      vec_rsc_0_9_i_wea_d_pff, vec_rsc_0_10_i_wea_d_pff, vec_rsc_0_11_i_wea_d_pff,
      vec_rsc_0_12_i_wea_d_pff, vec_rsc_0_13_i_wea_d_pff, vec_rsc_0_14_i_wea_d_pff,
      vec_rsc_0_15_i_wea_d_pff
);
  input clk;
  input rst;
  output vec_rsc_triosy_0_0_lz;
  output vec_rsc_triosy_0_1_lz;
  output vec_rsc_triosy_0_2_lz;
  output vec_rsc_triosy_0_3_lz;
  output vec_rsc_triosy_0_4_lz;
  output vec_rsc_triosy_0_5_lz;
  output vec_rsc_triosy_0_6_lz;
  output vec_rsc_triosy_0_7_lz;
  output vec_rsc_triosy_0_8_lz;
  output vec_rsc_triosy_0_9_lz;
  output vec_rsc_triosy_0_10_lz;
  output vec_rsc_triosy_0_11_lz;
  output vec_rsc_triosy_0_12_lz;
  output vec_rsc_triosy_0_13_lz;
  output vec_rsc_triosy_0_14_lz;
  output vec_rsc_triosy_0_15_lz;
  input [63:0] p_rsc_dat;
  output p_rsc_triosy_lz;
  input [63:0] r_rsc_dat;
  output r_rsc_triosy_lz;
  input [63:0] vec_rsc_0_0_i_qa_d;
  output vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_1_i_qa_d;
  output vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_2_i_qa_d;
  output vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_3_i_qa_d;
  output vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_4_i_qa_d;
  output vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_5_i_qa_d;
  output vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_6_i_qa_d;
  output vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_7_i_qa_d;
  output vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_8_i_qa_d;
  output vec_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_9_i_qa_d;
  output vec_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_10_i_qa_d;
  output vec_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_11_i_qa_d;
  output vec_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_12_i_qa_d;
  output vec_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_13_i_qa_d;
  output vec_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_14_i_qa_d;
  output vec_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_15_i_qa_d;
  output vec_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [5:0] vec_rsc_0_0_i_adra_d_pff;
  output [63:0] vec_rsc_0_0_i_da_d_pff;
  output vec_rsc_0_0_i_wea_d_pff;
  output vec_rsc_0_1_i_wea_d_pff;
  output vec_rsc_0_2_i_wea_d_pff;
  output vec_rsc_0_3_i_wea_d_pff;
  output vec_rsc_0_4_i_wea_d_pff;
  output vec_rsc_0_5_i_wea_d_pff;
  output vec_rsc_0_6_i_wea_d_pff;
  output vec_rsc_0_7_i_wea_d_pff;
  output vec_rsc_0_8_i_wea_d_pff;
  output vec_rsc_0_9_i_wea_d_pff;
  output vec_rsc_0_10_i_wea_d_pff;
  output vec_rsc_0_11_i_wea_d_pff;
  output vec_rsc_0_12_i_wea_d_pff;
  output vec_rsc_0_13_i_wea_d_pff;
  output vec_rsc_0_14_i_wea_d_pff;
  output vec_rsc_0_15_i_wea_d_pff;


  // Interconnect Declarations
  wire [63:0] p_rsci_idat;
  wire [63:0] r_rsci_idat;
  wire [63:0] COMP_LOOP_1_modulo_dev_cmp_return_rsc_z;
  wire COMP_LOOP_1_modulo_dev_cmp_ccs_ccore_en;
  reg [63:0] modExp_dev_while_rem_cmp_a;
  wire [63:0] modExp_dev_while_rem_cmp_z;
  reg [63:0] STAGE_MAIN_LOOP_div_cmp_a;
  reg [9:0] STAGE_MAIN_LOOP_div_cmp_b;
  wire [63:0] STAGE_MAIN_LOOP_div_cmp_z;
  wire [9:0] fsm_output;
  wire [9:0] COMP_LOOP_1_operator_64_false_acc_tmp;
  wire [11:0] nl_COMP_LOOP_1_operator_64_false_acc_tmp;
  wire or_tmp;
  wire nor_tmp_1;
  wire nor_tmp_3;
  wire and_dcpl;
  wire and_dcpl_5;
  wire or_tmp_33;
  wire mux_tmp_79;
  wire nor_tmp_87;
  wire mux_tmp_302;
  wire or_tmp_235;
  wire nor_tmp_130;
  wire and_tmp_11;
  wire and_dcpl_44;
  wire and_dcpl_70;
  wire not_tmp_266;
  wire and_dcpl_91;
  wire and_dcpl_92;
  wire and_dcpl_93;
  wire and_dcpl_94;
  wire and_dcpl_95;
  wire and_dcpl_96;
  wire and_dcpl_97;
  wire and_dcpl_98;
  wire or_tmp_546;
  wire and_dcpl_105;
  wire and_dcpl_106;
  wire and_dcpl_109;
  wire xor_dcpl;
  wire and_dcpl_113;
  wire not_tmp_280;
  wire and_dcpl_125;
  wire and_dcpl_131;
  wire and_dcpl_135;
  wire and_dcpl_143;
  wire and_dcpl_146;
  wire and_dcpl_147;
  wire and_dcpl_158;
  wire and_dcpl_159;
  wire not_tmp_292;
  wire and_dcpl_176;
  wire and_dcpl_192;
  wire and_dcpl_199;
  wire or_tmp_591;
  wire and_dcpl_225;
  wire not_tmp_311;
  wire not_tmp_312;
  wire nand_tmp_16;
  wire or_tmp_669;
  wire nand_tmp_19;
  wire not_tmp_322;
  wire nand_tmp_22;
  wire nand_tmp_28;
  wire nand_tmp_34;
  wire nand_tmp_40;
  wire nand_tmp_46;
  wire nand_tmp_52;
  wire nand_tmp_58;
  wire nand_tmp_64;
  wire nand_tmp_70;
  wire nand_tmp_76;
  wire nand_tmp_82;
  wire nand_tmp_88;
  wire nand_tmp_94;
  wire nand_tmp_100;
  wire nand_tmp_106;
  wire or_tmp_2322;
  wire mux_tmp_2110;
  wire mux_tmp_2111;
  wire mux_tmp_2112;
  wire mux_tmp_2113;
  wire or_tmp_2324;
  wire mux_tmp_2114;
  wire mux_tmp_2118;
  wire mux_tmp_2124;
  wire mux_tmp_2127;
  wire mux_tmp_2129;
  wire mux_tmp_2130;
  wire mux_tmp_2131;
  wire mux_tmp_2132;
  wire mux_tmp_2135;
  wire mux_tmp_2139;
  wire mux_tmp_2142;
  wire nor_tmp_357;
  wire mux_tmp_2161;
  wire and_dcpl_239;
  wire and_dcpl_240;
  wire or_tmp_2348;
  wire or_tmp_2352;
  wire or_tmp_2355;
  wire and_dcpl_241;
  wire and_dcpl_242;
  wire and_dcpl_243;
  wire and_dcpl_244;
  wire and_dcpl_245;
  wire and_dcpl_246;
  wire and_dcpl_248;
  wire and_dcpl_249;
  wire and_dcpl_251;
  wire and_dcpl_252;
  wire and_dcpl_253;
  wire and_dcpl_254;
  wire and_dcpl_255;
  wire and_dcpl_256;
  wire and_dcpl_257;
  wire and_dcpl_258;
  wire and_dcpl_259;
  wire and_dcpl_260;
  wire and_dcpl_261;
  wire and_dcpl_262;
  wire and_dcpl_263;
  wire and_dcpl_264;
  wire and_dcpl_265;
  wire and_dcpl_266;
  wire and_dcpl_267;
  wire and_dcpl_268;
  wire and_dcpl_269;
  wire and_dcpl_270;
  wire and_dcpl_271;
  wire and_dcpl_273;
  wire and_dcpl_275;
  wire and_dcpl_276;
  wire and_dcpl_278;
  wire and_dcpl_279;
  wire and_dcpl_280;
  wire and_dcpl_282;
  wire and_dcpl_283;
  wire and_dcpl_284;
  wire and_dcpl_285;
  wire and_dcpl_286;
  wire and_dcpl_287;
  wire and_dcpl_288;
  wire and_dcpl_289;
  wire or_tmp_2368;
  wire mux_tmp_2215;
  wire mux_tmp_2216;
  wire or_tmp_2373;
  wire or_tmp_2381;
  wire mux_tmp_2223;
  wire mux_tmp_2226;
  wire and_dcpl_290;
  wire or_tmp_2391;
  wire or_tmp_2393;
  wire or_tmp_2395;
  wire mux_tmp_2244;
  wire or_tmp_2401;
  wire or_tmp_2402;
  wire mux_tmp_2247;
  wire or_tmp_2406;
  wire mux_tmp_2250;
  wire not_tmp_572;
  wire or_tmp_2409;
  wire mux_tmp_2276;
  wire and_dcpl_293;
  wire and_dcpl_294;
  wire and_dcpl_295;
  wire or_tmp_2439;
  wire and_tmp_24;
  wire nor_tmp_388;
  wire or_tmp_2447;
  wire or_tmp_2451;
  wire not_tmp_597;
  wire mux_tmp_2377;
  wire or_tmp_2548;
  wire or_tmp_2549;
  wire mux_tmp_2380;
  wire nor_tmp_399;
  wire mux_tmp_2381;
  wire mux_tmp_2382;
  wire not_tmp_617;
  wire mux_tmp_2389;
  wire or_tmp_2551;
  wire or_tmp_2552;
  wire mux_tmp_2400;
  wire nor_tmp_403;
  wire and_dcpl_307;
  wire and_dcpl_311;
  wire and_dcpl_313;
  wire and_dcpl_317;
  wire and_dcpl_319;
  wire and_dcpl_321;
  wire and_dcpl_323;
  wire and_dcpl_329;
  wire and_dcpl_331;
  wire and_dcpl_345;
  wire and_dcpl_346;
  wire mux_tmp_2449;
  wire mux_tmp_2450;
  wire or_dcpl_72;
  wire mux_tmp_2457;
  wire mux_tmp_2458;
  wire mux_tmp_2459;
  wire or_tmp_2585;
  wire mux_tmp_2461;
  wire mux_tmp_2462;
  wire mux_tmp_2467;
  wire mux_tmp_2468;
  wire or_tmp_2587;
  wire mux_tmp_2469;
  wire mux_tmp_2470;
  wire or_tmp_2588;
  wire mux_tmp_2474;
  wire nand_tmp_140;
  wire nor_tmp_417;
  wire mux_tmp_2529;
  wire not_tmp_662;
  wire mux_tmp_2538;
  wire not_tmp_664;
  wire and_dcpl_354;
  wire and_dcpl_357;
  wire and_dcpl_359;
  wire nor_tmp_427;
  wire and_dcpl_361;
  wire mux_tmp_2574;
  wire or_tmp_2638;
  wire mux_tmp_2583;
  wire and_dcpl_364;
  wire and_dcpl_367;
  wire and_dcpl_370;
  wire not_tmp_696;
  wire not_tmp_698;
  wire and_dcpl_372;
  wire mux_tmp_2612;
  wire not_tmp_703;
  wire mux_tmp_2614;
  wire not_tmp_706;
  wire or_tmp_2668;
  wire and_tmp_32;
  wire mux_tmp_2625;
  wire mux_tmp_2626;
  wire nor_tmp_459;
  wire mux_tmp_2653;
  wire nor_tmp_463;
  wire nor_tmp_467;
  wire mux_tmp_2666;
  wire not_tmp_729;
  wire mux_tmp_2689;
  wire mux_tmp_2713;
  wire mux_tmp_2714;
  wire mux_tmp_2720;
  wire or_tmp_2733;
  wire or_tmp_2734;
  wire mux_tmp_2721;
  wire or_tmp_2735;
  wire or_tmp_2736;
  wire mux_tmp_2724;
  wire nand_tmp_148;
  reg COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm;
  reg operator_64_false_1_slc_operator_64_false_1_acc_5_itm;
  wire [7:0] COMP_LOOP_acc_8_psp_sva_1;
  wire [8:0] nl_COMP_LOOP_acc_8_psp_sva_1;
  reg [4:0] COMP_LOOP_k_9_4_sva_4_0;
  wire [9:0] COMP_LOOP_acc_cse_4_sva_1;
  wire [10:0] nl_COMP_LOOP_acc_cse_4_sva_1;
  reg [9:0] STAGE_VEC_LOOP_j_sva_9_0;
  reg operator_64_false_slc_operator_64_false_acc_1_60_itm;
  reg [9:0] operator_64_false_acc_cse_sva;
  reg [9:0] operator_64_false_acc_cse_12_sva;
  reg [7:0] COMP_LOOP_acc_12_psp_sva;
  reg [8:0] COMP_LOOP_acc_7_psp_sva;
  wire [9:0] nl_COMP_LOOP_acc_7_psp_sva;
  reg [9:0] operator_64_false_acc_cse_2_sva;
  reg [9:0] operator_64_false_acc_cse_8_sva;
  reg [6:0] COMP_LOOP_acc_10_psp_sva;
  wire [7:0] nl_COMP_LOOP_acc_10_psp_sva;
  reg [9:0] operator_64_false_acc_cse_4_sva;
  reg [8:0] COMP_LOOP_acc_13_psp_sva;
  wire [9:0] nl_COMP_LOOP_acc_13_psp_sva;
  reg [9:0] operator_64_false_acc_cse_14_sva;
  reg [8:0] COMP_LOOP_acc_11_psp_sva;
  wire [9:0] nl_COMP_LOOP_acc_11_psp_sva;
  reg [9:0] operator_64_false_acc_cse_10_sva;
  reg [8:0] COMP_LOOP_acc_9_psp_sva;
  wire [9:0] nl_COMP_LOOP_acc_9_psp_sva;
  reg [9:0] operator_64_false_acc_cse_6_sva;
  reg [7:0] COMP_LOOP_acc_8_psp_sva;
  reg [9:0] operator_64_false_acc_cse_13_sva;
  reg [9:0] COMP_LOOP_acc_cse_12_sva;
  wire [10:0] nl_COMP_LOOP_acc_cse_12_sva;
  reg [9:0] operator_64_false_acc_cse_11_sva;
  reg [9:0] COMP_LOOP_acc_cse_8_sva;
  wire [10:0] nl_COMP_LOOP_acc_cse_8_sva;
  reg [9:0] operator_64_false_acc_cse_7_sva;
  reg [9:0] operator_64_false_acc_cse_3_sva;
  reg [9:0] COMP_LOOP_acc_cse_4_sva;
  reg [9:0] COMP_LOOP_acc_cse_14_sva;
  wire [10:0] nl_COMP_LOOP_acc_cse_14_sva;
  reg [9:0] operator_64_false_acc_cse_9_sva;
  reg [9:0] COMP_LOOP_acc_cse_10_sva;
  wire [10:0] nl_COMP_LOOP_acc_cse_10_sva;
  reg [9:0] COMP_LOOP_acc_cse_sva;
  wire [10:0] nl_COMP_LOOP_acc_cse_sva;
  reg [9:0] operator_64_false_acc_cse_15_sva;
  reg [9:0] COMP_LOOP_acc_cse_6_sva;
  reg [9:0] operator_64_false_acc_cse_5_sva;
  reg [9:0] COMP_LOOP_acc_cse_2_sva;
  reg [9:0] operator_64_false_acc_cse_1_sva;
  reg [9:0] STAGE_MAIN_LOOP_lshift_psp_1_sva;
  wire [9:0] COMP_LOOP_acc_cse_2_sva_1;
  wire [10:0] nl_COMP_LOOP_acc_cse_2_sva_1;
  wire [9:0] operator_64_false_acc_cse_2_sva_mx0w0;
  wire [11:0] nl_operator_64_false_acc_cse_2_sva_mx0w0;
  wire [9:0] operator_64_false_acc_cse_3_sva_mx0w0;
  wire [11:0] nl_operator_64_false_acc_cse_3_sva_mx0w0;
  wire [9:0] operator_64_false_acc_cse_4_sva_mx0w0;
  wire [11:0] nl_operator_64_false_acc_cse_4_sva_mx0w0;
  wire [9:0] operator_64_false_acc_cse_5_sva_mx0w0;
  wire [11:0] nl_operator_64_false_acc_cse_5_sva_mx0w0;
  wire [9:0] operator_64_false_acc_cse_6_sva_mx0w0;
  wire [11:0] nl_operator_64_false_acc_cse_6_sva_mx0w0;
  wire [9:0] operator_64_false_acc_cse_7_sva_mx0w0;
  wire [11:0] nl_operator_64_false_acc_cse_7_sva_mx0w0;
  wire [9:0] operator_64_false_acc_cse_8_sva_mx0w0;
  wire [11:0] nl_operator_64_false_acc_cse_8_sva_mx0w0;
  wire [9:0] operator_64_false_acc_cse_9_sva_mx0w0;
  wire [11:0] nl_operator_64_false_acc_cse_9_sva_mx0w0;
  wire [9:0] operator_64_false_acc_cse_10_sva_mx0w0;
  wire [11:0] nl_operator_64_false_acc_cse_10_sva_mx0w0;
  wire [9:0] operator_64_false_acc_cse_11_sva_mx0w0;
  wire [11:0] nl_operator_64_false_acc_cse_11_sva_mx0w0;
  wire [9:0] operator_64_false_acc_cse_12_sva_mx0w0;
  wire [11:0] nl_operator_64_false_acc_cse_12_sva_mx0w0;
  wire [9:0] operator_64_false_acc_cse_13_sva_mx0w0;
  wire [11:0] nl_operator_64_false_acc_cse_13_sva_mx0w0;
  wire [9:0] operator_64_false_acc_cse_14_sva_mx0w0;
  wire [11:0] nl_operator_64_false_acc_cse_14_sva_mx0w0;
  wire [9:0] operator_64_false_acc_cse_15_sva_mx0w0;
  wire [11:0] nl_operator_64_false_acc_cse_15_sva_mx0w0;
  wire [9:0] operator_64_false_acc_cse_sva_mx0w0;
  wire [11:0] nl_operator_64_false_acc_cse_sva_mx0w0;
  wire and_332_m1c;
  wire and_334_m1c;
  wire and_335_m1c;
  wire and_338_m1c;
  wire and_340_m1c;
  wire and_342_m1c;
  wire and_344_m1c;
  wire and_346_m1c;
  wire and_348_m1c;
  wire and_350_m1c;
  wire and_351_m1c;
  wire and_352_m1c;
  wire and_354_m1c;
  wire and_356_m1c;
  wire and_358_m1c;
  wire nand_437_cse;
  reg reg_vec_rsc_triosy_0_15_obj_ld_cse;
  reg reg_ensig_cgo_cse;
  wire nor_368_cse;
  wire and_516_cse;
  wire and_515_cse;
  reg [63:0] reg_COMP_LOOP_1_modulo_dev_cmp_m_rsc_dat_cse;
  wire or_602_cse;
  wire or_2500_cse;
  wire or_2700_cse;
  wire or_598_cse;
  wire and_697_cse;
  wire and_711_cse;
  wire or_111_cse;
  wire and_581_cse;
  wire or_307_cse;
  wire or_165_cse;
  wire nor_813_cse;
  wire or_420_cse;
  wire and_459_cse;
  wire and_623_cse;
  wire and_679_cse;
  wire or_2733_cse;
  wire and_756_cse;
  wire nor_936_cse;
  wire and_475_cse;
  wire and_613_cse;
  wire nor_832_cse;
  wire nand_442_cse;
  wire or_694_cse;
  wire or_803_cse;
  wire or_909_cse;
  wire or_1018_cse;
  wire or_1124_cse;
  wire or_1233_cse;
  wire or_1339_cse;
  wire or_1448_cse;
  wire nand_169_cse;
  wire nand_445_cse;
  wire mux_2252_cse;
  wire or_2573_cse;
  wire or_204_cse;
  wire mux_156_cse;
  wire nor_510_cse;
  wire mux_494_cse;
  wire nor_569_cse;
  wire nor_497_cse;
  wire mux_2374_cse;
  wire or_2549_cse;
  wire nor_558_cse;
  wire mux_792_cse;
  wire mux_79_cse;
  wire mux_1112_cse;
  wire mux_1031_cse;
  reg COMP_LOOP_COMP_LOOP_nor_itm;
  reg COMP_LOOP_COMP_LOOP_and_244_itm;
  reg COMP_LOOP_COMP_LOOP_and_62_itm;
  reg COMP_LOOP_COMP_LOOP_and_185_itm;
  reg COMP_LOOP_COMP_LOOP_and_64_itm;
  reg COMP_LOOP_COMP_LOOP_and_65_itm;
  reg COMP_LOOP_COMP_LOOP_and_66_itm;
  reg COMP_LOOP_COMP_LOOP_and_6_itm;
  reg COMP_LOOP_COMP_LOOP_and_68_itm;
  reg COMP_LOOP_COMP_LOOP_and_69_itm;
  reg COMP_LOOP_COMP_LOOP_and_70_itm;
  reg COMP_LOOP_COMP_LOOP_and_10_itm;
  reg COMP_LOOP_COMP_LOOP_and_72_itm;
  reg COMP_LOOP_COMP_LOOP_and_12_itm;
  reg COMP_LOOP_COMP_LOOP_and_13_itm;
  reg COMP_LOOP_COMP_LOOP_and_14_itm;
  reg [63:0] tmp_1_lpi_4_dfm;
  reg [63:0] tmp_10_lpi_4_dfm;
  reg [63:0] COMP_LOOP_10_modExp_dev_1_while_mul_mut;
  reg COMP_LOOP_COMP_LOOP_nor_5_itm;
  reg COMP_LOOP_nor_51_itm;
  reg COMP_LOOP_nor_52_itm;
  reg COMP_LOOP_COMP_LOOP_and_77_itm;
  reg COMP_LOOP_nor_54_itm;
  reg COMP_LOOP_COMP_LOOP_and_79_itm;
  reg COMP_LOOP_COMP_LOOP_and_80_itm;
  reg COMP_LOOP_COMP_LOOP_and_81_itm;
  reg COMP_LOOP_nor_57_itm;
  reg COMP_LOOP_COMP_LOOP_and_83_itm;
  reg COMP_LOOP_COMP_LOOP_and_84_itm;
  reg COMP_LOOP_COMP_LOOP_and_85_itm;
  reg COMP_LOOP_COMP_LOOP_and_86_itm;
  reg COMP_LOOP_COMP_LOOP_and_87_itm;
  reg COMP_LOOP_COMP_LOOP_and_88_itm;
  reg COMP_LOOP_COMP_LOOP_and_89_itm;
  reg COMP_LOOP_COMP_LOOP_nor_9_itm;
  reg COMP_LOOP_nor_91_itm;
  reg COMP_LOOP_nor_92_itm;
  reg COMP_LOOP_COMP_LOOP_and_137_itm;
  reg COMP_LOOP_nor_94_itm;
  reg COMP_LOOP_COMP_LOOP_and_139_itm;
  reg COMP_LOOP_COMP_LOOP_and_140_itm;
  reg COMP_LOOP_COMP_LOOP_and_141_itm;
  reg COMP_LOOP_nor_97_itm;
  reg COMP_LOOP_COMP_LOOP_and_143_itm;
  reg COMP_LOOP_COMP_LOOP_and_144_itm;
  reg COMP_LOOP_COMP_LOOP_and_145_itm;
  reg COMP_LOOP_COMP_LOOP_and_146_itm;
  reg COMP_LOOP_COMP_LOOP_and_147_itm;
  reg COMP_LOOP_COMP_LOOP_and_148_itm;
  reg COMP_LOOP_COMP_LOOP_and_149_itm;
  reg COMP_LOOP_COMP_LOOP_nor_13_itm;
  reg COMP_LOOP_nor_131_itm;
  reg COMP_LOOP_nor_132_itm;
  reg COMP_LOOP_COMP_LOOP_and_197_itm;
  reg COMP_LOOP_nor_134_itm;
  reg COMP_LOOP_COMP_LOOP_and_199_itm;
  reg COMP_LOOP_COMP_LOOP_and_200_itm;
  reg COMP_LOOP_COMP_LOOP_and_201_itm;
  reg COMP_LOOP_nor_137_itm;
  reg COMP_LOOP_COMP_LOOP_and_203_itm;
  reg COMP_LOOP_COMP_LOOP_and_204_itm;
  reg COMP_LOOP_COMP_LOOP_and_205_itm;
  reg COMP_LOOP_COMP_LOOP_and_206_itm;
  reg COMP_LOOP_COMP_LOOP_and_207_itm;
  reg COMP_LOOP_COMP_LOOP_and_208_itm;
  reg COMP_LOOP_COMP_LOOP_and_209_itm;
  reg COMP_LOOP_COMP_LOOP_nor_17_itm;
  reg COMP_LOOP_nor_171_itm;
  reg COMP_LOOP_nor_172_itm;
  reg COMP_LOOP_COMP_LOOP_and_257_itm;
  reg COMP_LOOP_nor_174_itm;
  reg COMP_LOOP_COMP_LOOP_and_259_itm;
  reg COMP_LOOP_COMP_LOOP_and_260_itm;
  reg COMP_LOOP_COMP_LOOP_and_261_itm;
  reg COMP_LOOP_nor_177_itm;
  reg COMP_LOOP_COMP_LOOP_and_263_itm;
  reg COMP_LOOP_COMP_LOOP_and_264_itm;
  reg COMP_LOOP_COMP_LOOP_and_265_itm;
  reg COMP_LOOP_COMP_LOOP_and_266_itm;
  reg COMP_LOOP_COMP_LOOP_and_267_itm;
  reg COMP_LOOP_COMP_LOOP_and_268_itm;
  reg COMP_LOOP_COMP_LOOP_and_269_itm;
  reg COMP_LOOP_COMP_LOOP_nor_21_itm;
  reg COMP_LOOP_nor_211_itm;
  reg COMP_LOOP_nor_212_itm;
  reg COMP_LOOP_COMP_LOOP_and_317_itm;
  reg COMP_LOOP_nor_214_itm;
  reg COMP_LOOP_COMP_LOOP_and_319_itm;
  reg COMP_LOOP_COMP_LOOP_and_320_itm;
  reg COMP_LOOP_COMP_LOOP_and_321_itm;
  reg COMP_LOOP_nor_217_itm;
  reg COMP_LOOP_COMP_LOOP_and_323_itm;
  reg COMP_LOOP_COMP_LOOP_and_324_itm;
  reg COMP_LOOP_COMP_LOOP_and_325_itm;
  reg COMP_LOOP_COMP_LOOP_and_326_itm;
  reg COMP_LOOP_COMP_LOOP_and_327_itm;
  reg COMP_LOOP_COMP_LOOP_and_328_itm;
  reg COMP_LOOP_COMP_LOOP_and_329_itm;
  reg COMP_LOOP_COMP_LOOP_nor_25_itm;
  reg COMP_LOOP_nor_251_itm;
  reg COMP_LOOP_nor_252_itm;
  reg COMP_LOOP_COMP_LOOP_and_377_itm;
  reg COMP_LOOP_nor_254_itm;
  reg COMP_LOOP_COMP_LOOP_and_379_itm;
  reg COMP_LOOP_COMP_LOOP_and_380_itm;
  reg COMP_LOOP_COMP_LOOP_and_381_itm;
  reg COMP_LOOP_nor_257_itm;
  reg COMP_LOOP_COMP_LOOP_and_383_itm;
  reg COMP_LOOP_COMP_LOOP_and_384_itm;
  reg COMP_LOOP_COMP_LOOP_and_385_itm;
  reg COMP_LOOP_COMP_LOOP_and_386_itm;
  reg COMP_LOOP_COMP_LOOP_and_387_itm;
  reg COMP_LOOP_COMP_LOOP_and_388_itm;
  reg COMP_LOOP_COMP_LOOP_and_389_itm;
  reg COMP_LOOP_COMP_LOOP_nor_29_itm;
  reg COMP_LOOP_nor_291_itm;
  reg COMP_LOOP_nor_292_itm;
  reg COMP_LOOP_COMP_LOOP_and_437_itm;
  reg COMP_LOOP_nor_294_itm;
  reg COMP_LOOP_COMP_LOOP_and_439_itm;
  reg COMP_LOOP_COMP_LOOP_and_440_itm;
  reg COMP_LOOP_COMP_LOOP_and_441_itm;
  reg COMP_LOOP_nor_297_itm;
  reg COMP_LOOP_COMP_LOOP_and_443_itm;
  reg COMP_LOOP_COMP_LOOP_and_444_itm;
  reg COMP_LOOP_COMP_LOOP_and_445_itm;
  reg COMP_LOOP_COMP_LOOP_and_446_itm;
  reg COMP_LOOP_COMP_LOOP_and_447_itm;
  reg COMP_LOOP_COMP_LOOP_and_448_itm;
  reg COMP_LOOP_COMP_LOOP_and_449_itm;
  reg COMP_LOOP_COMP_LOOP_nor_33_itm;
  reg COMP_LOOP_nor_331_itm;
  reg COMP_LOOP_nor_332_itm;
  reg COMP_LOOP_COMP_LOOP_and_497_itm;
  reg COMP_LOOP_nor_334_itm;
  reg COMP_LOOP_COMP_LOOP_and_499_itm;
  reg COMP_LOOP_COMP_LOOP_and_500_itm;
  reg COMP_LOOP_COMP_LOOP_and_501_itm;
  reg COMP_LOOP_nor_337_itm;
  reg COMP_LOOP_COMP_LOOP_and_503_itm;
  reg COMP_LOOP_COMP_LOOP_and_504_itm;
  reg COMP_LOOP_COMP_LOOP_and_505_itm;
  reg COMP_LOOP_COMP_LOOP_and_506_itm;
  reg COMP_LOOP_COMP_LOOP_and_507_itm;
  reg COMP_LOOP_COMP_LOOP_and_508_itm;
  reg COMP_LOOP_COMP_LOOP_and_509_itm;
  reg COMP_LOOP_COMP_LOOP_nor_37_itm;
  reg COMP_LOOP_nor_371_itm;
  reg COMP_LOOP_nor_372_itm;
  reg COMP_LOOP_COMP_LOOP_and_557_itm;
  reg COMP_LOOP_nor_374_itm;
  reg COMP_LOOP_COMP_LOOP_and_559_itm;
  reg COMP_LOOP_COMP_LOOP_and_560_itm;
  reg COMP_LOOP_COMP_LOOP_and_561_itm;
  reg COMP_LOOP_nor_377_itm;
  reg COMP_LOOP_COMP_LOOP_and_563_itm;
  reg COMP_LOOP_COMP_LOOP_and_564_itm;
  reg COMP_LOOP_COMP_LOOP_and_565_itm;
  reg COMP_LOOP_COMP_LOOP_and_566_itm;
  reg COMP_LOOP_COMP_LOOP_and_567_itm;
  reg COMP_LOOP_COMP_LOOP_and_568_itm;
  reg COMP_LOOP_COMP_LOOP_and_569_itm;
  reg COMP_LOOP_COMP_LOOP_nor_41_itm;
  reg COMP_LOOP_nor_411_itm;
  reg COMP_LOOP_nor_412_itm;
  reg COMP_LOOP_COMP_LOOP_and_617_itm;
  reg COMP_LOOP_nor_414_itm;
  reg COMP_LOOP_COMP_LOOP_and_619_itm;
  reg COMP_LOOP_COMP_LOOP_and_620_itm;
  reg COMP_LOOP_COMP_LOOP_and_621_itm;
  reg COMP_LOOP_nor_417_itm;
  reg COMP_LOOP_COMP_LOOP_and_623_itm;
  reg COMP_LOOP_COMP_LOOP_and_624_itm;
  reg COMP_LOOP_COMP_LOOP_and_625_itm;
  reg COMP_LOOP_COMP_LOOP_and_626_itm;
  reg COMP_LOOP_COMP_LOOP_and_627_itm;
  reg COMP_LOOP_COMP_LOOP_and_628_itm;
  reg COMP_LOOP_COMP_LOOP_and_629_itm;
  reg COMP_LOOP_COMP_LOOP_nor_45_itm;
  reg COMP_LOOP_nor_451_itm;
  reg COMP_LOOP_nor_452_itm;
  reg COMP_LOOP_COMP_LOOP_and_677_itm;
  reg COMP_LOOP_nor_454_itm;
  reg COMP_LOOP_COMP_LOOP_and_679_itm;
  reg COMP_LOOP_COMP_LOOP_and_680_itm;
  reg COMP_LOOP_COMP_LOOP_and_681_itm;
  reg COMP_LOOP_nor_457_itm;
  reg COMP_LOOP_COMP_LOOP_and_683_itm;
  reg COMP_LOOP_COMP_LOOP_and_684_itm;
  reg COMP_LOOP_COMP_LOOP_and_685_itm;
  reg COMP_LOOP_COMP_LOOP_and_686_itm;
  reg COMP_LOOP_COMP_LOOP_and_687_itm;
  reg COMP_LOOP_COMP_LOOP_and_688_itm;
  reg COMP_LOOP_COMP_LOOP_and_689_itm;
  reg COMP_LOOP_COMP_LOOP_nor_49_itm;
  reg COMP_LOOP_nor_491_itm;
  reg COMP_LOOP_nor_492_itm;
  reg COMP_LOOP_COMP_LOOP_and_737_itm;
  reg COMP_LOOP_nor_494_itm;
  reg COMP_LOOP_COMP_LOOP_and_739_itm;
  reg COMP_LOOP_COMP_LOOP_and_740_itm;
  reg COMP_LOOP_COMP_LOOP_and_741_itm;
  reg COMP_LOOP_nor_497_itm;
  reg COMP_LOOP_COMP_LOOP_and_743_itm;
  reg COMP_LOOP_COMP_LOOP_and_744_itm;
  reg COMP_LOOP_COMP_LOOP_and_745_itm;
  reg COMP_LOOP_COMP_LOOP_and_746_itm;
  reg COMP_LOOP_COMP_LOOP_and_747_itm;
  reg COMP_LOOP_COMP_LOOP_and_748_itm;
  reg COMP_LOOP_COMP_LOOP_and_749_itm;
  reg COMP_LOOP_COMP_LOOP_nor_53_itm;
  reg COMP_LOOP_nor_531_itm;
  reg COMP_LOOP_nor_532_itm;
  reg COMP_LOOP_COMP_LOOP_and_797_itm;
  reg COMP_LOOP_nor_534_itm;
  reg COMP_LOOP_COMP_LOOP_and_799_itm;
  reg COMP_LOOP_COMP_LOOP_and_800_itm;
  reg COMP_LOOP_COMP_LOOP_and_801_itm;
  reg COMP_LOOP_nor_537_itm;
  reg COMP_LOOP_COMP_LOOP_and_803_itm;
  reg COMP_LOOP_COMP_LOOP_and_804_itm;
  reg COMP_LOOP_COMP_LOOP_and_805_itm;
  reg COMP_LOOP_COMP_LOOP_and_806_itm;
  reg COMP_LOOP_COMP_LOOP_and_807_itm;
  reg COMP_LOOP_COMP_LOOP_and_808_itm;
  reg COMP_LOOP_COMP_LOOP_and_809_itm;
  reg COMP_LOOP_COMP_LOOP_nor_57_itm;
  reg COMP_LOOP_nor_571_itm;
  reg COMP_LOOP_nor_572_itm;
  reg COMP_LOOP_COMP_LOOP_and_857_itm;
  reg COMP_LOOP_nor_574_itm;
  reg COMP_LOOP_COMP_LOOP_and_859_itm;
  reg COMP_LOOP_COMP_LOOP_and_860_itm;
  reg COMP_LOOP_COMP_LOOP_and_861_itm;
  reg COMP_LOOP_nor_577_itm;
  reg COMP_LOOP_COMP_LOOP_and_863_itm;
  reg COMP_LOOP_COMP_LOOP_and_864_itm;
  reg COMP_LOOP_COMP_LOOP_and_865_itm;
  reg COMP_LOOP_COMP_LOOP_and_866_itm;
  reg COMP_LOOP_COMP_LOOP_and_867_itm;
  reg COMP_LOOP_COMP_LOOP_and_868_itm;
  reg COMP_LOOP_COMP_LOOP_and_869_itm;
  reg COMP_LOOP_COMP_LOOP_nor_61_itm;
  reg COMP_LOOP_nor_611_itm;
  reg COMP_LOOP_nor_612_itm;
  reg COMP_LOOP_COMP_LOOP_and_917_itm;
  reg COMP_LOOP_nor_614_itm;
  reg COMP_LOOP_COMP_LOOP_and_919_itm;
  reg COMP_LOOP_COMP_LOOP_and_920_itm;
  reg COMP_LOOP_COMP_LOOP_and_921_itm;
  reg COMP_LOOP_nor_617_itm;
  reg COMP_LOOP_COMP_LOOP_and_923_itm;
  reg COMP_LOOP_COMP_LOOP_and_924_itm;
  reg COMP_LOOP_COMP_LOOP_and_925_itm;
  reg COMP_LOOP_COMP_LOOP_and_926_itm;
  reg COMP_LOOP_COMP_LOOP_and_927_itm;
  reg COMP_LOOP_COMP_LOOP_and_928_itm;
  reg COMP_LOOP_COMP_LOOP_and_929_itm;
  reg [5:0] COMP_LOOP_acc_psp_sva;
  reg [63:0] p_sva;
  wire mux_2240_itm;
  wire mux_2232_itm;
  wire mux_2336_itm;
  wire mux_2586_itm;
  wire mux_2688_itm;
  wire mux_2703_itm;
  wire mux_2715_itm;
  wire mux_2727_itm;
  wire mux_2734_itm;
  wire mux_2745_itm;
  wire or_tmp_2740;
  wire or_tmp_2743;
  wire mux_tmp_2749;
  wire nand_tmp_150;
  wire and_dcpl_402;
  wire [63:0] z_out;
  wire [127:0] nl_z_out;
  wire and_dcpl_418;
  wire [10:0] z_out_1;
  wire [11:0] nl_z_out_1;
  wire and_dcpl_419;
  wire and_dcpl_421;
  wire and_dcpl_423;
  wire and_dcpl_424;
  wire and_dcpl_427;
  wire and_dcpl_429;
  wire and_dcpl_431;
  wire and_dcpl_432;
  wire and_dcpl_433;
  wire and_dcpl_434;
  wire and_dcpl_435;
  wire and_dcpl_436;
  wire and_dcpl_437;
  wire and_dcpl_439;
  wire and_dcpl_440;
  wire and_dcpl_441;
  wire and_dcpl_442;
  wire and_dcpl_444;
  wire and_dcpl_445;
  wire and_dcpl_449;
  wire and_dcpl_451;
  wire and_dcpl_452;
  wire and_dcpl_453;
  wire and_dcpl_454;
  wire and_dcpl_456;
  wire and_dcpl_457;
  wire and_dcpl_458;
  wire and_dcpl_462;
  wire and_dcpl_464;
  wire and_dcpl_465;
  wire and_dcpl_466;
  wire and_dcpl_468;
  wire and_dcpl_469;
  wire and_dcpl_470;
  wire and_dcpl_471;
  wire and_dcpl_474;
  wire and_dcpl_476;
  wire and_dcpl_478;
  wire and_dcpl_481;
  wire and_dcpl_483;
  wire and_dcpl_484;
  wire and_dcpl_487;
  wire and_dcpl_489;
  wire and_dcpl_490;
  wire and_dcpl_491;
  wire and_dcpl_493;
  wire and_dcpl_495;
  wire and_dcpl_496;
  wire and_dcpl_498;
  wire [64:0] z_out_2;
  wire and_dcpl_505;
  wire and_dcpl_507;
  wire and_dcpl_508;
  wire and_dcpl_509;
  wire and_dcpl_510;
  wire and_dcpl_511;
  wire and_dcpl_523;
  wire and_dcpl_525;
  wire and_dcpl_530;
  wire and_dcpl_534;
  wire and_dcpl_543;
  wire and_dcpl_544;
  wire [63:0] z_out_3;
  wire and_dcpl_582;
  wire and_dcpl_584;
  wire and_dcpl_589;
  wire and_dcpl_593;
  wire and_dcpl_599;
  wire and_dcpl_621;
  wire [63:0] z_out_5;
  reg [63:0] r_sva;
  reg [3:0] STAGE_MAIN_LOOP_acc_1_psp_sva;
  reg [63:0] modExp_dev_result_sva;
  reg COMP_LOOP_COMP_LOOP_nor_1_itm;
  reg COMP_LOOP_nor_12_itm;
  reg COMP_LOOP_nor_14_itm;
  reg COMP_LOOP_COMP_LOOP_and_19_itm;
  reg COMP_LOOP_COMP_LOOP_and_20_itm;
  reg COMP_LOOP_COMP_LOOP_and_21_itm;
  reg COMP_LOOP_nor_17_itm;
  reg COMP_LOOP_COMP_LOOP_and_23_itm;
  reg COMP_LOOP_COMP_LOOP_and_24_itm;
  reg COMP_LOOP_COMP_LOOP_and_25_itm;
  reg COMP_LOOP_COMP_LOOP_and_26_itm;
  reg COMP_LOOP_COMP_LOOP_and_27_itm;
  reg COMP_LOOP_COMP_LOOP_and_28_itm;
  reg COMP_LOOP_COMP_LOOP_and_29_itm;
  reg [54:0] modExp_dev_exp_1_sva_63_9;
  reg [4:0] modExp_dev_exp_1_sva_8_4;
  wire [9:0] STAGE_MAIN_LOOP_lshift_psp_1_sva_mx0w0;
  wire COMP_LOOP_10_modExp_dev_1_while_mul_mut_mx0c4;
  wire COMP_LOOP_10_modExp_dev_1_while_mul_mut_mx0c5;
  wire STAGE_VEC_LOOP_j_sva_9_0_mx0c1;
  wire COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c3;
  wire COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c4;
  wire COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c5;
  wire COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c6;
  wire COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c7;
  wire COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c8;
  wire COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c9;
  wire COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c10;
  wire COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c11;
  wire COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c12;
  wire COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c13;
  wire operator_64_false_slc_operator_64_false_acc_1_60_itm_mx0c1;
  wire operator_64_false_slc_operator_64_false_acc_1_60_itm_mx0c2;
  wire operator_64_false_slc_operator_64_false_acc_1_60_itm_mx0c3;
  wire operator_64_false_slc_operator_64_false_acc_1_60_itm_mx0c4;
  wire tmp_1_lpi_4_dfm_mx0c0;
  wire and_330_rgt;
  wire or_2938_cse;
  wire nor_554_cse;
  wire or_2955_cse;
  wire mux_2332_cse;
  wire mux_2326_cse;
  wire or_2929_cse;
  wire mux_2829_cse;
  wire nand_176_cse;
  wire mux_2830_cse;
  wire and_920_cse;
  wire and_936_cse;
  wire and_945_cse;
  wire and_950_cse;
  wire and_953_cse;
  wire and_957_cse;
  wire and_964_cse;
  wire and_966_cse;
  wire and_973_cse;
  wire and_975_cse;
  wire and_978_cse;
  wire mux_2835_cse;
  wire or_2960_cse;
  wire and_925_cse;
  wire and_940_cse;
  wire and_960_cse;
  wire and_970_cse;
  wire mux_tmp_2812;
  wire mux_tmp_2813;
  wire mux_tmp_2815;
  wire mux_tmp_2823;
  wire mux_tmp_2824;
  wire nand_490_cse;
  wire nor_1040_cse;
  wire or_3018_cse;
  wire nor_1039_cse;
  wire and_694_cse;
  wire mux_2797_itm;
  wire mux_2545_itm;
  wire mux_2863_itm;
  wire operator_64_false_or_120_itm;
  wire operator_64_false_or_121_cse;
  wire operator_64_false_operator_64_false_or_1_cse;
  wire [11:0] COMP_LOOP_slc_acc_3_12_1_slc;

  wire[0:0] mux_2239_nl;
  wire[0:0] mux_2238_nl;
  wire[0:0] mux_2237_nl;
  wire[0:0] mux_2236_nl;
  wire[0:0] mux_2235_nl;
  wire[0:0] mux_2234_nl;
  wire[0:0] mux_2233_nl;
  wire[0:0] mux_2231_nl;
  wire[0:0] mux_2230_nl;
  wire[0:0] mux_2229_nl;
  wire[0:0] mux_2228_nl;
  wire[0:0] mux_2227_nl;
  wire[0:0] mux_2226_nl;
  wire[0:0] mux_2225_nl;
  wire[0:0] mux_2224_nl;
  wire[0:0] mux_2223_nl;
  wire[0:0] mux_2222_nl;
  wire[0:0] mux_2221_nl;
  wire[0:0] mux_2220_nl;
  wire[0:0] mux_2219_nl;
  wire[0:0] mux_2218_nl;
  wire[0:0] mux_2217_nl;
  wire[0:0] mux_2216_nl;
  wire[0:0] mux_2215_nl;
  wire[0:0] mux_2214_nl;
  wire[0:0] mux_2213_nl;
  wire[0:0] mux_2211_nl;
  wire[0:0] mux_2210_nl;
  wire[0:0] mux_2209_nl;
  wire[0:0] mux_2208_nl;
  wire[0:0] or_2841_nl;
  wire[0:0] mux_2207_nl;
  wire[0:0] mux_2206_nl;
  wire[0:0] mux_2205_nl;
  wire[0:0] mux_2204_nl;
  wire[0:0] mux_2203_nl;
  wire[0:0] mux_2202_nl;
  wire[0:0] mux_2201_nl;
  wire[0:0] mux_2200_nl;
  wire[0:0] or_2392_nl;
  wire[0:0] mux_2199_nl;
  wire[0:0] mux_2198_nl;
  wire[0:0] mux_2197_nl;
  wire[0:0] mux_2196_nl;
  wire[0:0] mux_2195_nl;
  wire[0:0] mux_2194_nl;
  wire[0:0] mux_2192_nl;
  wire[0:0] mux_2191_nl;
  wire[0:0] mux_2189_nl;
  wire[0:0] mux_2188_nl;
  wire[0:0] mux_2187_nl;
  wire[0:0] mux_2185_nl;
  wire[0:0] mux_2184_nl;
  wire[0:0] mux_2179_nl;
  wire[0:0] mux_2173_nl;
  wire[0:0] mux_2172_nl;
  wire[0:0] mux_2171_nl;
  wire[0:0] mux_2170_nl;
  wire[0:0] mux_2168_nl;
  wire[0:0] mux_2167_nl;
  wire[0:0] mux_2166_nl;
  wire[0:0] mux_2323_nl;
  wire[0:0] mux_2322_nl;
  wire[0:0] mux_2321_nl;
  wire[0:0] mux_2320_nl;
  wire[0:0] mux_2319_nl;
  wire[0:0] mux_2318_nl;
  wire[0:0] or_2479_nl;
  wire[0:0] mux_2317_nl;
  wire[0:0] mux_2316_nl;
  wire[0:0] mux_2315_nl;
  wire[0:0] mux_2314_nl;
  wire[0:0] nand_177_nl;
  wire[0:0] mux_2313_nl;
  wire[0:0] or_2477_nl;
  wire[0:0] mux_2312_nl;
  wire[0:0] mux_2311_nl;
  wire[0:0] mux_2310_nl;
  wire[0:0] or_2476_nl;
  wire[0:0] mux_2309_nl;
  wire[0:0] nand_178_nl;
  wire[0:0] mux_2308_nl;
  wire[0:0] mux_2307_nl;
  wire[0:0] mux_2306_nl;
  wire[0:0] mux_2305_nl;
  wire[0:0] mux_2304_nl;
  wire[0:0] mux_2303_nl;
  wire[0:0] mux_2302_nl;
  wire[0:0] mux_2300_nl;
  wire[0:0] mux_2299_nl;
  wire[0:0] or_2468_nl;
  wire[0:0] mux_2297_nl;
  wire[0:0] mux_2296_nl;
  wire[0:0] or_2461_nl;
  wire[0:0] mux_2294_nl;
  wire[0:0] mux_2293_nl;
  wire[0:0] mux_2292_nl;
  wire[0:0] or_2455_nl;
  wire[0:0] mux_2339_nl;
  wire[0:0] mux_2338_nl;
  wire[0:0] mux_2337_nl;
  wire[0:0] nor_549_nl;
  wire[0:0] and_511_nl;
  wire[0:0] and_512_nl;
  wire[0:0] and_513_nl;
  wire[0:0] mux_1016_nl;
  wire[0:0] nor_548_nl;
  wire[0:0] operator_64_false_or_2_nl;
  wire[0:0] mux_2427_nl;
  wire[0:0] nor_524_nl;
  wire[0:0] and_331_nl;
  wire[0:0] COMP_LOOP_or_2_nl;
  wire[0:0] COMP_LOOP_or_3_nl;
  wire[0:0] COMP_LOOP_or_4_nl;
  wire[0:0] COMP_LOOP_or_5_nl;
  wire[0:0] COMP_LOOP_or_6_nl;
  wire[0:0] COMP_LOOP_or_7_nl;
  wire[0:0] COMP_LOOP_or_8_nl;
  wire[0:0] COMP_LOOP_or_9_nl;
  wire[0:0] COMP_LOOP_or_10_nl;
  wire[0:0] COMP_LOOP_or_11_nl;
  wire[0:0] COMP_LOOP_or_12_nl;
  wire[0:0] COMP_LOOP_or_13_nl;
  wire[0:0] COMP_LOOP_or_14_nl;
  wire[0:0] COMP_LOOP_or_15_nl;
  wire[0:0] COMP_LOOP_or_16_nl;
  wire[0:0] COMP_LOOP_or_17_nl;
  wire[0:0] mux_2475_nl;
  wire[0:0] mux_2474_nl;
  wire[0:0] mux_2473_nl;
  wire[0:0] mux_2472_nl;
  wire[0:0] mux_2471_nl;
  wire[0:0] mux_2470_nl;
  wire[0:0] or_2623_nl;
  wire[0:0] mux_2469_nl;
  wire[0:0] or_2622_nl;
  wire[0:0] mux_2468_nl;
  wire[0:0] mux_2467_nl;
  wire[0:0] mux_2466_nl;
  wire[0:0] mux_2465_nl;
  wire[0:0] mux_2464_nl;
  wire[0:0] mux_2463_nl;
  wire[0:0] mux_2462_nl;
  wire[0:0] mux_2461_nl;
  wire[0:0] mux_2460_nl;
  wire[0:0] mux_2459_nl;
  wire[0:0] mux_2458_nl;
  wire[0:0] or_2621_nl;
  wire[0:0] mux_2457_nl;
  wire[0:0] mux_2456_nl;
  wire[0:0] mux_2455_nl;
  wire[0:0] mux_2454_nl;
  wire[0:0] mux_2453_nl;
  wire[0:0] mux_2452_nl;
  wire[0:0] mux_2450_nl;
  wire[0:0] mux_2449_nl;
  wire[0:0] mux_2448_nl;
  wire[0:0] mux_2447_nl;
  wire[0:0] mux_2446_nl;
  wire[0:0] mux_2445_nl;
  wire[0:0] mux_2444_nl;
  wire[0:0] mux_2443_nl;
  wire[0:0] mux_2442_nl;
  wire[0:0] mux_2441_nl;
  wire[0:0] mux_2437_nl;
  wire[0:0] mux_2436_nl;
  wire[0:0] mux_2435_nl;
  wire[0:0] mux_2434_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_17_nl;
  wire[0:0] modExp_dev_while_or_nl;
  wire[0:0] modExp_dev_while_or_1_nl;
  wire[0:0] nand_486_nl;
  wire[0:0] mux_2864_nl;
  wire[0:0] nor_nl;
  wire[0:0] nor_1038_nl;
  wire[3:0] operator_64_false_or_2_nl_1;
  wire[3:0] operator_64_false_and_nl;
  wire[3:0] operator_64_false_mux1h_nl;
  wire[0:0] and_421_nl;
  wire[0:0] and_422_nl;
  wire[0:0] and_423_nl;
  wire[0:0] and_424_nl;
  wire[0:0] and_425_nl;
  wire[0:0] and_426_nl;
  wire[0:0] and_427_nl;
  wire[0:0] and_428_nl;
  wire[0:0] and_429_nl;
  wire[0:0] and_430_nl;
  wire[0:0] and_431_nl;
  wire[0:0] and_432_nl;
  wire[0:0] and_433_nl;
  wire[0:0] and_434_nl;
  wire[0:0] COMP_LOOP_nand_nl;
  wire[0:0] and_435_nl;
  wire[5:0] operator_64_false_1_acc_nl;
  wire[6:0] nl_operator_64_false_1_acc_nl;
  wire[0:0] mux_2590_nl;
  wire[0:0] or_2696_nl;
  wire[0:0] mux_2587_nl;
  wire[0:0] mux_2592_nl;
  wire[0:0] mux_2591_nl;
  wire[0:0] or_2699_nl;
  wire[0:0] mux_2599_nl;
  wire[0:0] mux_2598_nl;
  wire[0:0] mux_2597_nl;
  wire[0:0] mux_2596_nl;
  wire[0:0] mux_2594_nl;
  wire[0:0] mux_2593_nl;
  wire[0:0] mux_2601_nl;
  wire[0:0] mux_2600_nl;
  wire[0:0] or_2701_nl;
  wire[0:0] mux_2612_nl;
  wire[0:0] mux_2611_nl;
  wire[0:0] and_485_nl;
  wire[0:0] mux_2616_nl;
  wire[0:0] or_2824_nl;
  wire[0:0] mux_2615_nl;
  wire[0:0] mux_2614_nl;
  wire[0:0] or_2825_nl;
  wire[0:0] nand_161_nl;
  wire[0:0] nand_162_nl;
  wire[0:0] mux_2621_nl;
  wire[0:0] or_2707_nl;
  wire[0:0] mux_2620_nl;
  wire[0:0] mux_2619_nl;
  wire[0:0] and_482_nl;
  wire[0:0] mux_2624_nl;
  wire[0:0] or_2708_nl;
  wire[0:0] mux_2623_nl;
  wire[0:0] and_480_nl;
  wire[0:0] mux_2633_nl;
  wire[0:0] mux_2632_nl;
  wire[0:0] mux_2631_nl;
  wire[0:0] mux_2630_nl;
  wire[0:0] mux_2629_nl;
  wire[0:0] mux_2628_nl;
  wire[0:0] mux_2627_nl;
  wire[0:0] mux_2626_nl;
  wire[0:0] mux_2640_nl;
  wire[0:0] mux_2639_nl;
  wire[0:0] mux_2638_nl;
  wire[0:0] mux_2637_nl;
  wire[0:0] nor_511_nl;
  wire[0:0] and_473_nl;
  wire[0:0] mux_2641_nl;
  wire[0:0] and_393_nl;
  wire[0:0] mux_2645_nl;
  wire[0:0] and_397_nl;
  wire[0:0] mux_2649_nl;
  wire[0:0] mux_2648_nl;
  wire[0:0] mux_2647_nl;
  wire[0:0] mux_2646_nl;
  wire[0:0] nor_937_nl;
  wire[0:0] and_754_nl;
  wire[0:0] and_755_nl;
  wire[0:0] mux_2657_nl;
  wire[0:0] mux_2656_nl;
  wire[0:0] mux_2655_nl;
  wire[0:0] or_196_nl;
  wire[0:0] mux_2654_nl;
  wire[0:0] mux_2653_nl;
  wire[0:0] or_2651_nl;
  wire[0:0] or_2732_nl;
  wire[0:0] mux_2670_nl;
  wire[0:0] mux_2669_nl;
  wire[0:0] mux_2668_nl;
  wire[0:0] mux_2667_nl;
  wire[0:0] mux_2666_nl;
  wire[0:0] mux_2681_nl;
  wire[0:0] mux_2680_nl;
  wire[0:0] mux_2679_nl;
  wire[0:0] mux_2678_nl;
  wire[0:0] or_2743_nl;
  wire[0:0] or_2748_nl;
  wire[0:0] mux_2692_nl;
  wire[0:0] mux_2691_nl;
  wire[0:0] nor_503_nl;
  wire[0:0] mux_2690_nl;
  wire[0:0] nor_504_nl;
  wire[0:0] and_409_nl;
  wire[0:0] mux_2708_nl;
  wire[0:0] mux_2707_nl;
  wire[0:0] mux_2706_nl;
  wire[0:0] nor_500_nl;
  wire[0:0] and_452_nl;
  wire[0:0] mux_2705_nl;
  wire[0:0] or_2755_nl;
  wire[0:0] mux_2713_nl;
  wire[0:0] mux_2712_nl;
  wire[0:0] mux_2711_nl;
  wire[0:0] nor_498_nl;
  wire[0:0] mux_2710_nl;
  wire[0:0] nor_499_nl;
  wire[0:0] and_410_nl;
  wire[0:0] mux_2722_nl;
  wire[0:0] mux_2721_nl;
  wire[0:0] mux_2720_nl;
  wire[0:0] mux_2719_nl;
  wire[0:0] mux_2718_nl;
  wire[0:0] and_636_nl;
  wire[0:0] mux_2730_nl;
  wire[0:0] mux_2729_nl;
  wire[0:0] or_2814_nl;
  wire[0:0] mux_2728_nl;
  wire[0:0] or_2815_nl;
  wire[0:0] nand_156_nl;
  wire[0:0] mux_2733_nl;
  wire[0:0] mux_2732_nl;
  wire[0:0] or_2812_nl;
  wire[0:0] mux_2731_nl;
  wire[0:0] or_411_nl;
  wire[0:0] or_2777_nl;
  wire[0:0] nand_154_nl;
  wire[0:0] and_413_nl;
  wire[0:0] and_414_nl;
  wire[0:0] mux_2736_nl;
  wire[0:0] or_2891_nl;
  wire[0:0] COMP_LOOP_nor_11_nl;
  wire[0:0] COMP_LOOP_or_35_nl;
  wire[0:0] COMP_LOOP_or_18_nl;
  wire[0:0] COMP_LOOP_or_19_nl;
  wire[0:0] COMP_LOOP_or_20_nl;
  wire[0:0] COMP_LOOP_or_21_nl;
  wire[0:0] COMP_LOOP_or_22_nl;
  wire[0:0] COMP_LOOP_or_23_nl;
  wire[0:0] COMP_LOOP_or_24_nl;
  wire[0:0] COMP_LOOP_or_25_nl;
  wire[0:0] COMP_LOOP_or_26_nl;
  wire[0:0] COMP_LOOP_or_27_nl;
  wire[0:0] COMP_LOOP_or_28_nl;
  wire[0:0] COMP_LOOP_or_29_nl;
  wire[0:0] COMP_LOOP_or_30_nl;
  wire[0:0] COMP_LOOP_or_31_nl;
  wire[0:0] COMP_LOOP_or_32_nl;
  wire[0:0] COMP_LOOP_or_33_nl;
  wire[0:0] not_7089_nl;
  wire[0:0] mux_2893_nl;
  wire[0:0] mux_2892_nl;
  wire[0:0] nand_nl;
  wire[0:0] mux_2891_nl;
  wire[0:0] mux_2890_nl;
  wire[0:0] nor_1035_nl;
  wire[0:0] mux_2889_nl;
  wire[0:0] mux_2896_nl;
  wire[0:0] or_3019_nl;
  wire[0:0] mux_2888_nl;
  wire[0:0] mux_2887_nl;
  wire[0:0] mux_2895_nl;
  wire[0:0] mux_2885_nl;
  wire[0:0] or_3017_nl;
  wire[0:0] mux_2884_nl;
  wire[0:0] mux_2883_nl;
  wire[0:0] mux_2882_nl;
  wire[0:0] mux_2881_nl;
  wire[0:0] mux_2880_nl;
  wire[0:0] mux_2879_nl;
  wire[0:0] mux_2878_nl;
  wire[0:0] mux_2875_nl;
  wire[0:0] mux_2874_nl;
  wire[0:0] or_3011_nl;
  wire[0:0] mux_2873_nl;
  wire[0:0] or_3008_nl;
  wire[0:0] mux_2872_nl;
  wire[0:0] mux_2871_nl;
  wire[0:0] mux_2870_nl;
  wire[0:0] mux_2869_nl;
  wire[0:0] or_3006_nl;
  wire[0:0] mux_2867_nl;
  wire[0:0] or_3005_nl;
  wire[0:0] or_3004_nl;
  wire[0:0] or_424_nl;
  wire[0:0] or_444_nl;
  wire[0:0] or_533_nl;
  wire[0:0] mux_1049_nl;
  wire[0:0] mux_1048_nl;
  wire[0:0] or_2836_nl;
  wire[0:0] nand_389_nl;
  wire[0:0] nand_390_nl;
  wire[0:0] nand_391_nl;
  wire[0:0] nor_809_nl;
  wire[0:0] nor_810_nl;
  wire[0:0] and_741_nl;
  wire[0:0] nor_797_nl;
  wire[0:0] mux_1085_nl;
  wire[0:0] nor_775_nl;
  wire[0:0] nor_776_nl;
  wire[0:0] mux_1111_nl;
  wire[0:0] or_735_nl;
  wire[0:0] mux_1153_nl;
  wire[0:0] nor_763_nl;
  wire[0:0] nor_764_nl;
  wire[0:0] mux_1221_nl;
  wire[0:0] nor_751_nl;
  wire[0:0] nor_752_nl;
  wire[0:0] mux_1289_nl;
  wire[0:0] nor_739_nl;
  wire[0:0] nor_740_nl;
  wire[0:0] mux_1357_nl;
  wire[0:0] nor_727_nl;
  wire[0:0] nor_728_nl;
  wire[0:0] mux_1425_nl;
  wire[0:0] nor_715_nl;
  wire[0:0] nor_716_nl;
  wire[0:0] mux_1493_nl;
  wire[0:0] nor_703_nl;
  wire[0:0] nor_704_nl;
  wire[0:0] mux_1561_nl;
  wire[0:0] nor_691_nl;
  wire[0:0] nor_692_nl;
  wire[0:0] mux_1629_nl;
  wire[0:0] nor_679_nl;
  wire[0:0] nor_680_nl;
  wire[0:0] mux_1697_nl;
  wire[0:0] nor_667_nl;
  wire[0:0] nor_668_nl;
  wire[0:0] mux_1765_nl;
  wire[0:0] nor_655_nl;
  wire[0:0] nor_656_nl;
  wire[0:0] mux_1833_nl;
  wire[0:0] nor_643_nl;
  wire[0:0] nor_644_nl;
  wire[0:0] mux_1901_nl;
  wire[0:0] nor_631_nl;
  wire[0:0] nor_632_nl;
  wire[0:0] mux_1969_nl;
  wire[0:0] nor_619_nl;
  wire[0:0] nor_620_nl;
  wire[0:0] mux_2037_nl;
  wire[0:0] nor_607_nl;
  wire[0:0] nor_608_nl;
  wire[0:0] mux_2105_nl;
  wire[0:0] nor_595_nl;
  wire[0:0] nor_596_nl;
  wire[0:0] or_2390_nl;
  wire[0:0] mux_2174_nl;
  wire[0:0] mux_2177_nl;
  wire[0:0] mux_2176_nl;
  wire[0:0] or_2412_nl;
  wire[0:0] or_2411_nl;
  wire[0:0] or_2634_nl;
  wire[0:0] or_2431_nl;
  wire[0:0] nand_180_nl;
  wire[0:0] or_2464_nl;
  wire[0:0] or_2462_nl;
  wire[0:0] nor_552_nl;
  wire[0:0] or_2486_nl;
  wire[0:0] or_2484_nl;
  wire[0:0] nor_550_nl;
  wire[0:0] nor_551_nl;
  wire[0:0] mux_2335_nl;
  wire[0:0] or_2498_nl;
  wire[0:0] mux_2334_nl;
  wire[0:0] or_2497_nl;
  wire[0:0] or_2495_nl;
  wire[0:0] mux_2333_nl;
  wire[0:0] nand_120_nl;
  wire[0:0] or_2492_nl;
  wire[0:0] mux_2331_nl;
  wire[0:0] or_2491_nl;
  wire[0:0] mux_2330_nl;
  wire[0:0] mux_2329_nl;
  wire[0:0] mux_2328_nl;
  wire[0:0] or_2489_nl;
  wire[0:0] or_2488_nl;
  wire[0:0] mux_2325_nl;
  wire[0:0] nand_175_nl;
  wire[0:0] mux_2324_nl;
  wire[0:0] or_2482_nl;
  wire[0:0] or_2480_nl;
  wire[0:0] mux_2358_nl;
  wire[0:0] mux_2357_nl;
  wire[0:0] nor_541_nl;
  wire[0:0] nor_542_nl;
  wire[0:0] mux_2356_nl;
  wire[0:0] and_506_nl;
  wire[0:0] mux_2355_nl;
  wire[0:0] or_2521_nl;
  wire[0:0] mux_2354_nl;
  wire[0:0] nor_825_nl;
  wire[0:0] nor_544_nl;
  wire[0:0] mux_2353_nl;
  wire[0:0] or_2518_nl;
  wire[0:0] mux_2352_nl;
  wire[0:0] mux_2351_nl;
  wire[0:0] nor_545_nl;
  wire[0:0] mux_2350_nl;
  wire[0:0] or_2831_nl;
  wire[0:0] and_507_nl;
  wire[0:0] mux_2348_nl;
  wire[0:0] or_2510_nl;
  wire[0:0] and_508_nl;
  wire[0:0] mux_2347_nl;
  wire[0:0] nor_546_nl;
  wire[0:0] nor_547_nl;
  wire[0:0] or_2555_nl;
  wire[0:0] nand_420_nl;
  wire[0:0] or_2612_nl;
  wire[0:0] mux_2439_nl;
  wire[0:0] mux_2438_nl;
  wire[0:0] mux_2511_nl;
  wire[0:0] mux_2507_nl;
  wire[0:0] nand_137_nl;
  wire[0:0] mux_2524_nl;
  wire[0:0] mux_2531_nl;
  wire[0:0] and_494_nl;
  wire[0:0] nor_516_nl;
  wire[0:0] and_489_nl;
  wire[0:0] mux_2585_nl;
  wire[0:0] mux_2584_nl;
  wire[0:0] mux_2583_nl;
  wire[0:0] mux_2582_nl;
  wire[0:0] mux_2581_nl;
  wire[0:0] mux_2610_nl;
  wire[0:0] mux_2609_nl;
  wire[0:0] mux_2608_nl;
  wire[0:0] mux_2607_nl;
  wire[0:0] mux_2606_nl;
  wire[0:0] or_2877_nl;
  wire[0:0] mux_2605_nl;
  wire[0:0] mux_2604_nl;
  wire[0:0] mux_2603_nl;
  wire[0:0] mux_2602_nl;
  wire[0:0] or_2604_nl;
  wire[0:0] mux_2613_nl;
  wire[0:0] mux_2618_nl;
  wire[0:0] mux_2617_nl;
  wire[0:0] and_483_nl;
  wire[0:0] mux_2622_nl;
  wire[0:0] nor_871_nl;
  wire[0:0] and_684_nl;
  wire[0:0] mux_2636_nl;
  wire[0:0] or_2712_nl;
  wire[0:0] mux_2635_nl;
  wire[0:0] mux_2644_nl;
  wire[0:0] nor_940_nl;
  wire[0:0] mux_2643_nl;
  wire[0:0] or_2719_nl;
  wire[0:0] or_2900_nl;
  wire[0:0] mux_2642_nl;
  wire[0:0] and_395_nl;
  wire[0:0] mux_2651_nl;
  wire[0:0] and_400_nl;
  wire[0:0] mux_2650_nl;
  wire[0:0] mux_2661_nl;
  wire[0:0] and_403_nl;
  wire[0:0] mux_2660_nl;
  wire[0:0] mux_2659_nl;
  wire[0:0] mux_2664_nl;
  wire[0:0] mux_2674_nl;
  wire[0:0] or_2740_nl;
  wire[0:0] mux_2673_nl;
  wire[0:0] or_2737_nl;
  wire[0:0] mux_2672_nl;
  wire[0:0] or_2735_nl;
  wire[0:0] mux_2687_nl;
  wire[0:0] mux_2686_nl;
  wire[0:0] mux_2685_nl;
  wire[0:0] or_2747_nl;
  wire[0:0] mux_2684_nl;
  wire[0:0] and_461_nl;
  wire[0:0] mux_2702_nl;
  wire[0:0] mux_2701_nl;
  wire[0:0] mux_2700_nl;
  wire[0:0] mux_2699_nl;
  wire[0:0] mux_2698_nl;
  wire[0:0] mux_2697_nl;
  wire[0:0] mux_2696_nl;
  wire[0:0] mux_2695_nl;
  wire[0:0] or_2762_nl;
  wire[0:0] mux_2726_nl;
  wire[0:0] mux_2725_nl;
  wire[0:0] mux_2724_nl;
  wire[0:0] nor_494_nl;
  wire[0:0] and_444_nl;
  wire[0:0] and_445_nl;
  wire[0:0] and_412_nl;
  wire[0:0] mux_2739_nl;
  wire[0:0] mux_2744_nl;
  wire[0:0] mux_2743_nl;
  wire[0:0] mux_2742_nl;
  wire[0:0] mux_2741_nl;
  wire[0:0] nor_490_nl;
  wire[0:0] mux_2763_nl;
  wire[0:0] mux_2762_nl;
  wire[0:0] nand_145_nl;
  wire[0:0] mux_2783_nl;
  wire[0:0] mux_2782_nl;
  wire[0:0] mux_2796_nl;
  wire[0:0] mux_2795_nl;
  wire[0:0] mux_2794_nl;
  wire[0:0] mux_2793_nl;
  wire[0:0] mux_2792_nl;
  wire[0:0] mux_2791_nl;
  wire[0:0] mux_2790_nl;
  wire[0:0] mux_2789_nl;
  wire[0:0] mux_2788_nl;
  wire[0:0] mux_2787_nl;
  wire[0:0] mux_2786_nl;
  wire[0:0] mux_2785_nl;
  wire[0:0] mux_2784_nl;
  wire[0:0] mux_2781_nl;
  wire[0:0] nand_147_nl;
  wire[0:0] mux_2780_nl;
  wire[0:0] mux_2779_nl;
  wire[0:0] mux_2778_nl;
  wire[0:0] mux_2777_nl;
  wire[0:0] mux_2776_nl;
  wire[0:0] nand_146_nl;
  wire[0:0] mux_2774_nl;
  wire[0:0] mux_2773_nl;
  wire[0:0] mux_2770_nl;
  wire[0:0] mux_2769_nl;
  wire[0:0] mux_2768_nl;
  wire[0:0] nor_489_nl;
  wire[0:0] mux_2767_nl;
  wire[0:0] mux_2371_nl;
  wire[0:0] mux_2370_nl;
  wire[0:0] and_504_nl;
  wire[0:0] nor_534_nl;
  wire[0:0] mux_2369_nl;
  wire[0:0] or_2547_nl;
  wire[0:0] nand_126_nl;
  wire[0:0] and_505_nl;
  wire[0:0] mux_2367_nl;
  wire[0:0] nor_535_nl;
  wire[0:0] nor_536_nl;
  wire[0:0] mux_2366_nl;
  wire[0:0] nor_537_nl;
  wire[0:0] mux_2365_nl;
  wire[0:0] or_2539_nl;
  wire[0:0] mux_2364_nl;
  wire[0:0] mux_2362_nl;
  wire[0:0] nor_538_nl;
  wire[0:0] mux_2361_nl;
  wire[0:0] or_2531_nl;
  wire[0:0] or_2530_nl;
  wire[0:0] mux_2360_nl;
  wire[0:0] nor_539_nl;
  wire[0:0] nor_540_nl;
  wire[0:0] mux_2385_nl;
  wire[0:0] mux_2384_nl;
  wire[0:0] nor_525_nl;
  wire[0:0] mux_2383_nl;
  wire[0:0] mux_2382_nl;
  wire[0:0] or_2571_nl;
  wire[0:0] or_2625_nl;
  wire[0:0] nand_172_nl;
  wire[0:0] and_501_nl;
  wire[0:0] mux_2381_nl;
  wire[0:0] nor_526_nl;
  wire[0:0] nor_527_nl;
  wire[0:0] mux_2380_nl;
  wire[0:0] nor_528_nl;
  wire[0:0] and_502_nl;
  wire[0:0] mux_2379_nl;
  wire[0:0] or_2560_nl;
  wire[0:0] mux_2378_nl;
  wire[0:0] mux_2377_nl;
  wire[0:0] and_503_nl;
  wire[0:0] mux_2376_nl;
  wire[0:0] nor_529_nl;
  wire[0:0] nor_530_nl;
  wire[0:0] mux_2375_nl;
  wire[0:0] nor_532_nl;
  wire[0:0] nor_533_nl;
  wire[0:0] mux_2373_nl;
  wire[0:0] or_2550_nl;
  wire[0:0] mux_2544_nl;
  wire[0:0] mux_2543_nl;
  wire[0:0] mux_2542_nl;
  wire[0:0] mux_2541_nl;
  wire[0:0] or_2664_nl;
  wire[0:0] mux_2540_nl;
  wire[0:0] mux_2539_nl;
  wire[0:0] mux_2538_nl;
  wire[0:0] mux_2537_nl;
  wire[0:0] mux_2536_nl;
  wire[0:0] mux_2535_nl;
  wire[0:0] mux_2534_nl;
  wire[0:0] mux_2533_nl;
  wire[0:0] mux_2532_nl;
  wire[0:0] mux_2530_nl;
  wire[0:0] nand_139_nl;
  wire[0:0] mux_2529_nl;
  wire[0:0] mux_2528_nl;
  wire[0:0] mux_2527_nl;
  wire[0:0] mux_2526_nl;
  wire[0:0] nand_138_nl;
  wire[0:0] mux_2523_nl;
  wire[0:0] mux_2522_nl;
  wire[0:0] mux_2517_nl;
  wire[0:0] mux_2516_nl;
  wire[0:0] mux_2515_nl;
  wire[0:0] nor_520_nl;
  wire[0:0] mux_2514_nl;
  wire[0:0] and_125_nl;
  wire[0:0] mux_1051_nl;
  wire[0:0] or_508_nl;
  wire[0:0] and_132_nl;
  wire[0:0] and_136_nl;
  wire[0:0] and_139_nl;
  wire[0:0] mux_1052_nl;
  wire[0:0] nor_811_nl;
  wire[0:0] nor_812_nl;
  wire[0:0] and_144_nl;
  wire[0:0] and_149_nl;
  wire[0:0] mux_1054_nl;
  wire[0:0] and_556_nl;
  wire[0:0] nor_808_nl;
  wire[0:0] and_151_nl;
  wire[0:0] mux_1055_nl;
  wire[0:0] nor_806_nl;
  wire[0:0] nor_807_nl;
  wire[0:0] and_156_nl;
  wire[0:0] mux_1056_nl;
  wire[0:0] nor_804_nl;
  wire[0:0] nor_805_nl;
  wire[0:0] and_159_nl;
  wire[0:0] mux_1057_nl;
  wire[0:0] nor_802_nl;
  wire[0:0] nor_803_nl;
  wire[0:0] and_163_nl;
  wire[0:0] mux_1058_nl;
  wire[0:0] and_555_nl;
  wire[0:0] nor_801_nl;
  wire[0:0] and_171_nl;
  wire[0:0] and_175_nl;
  wire[0:0] mux_1059_nl;
  wire[0:0] nor_799_nl;
  wire[0:0] nor_800_nl;
  wire[0:0] and_179_nl;
  wire[0:0] mux_1060_nl;
  wire[0:0] nor_798_nl;
  wire[0:0] and_554_nl;
  wire[0:0] and_184_nl;
  wire[0:0] and_188_nl;
  wire[0:0] and_191_nl;
  wire[0:0] mux_1062_nl;
  wire[0:0] nor_795_nl;
  wire[0:0] nor_796_nl;
  wire[0:0] and_196_nl;
  wire[0:0] mux_1063_nl;
  wire[0:0] nor_793_nl;
  wire[0:0] nor_794_nl;
  wire[0:0] and_200_nl;
  wire[0:0] mux_1064_nl;
  wire[0:0] and_552_nl;
  wire[0:0] nor_792_nl;
  wire[0:0] and_205_nl;
  wire[0:0] mux_1065_nl;
  wire[0:0] nor_790_nl;
  wire[0:0] nor_791_nl;
  wire[0:0] and_208_nl;
  wire[0:0] mux_1066_nl;
  wire[0:0] nor_788_nl;
  wire[0:0] nor_789_nl;
  wire[0:0] and_213_nl;
  wire[0:0] and_218_nl;
  wire[0:0] and_223_nl;
  wire[0:0] and_227_nl;
  wire[0:0] mux_1067_nl;
  wire[0:0] nor_786_nl;
  wire[0:0] and_762_nl;
  wire[0:0] and_231_nl;
  wire[0:0] mux_1068_nl;
  wire[0:0] and_551_nl;
  wire[0:0] nor_785_nl;
  wire[0:0] and_234_nl;
  wire[0:0] mux_1069_nl;
  wire[0:0] and_237_nl;
  wire[0:0] mux_1070_nl;
  wire[0:0] and_550_nl;
  wire[0:0] nor_784_nl;
  wire[0:0] and_240_nl;
  wire[0:0] mux_1071_nl;
  wire[0:0] nor_782_nl;
  wire[0:0] nor_783_nl;
  wire[0:0] and_245_nl;
  wire[0:0] mux_1072_nl;
  wire[0:0] nor_781_nl;
  wire[0:0] and_549_nl;
  wire[0:0] and_249_nl;
  wire[0:0] mux_1073_nl;
  wire[0:0] nor_779_nl;
  wire[0:0] nor_780_nl;
  wire[0:0] and_250_nl;
  wire[0:0] and_254_nl;
  wire[0:0] mux_1074_nl;
  wire[0:0] nor_777_nl;
  wire[0:0] nor_778_nl;
  wire[0:0] mux_1107_nl;
  wire[0:0] mux_1106_nl;
  wire[0:0] mux_1105_nl;
  wire[0:0] nand_18_nl;
  wire[0:0] mux_1104_nl;
  wire[0:0] mux_1103_nl;
  wire[0:0] nor_765_nl;
  wire[0:0] nor_766_nl;
  wire[0:0] mux_1102_nl;
  wire[0:0] nor_767_nl;
  wire[0:0] nor_768_nl;
  wire[0:0] mux_1101_nl;
  wire[0:0] nand_17_nl;
  wire[0:0] mux_1100_nl;
  wire[0:0] nor_769_nl;
  wire[0:0] nor_770_nl;
  wire[0:0] mux_1099_nl;
  wire[0:0] mux_1098_nl;
  wire[0:0] or_711_nl;
  wire[0:0] or_709_nl;
  wire[0:0] or_708_nl;
  wire[0:0] mux_1097_nl;
  wire[0:0] or_707_nl;
  wire[0:0] mux_1096_nl;
  wire[0:0] mux_1095_nl;
  wire[0:0] or_706_nl;
  wire[0:0] or_705_nl;
  wire[0:0] mux_1094_nl;
  wire[0:0] or_703_nl;
  wire[0:0] or_701_nl;
  wire[0:0] mux_1093_nl;
  wire[0:0] or_699_nl;
  wire[0:0] mux_1092_nl;
  wire[0:0] or_698_nl;
  wire[0:0] or_697_nl;
  wire[0:0] or_696_nl;
  wire[0:0] mux_1091_nl;
  wire[0:0] mux_1090_nl;
  wire[0:0] mux_1089_nl;
  wire[0:0] mux_1088_nl;
  wire[0:0] mux_1087_nl;
  wire[0:0] or_692_nl;
  wire[0:0] mux_1086_nl;
  wire[0:0] or_691_nl;
  wire[0:0] nand_15_nl;
  wire[0:0] mux_1084_nl;
  wire[0:0] mux_1083_nl;
  wire[0:0] nor_771_nl;
  wire[0:0] nor_772_nl;
  wire[0:0] mux_1082_nl;
  wire[0:0] nor_773_nl;
  wire[0:0] nor_774_nl;
  wire[0:0] mux_1081_nl;
  wire[0:0] mux_1080_nl;
  wire[0:0] mux_1079_nl;
  wire[0:0] or_680_nl;
  wire[0:0] mux_1078_nl;
  wire[0:0] or_678_nl;
  wire[0:0] or_676_nl;
  wire[0:0] or_675_nl;
  wire[0:0] mux_1077_nl;
  wire[0:0] or_674_nl;
  wire[0:0] or_673_nl;
  wire[0:0] or_672_nl;
  wire[0:0] mux_1076_nl;
  wire[0:0] mux_1075_nl;
  wire[0:0] or_671_nl;
  wire[0:0] or_670_nl;
  wire[0:0] or_668_nl;
  wire[0:0] mux_1142_nl;
  wire[0:0] mux_1141_nl;
  wire[0:0] mux_1140_nl;
  wire[0:0] mux_1139_nl;
  wire[0:0] or_775_nl;
  wire[0:0] mux_1138_nl;
  wire[0:0] or_773_nl;
  wire[0:0] mux_1137_nl;
  wire[0:0] or_772_nl;
  wire[0:0] or_771_nl;
  wire[0:0] mux_1136_nl;
  wire[0:0] mux_1135_nl;
  wire[0:0] mux_1134_nl;
  wire[0:0] or_770_nl;
  wire[0:0] or_768_nl;
  wire[0:0] or_766_nl;
  wire[0:0] or_764_nl;
  wire[0:0] mux_1133_nl;
  wire[0:0] mux_1132_nl;
  wire[0:0] mux_1131_nl;
  wire[0:0] mux_1130_nl;
  wire[0:0] or_763_nl;
  wire[0:0] or_762_nl;
  wire[0:0] or_761_nl;
  wire[0:0] or_760_nl;
  wire[0:0] mux_1129_nl;
  wire[0:0] mux_1128_nl;
  wire[0:0] or_758_nl;
  wire[0:0] mux_1127_nl;
  wire[0:0] or_757_nl;
  wire[0:0] or_756_nl;
  wire[0:0] or_755_nl;
  wire[0:0] mux_1126_nl;
  wire[0:0] mux_1125_nl;
  wire[0:0] mux_1124_nl;
  wire[0:0] mux_1123_nl;
  wire[0:0] mux_1122_nl;
  wire[0:0] or_754_nl;
  wire[0:0] or_752_nl;
  wire[0:0] or_750_nl;
  wire[0:0] nand_20_nl;
  wire[0:0] mux_1121_nl;
  wire[0:0] mux_1120_nl;
  wire[0:0] mux_1119_nl;
  wire[0:0] or_748_nl;
  wire[0:0] or_747_nl;
  wire[0:0] or_745_nl;
  wire[0:0] or_744_nl;
  wire[0:0] mux_1118_nl;
  wire[0:0] mux_1117_nl;
  wire[0:0] or_742_nl;
  wire[0:0] or_740_nl;
  wire[0:0] mux_1116_nl;
  wire[0:0] or_739_nl;
  wire[0:0] mux_1115_nl;
  wire[0:0] or_737_nl;
  wire[0:0] mux_1114_nl;
  wire[0:0] mux_1113_nl;
  wire[0:0] or_730_nl;
  wire[0:0] or_729_nl;
  wire[0:0] or_727_nl;
  wire[0:0] or_726_nl;
  wire[0:0] mux_1110_nl;
  wire[0:0] or_725_nl;
  wire[0:0] mux_1109_nl;
  wire[0:0] or_724_nl;
  wire[0:0] mux_1108_nl;
  wire[0:0] or_723_nl;
  wire[0:0] or_722_nl;
  wire[0:0] mux_1175_nl;
  wire[0:0] mux_1174_nl;
  wire[0:0] mux_1173_nl;
  wire[0:0] nand_24_nl;
  wire[0:0] mux_1172_nl;
  wire[0:0] mux_1171_nl;
  wire[0:0] nor_753_nl;
  wire[0:0] nor_754_nl;
  wire[0:0] mux_1170_nl;
  wire[0:0] nor_755_nl;
  wire[0:0] nor_756_nl;
  wire[0:0] mux_1169_nl;
  wire[0:0] nand_23_nl;
  wire[0:0] mux_1168_nl;
  wire[0:0] nor_757_nl;
  wire[0:0] nor_758_nl;
  wire[0:0] mux_1167_nl;
  wire[0:0] mux_1166_nl;
  wire[0:0] or_820_nl;
  wire[0:0] or_818_nl;
  wire[0:0] or_817_nl;
  wire[0:0] mux_1165_nl;
  wire[0:0] or_816_nl;
  wire[0:0] mux_1164_nl;
  wire[0:0] mux_1163_nl;
  wire[0:0] or_815_nl;
  wire[0:0] or_814_nl;
  wire[0:0] mux_1162_nl;
  wire[0:0] or_812_nl;
  wire[0:0] or_810_nl;
  wire[0:0] mux_1161_nl;
  wire[0:0] or_808_nl;
  wire[0:0] mux_1160_nl;
  wire[0:0] or_807_nl;
  wire[0:0] or_806_nl;
  wire[0:0] or_805_nl;
  wire[0:0] mux_1159_nl;
  wire[0:0] mux_1158_nl;
  wire[0:0] mux_1157_nl;
  wire[0:0] mux_1156_nl;
  wire[0:0] mux_1155_nl;
  wire[0:0] or_801_nl;
  wire[0:0] mux_1154_nl;
  wire[0:0] or_800_nl;
  wire[0:0] nand_21_nl;
  wire[0:0] mux_1152_nl;
  wire[0:0] mux_1151_nl;
  wire[0:0] nor_759_nl;
  wire[0:0] nor_760_nl;
  wire[0:0] mux_1150_nl;
  wire[0:0] nor_761_nl;
  wire[0:0] nor_762_nl;
  wire[0:0] mux_1149_nl;
  wire[0:0] mux_1148_nl;
  wire[0:0] mux_1147_nl;
  wire[0:0] or_789_nl;
  wire[0:0] mux_1146_nl;
  wire[0:0] or_787_nl;
  wire[0:0] or_785_nl;
  wire[0:0] or_784_nl;
  wire[0:0] mux_1145_nl;
  wire[0:0] or_783_nl;
  wire[0:0] or_782_nl;
  wire[0:0] or_781_nl;
  wire[0:0] mux_1144_nl;
  wire[0:0] mux_1143_nl;
  wire[0:0] or_780_nl;
  wire[0:0] or_779_nl;
  wire[0:0] or_777_nl;
  wire[0:0] mux_1210_nl;
  wire[0:0] mux_1209_nl;
  wire[0:0] mux_1208_nl;
  wire[0:0] mux_1207_nl;
  wire[0:0] or_881_nl;
  wire[0:0] mux_1206_nl;
  wire[0:0] or_879_nl;
  wire[0:0] mux_1205_nl;
  wire[0:0] or_878_nl;
  wire[0:0] or_877_nl;
  wire[0:0] mux_1204_nl;
  wire[0:0] mux_1203_nl;
  wire[0:0] mux_1202_nl;
  wire[0:0] or_876_nl;
  wire[0:0] or_874_nl;
  wire[0:0] or_872_nl;
  wire[0:0] or_870_nl;
  wire[0:0] mux_1201_nl;
  wire[0:0] mux_1200_nl;
  wire[0:0] mux_1199_nl;
  wire[0:0] mux_1198_nl;
  wire[0:0] or_869_nl;
  wire[0:0] or_868_nl;
  wire[0:0] or_867_nl;
  wire[0:0] or_866_nl;
  wire[0:0] mux_1197_nl;
  wire[0:0] mux_1196_nl;
  wire[0:0] or_864_nl;
  wire[0:0] mux_1195_nl;
  wire[0:0] or_863_nl;
  wire[0:0] or_862_nl;
  wire[0:0] or_861_nl;
  wire[0:0] mux_1194_nl;
  wire[0:0] mux_1193_nl;
  wire[0:0] mux_1192_nl;
  wire[0:0] mux_1191_nl;
  wire[0:0] mux_1190_nl;
  wire[0:0] or_860_nl;
  wire[0:0] or_858_nl;
  wire[0:0] or_856_nl;
  wire[0:0] nand_26_nl;
  wire[0:0] mux_1189_nl;
  wire[0:0] mux_1188_nl;
  wire[0:0] or_854_nl;
  wire[0:0] mux_1187_nl;
  wire[0:0] or_852_nl;
  wire[0:0] nor_277_nl;
  wire[0:0] or_851_nl;
  wire[0:0] mux_1186_nl;
  wire[0:0] mux_1185_nl;
  wire[0:0] or_849_nl;
  wire[0:0] or_847_nl;
  wire[0:0] mux_1184_nl;
  wire[0:0] or_846_nl;
  wire[0:0] mux_1183_nl;
  wire[0:0] or_844_nl;
  wire[0:0] mux_1182_nl;
  wire[0:0] or_842_nl;
  wire[0:0] mux_1181_nl;
  wire[0:0] nor_275_nl;
  wire[0:0] nor_274_nl;
  wire[0:0] or_835_nl;
  wire[0:0] mux_1178_nl;
  wire[0:0] or_834_nl;
  wire[0:0] mux_1177_nl;
  wire[0:0] or_833_nl;
  wire[0:0] mux_1176_nl;
  wire[0:0] or_832_nl;
  wire[0:0] or_831_nl;
  wire[0:0] mux_1243_nl;
  wire[0:0] mux_1242_nl;
  wire[0:0] mux_1241_nl;
  wire[0:0] nand_30_nl;
  wire[0:0] mux_1240_nl;
  wire[0:0] mux_1239_nl;
  wire[0:0] nor_741_nl;
  wire[0:0] nor_742_nl;
  wire[0:0] mux_1238_nl;
  wire[0:0] nor_743_nl;
  wire[0:0] nor_744_nl;
  wire[0:0] mux_1237_nl;
  wire[0:0] nand_29_nl;
  wire[0:0] mux_1236_nl;
  wire[0:0] nor_745_nl;
  wire[0:0] nor_746_nl;
  wire[0:0] mux_1235_nl;
  wire[0:0] mux_1234_nl;
  wire[0:0] or_926_nl;
  wire[0:0] or_924_nl;
  wire[0:0] or_923_nl;
  wire[0:0] mux_1233_nl;
  wire[0:0] or_922_nl;
  wire[0:0] mux_1232_nl;
  wire[0:0] mux_1231_nl;
  wire[0:0] or_921_nl;
  wire[0:0] or_920_nl;
  wire[0:0] mux_1230_nl;
  wire[0:0] or_918_nl;
  wire[0:0] or_916_nl;
  wire[0:0] mux_1229_nl;
  wire[0:0] or_914_nl;
  wire[0:0] mux_1228_nl;
  wire[0:0] or_913_nl;
  wire[0:0] or_912_nl;
  wire[0:0] or_911_nl;
  wire[0:0] mux_1227_nl;
  wire[0:0] mux_1226_nl;
  wire[0:0] mux_1225_nl;
  wire[0:0] mux_1224_nl;
  wire[0:0] mux_1223_nl;
  wire[0:0] or_907_nl;
  wire[0:0] mux_1222_nl;
  wire[0:0] or_906_nl;
  wire[0:0] nand_27_nl;
  wire[0:0] mux_1220_nl;
  wire[0:0] mux_1219_nl;
  wire[0:0] nor_747_nl;
  wire[0:0] nor_748_nl;
  wire[0:0] mux_1218_nl;
  wire[0:0] nor_749_nl;
  wire[0:0] nor_750_nl;
  wire[0:0] mux_1217_nl;
  wire[0:0] mux_1216_nl;
  wire[0:0] mux_1215_nl;
  wire[0:0] or_895_nl;
  wire[0:0] mux_1214_nl;
  wire[0:0] or_893_nl;
  wire[0:0] or_891_nl;
  wire[0:0] or_890_nl;
  wire[0:0] mux_1213_nl;
  wire[0:0] or_889_nl;
  wire[0:0] or_888_nl;
  wire[0:0] or_887_nl;
  wire[0:0] mux_1212_nl;
  wire[0:0] mux_1211_nl;
  wire[0:0] or_886_nl;
  wire[0:0] or_885_nl;
  wire[0:0] or_883_nl;
  wire[0:0] mux_1278_nl;
  wire[0:0] mux_1277_nl;
  wire[0:0] mux_1276_nl;
  wire[0:0] mux_1275_nl;
  wire[0:0] or_990_nl;
  wire[0:0] mux_1274_nl;
  wire[0:0] or_988_nl;
  wire[0:0] mux_1273_nl;
  wire[0:0] or_987_nl;
  wire[0:0] or_986_nl;
  wire[0:0] mux_1272_nl;
  wire[0:0] mux_1271_nl;
  wire[0:0] mux_1270_nl;
  wire[0:0] or_985_nl;
  wire[0:0] or_983_nl;
  wire[0:0] or_981_nl;
  wire[0:0] or_979_nl;
  wire[0:0] mux_1269_nl;
  wire[0:0] mux_1268_nl;
  wire[0:0] mux_1267_nl;
  wire[0:0] mux_1266_nl;
  wire[0:0] or_978_nl;
  wire[0:0] or_977_nl;
  wire[0:0] or_976_nl;
  wire[0:0] or_975_nl;
  wire[0:0] mux_1265_nl;
  wire[0:0] mux_1264_nl;
  wire[0:0] or_973_nl;
  wire[0:0] mux_1263_nl;
  wire[0:0] or_972_nl;
  wire[0:0] or_971_nl;
  wire[0:0] or_970_nl;
  wire[0:0] mux_1262_nl;
  wire[0:0] mux_1261_nl;
  wire[0:0] mux_1260_nl;
  wire[0:0] mux_1259_nl;
  wire[0:0] mux_1258_nl;
  wire[0:0] or_969_nl;
  wire[0:0] or_967_nl;
  wire[0:0] or_965_nl;
  wire[0:0] nand_32_nl;
  wire[0:0] mux_1257_nl;
  wire[0:0] mux_1256_nl;
  wire[0:0] mux_1255_nl;
  wire[0:0] or_963_nl;
  wire[0:0] or_962_nl;
  wire[0:0] or_960_nl;
  wire[0:0] or_959_nl;
  wire[0:0] mux_1254_nl;
  wire[0:0] mux_1253_nl;
  wire[0:0] or_957_nl;
  wire[0:0] or_955_nl;
  wire[0:0] mux_1252_nl;
  wire[0:0] or_954_nl;
  wire[0:0] mux_1251_nl;
  wire[0:0] or_952_nl;
  wire[0:0] mux_1250_nl;
  wire[0:0] mux_1249_nl;
  wire[0:0] or_945_nl;
  wire[0:0] or_944_nl;
  wire[0:0] or_942_nl;
  wire[0:0] or_941_nl;
  wire[0:0] mux_1246_nl;
  wire[0:0] or_940_nl;
  wire[0:0] mux_1245_nl;
  wire[0:0] or_939_nl;
  wire[0:0] mux_1244_nl;
  wire[0:0] or_938_nl;
  wire[0:0] or_937_nl;
  wire[0:0] mux_1311_nl;
  wire[0:0] mux_1310_nl;
  wire[0:0] mux_1309_nl;
  wire[0:0] nand_36_nl;
  wire[0:0] mux_1308_nl;
  wire[0:0] mux_1307_nl;
  wire[0:0] nor_729_nl;
  wire[0:0] nor_730_nl;
  wire[0:0] mux_1306_nl;
  wire[0:0] nor_731_nl;
  wire[0:0] nor_732_nl;
  wire[0:0] mux_1305_nl;
  wire[0:0] nand_35_nl;
  wire[0:0] mux_1304_nl;
  wire[0:0] nor_733_nl;
  wire[0:0] nor_734_nl;
  wire[0:0] mux_1303_nl;
  wire[0:0] mux_1302_nl;
  wire[0:0] or_1035_nl;
  wire[0:0] or_1033_nl;
  wire[0:0] or_1032_nl;
  wire[0:0] mux_1301_nl;
  wire[0:0] or_1031_nl;
  wire[0:0] mux_1300_nl;
  wire[0:0] mux_1299_nl;
  wire[0:0] or_1030_nl;
  wire[0:0] or_1029_nl;
  wire[0:0] mux_1298_nl;
  wire[0:0] or_1027_nl;
  wire[0:0] or_1025_nl;
  wire[0:0] mux_1297_nl;
  wire[0:0] or_1023_nl;
  wire[0:0] mux_1296_nl;
  wire[0:0] or_1022_nl;
  wire[0:0] or_1021_nl;
  wire[0:0] or_1020_nl;
  wire[0:0] mux_1295_nl;
  wire[0:0] mux_1294_nl;
  wire[0:0] mux_1293_nl;
  wire[0:0] mux_1292_nl;
  wire[0:0] mux_1291_nl;
  wire[0:0] or_1016_nl;
  wire[0:0] mux_1290_nl;
  wire[0:0] or_1015_nl;
  wire[0:0] nand_33_nl;
  wire[0:0] mux_1288_nl;
  wire[0:0] mux_1287_nl;
  wire[0:0] nor_735_nl;
  wire[0:0] nor_736_nl;
  wire[0:0] mux_1286_nl;
  wire[0:0] nor_737_nl;
  wire[0:0] nor_738_nl;
  wire[0:0] mux_1285_nl;
  wire[0:0] mux_1284_nl;
  wire[0:0] mux_1283_nl;
  wire[0:0] or_1004_nl;
  wire[0:0] mux_1282_nl;
  wire[0:0] or_1002_nl;
  wire[0:0] or_1000_nl;
  wire[0:0] or_999_nl;
  wire[0:0] mux_1281_nl;
  wire[0:0] or_998_nl;
  wire[0:0] or_997_nl;
  wire[0:0] or_996_nl;
  wire[0:0] mux_1280_nl;
  wire[0:0] mux_1279_nl;
  wire[0:0] or_995_nl;
  wire[0:0] or_994_nl;
  wire[0:0] or_992_nl;
  wire[0:0] mux_1346_nl;
  wire[0:0] mux_1345_nl;
  wire[0:0] mux_1344_nl;
  wire[0:0] mux_1343_nl;
  wire[0:0] or_1096_nl;
  wire[0:0] mux_1342_nl;
  wire[0:0] or_1094_nl;
  wire[0:0] mux_1341_nl;
  wire[0:0] or_1093_nl;
  wire[0:0] or_1092_nl;
  wire[0:0] mux_1340_nl;
  wire[0:0] mux_1339_nl;
  wire[0:0] mux_1338_nl;
  wire[0:0] or_1091_nl;
  wire[0:0] or_1089_nl;
  wire[0:0] or_1087_nl;
  wire[0:0] or_1085_nl;
  wire[0:0] mux_1337_nl;
  wire[0:0] mux_1336_nl;
  wire[0:0] mux_1335_nl;
  wire[0:0] mux_1334_nl;
  wire[0:0] or_1084_nl;
  wire[0:0] or_1083_nl;
  wire[0:0] or_1082_nl;
  wire[0:0] or_1081_nl;
  wire[0:0] mux_1333_nl;
  wire[0:0] mux_1332_nl;
  wire[0:0] nand_357_nl;
  wire[0:0] mux_1331_nl;
  wire[0:0] or_1078_nl;
  wire[0:0] or_1077_nl;
  wire[0:0] or_1076_nl;
  wire[0:0] mux_1330_nl;
  wire[0:0] mux_1329_nl;
  wire[0:0] mux_1328_nl;
  wire[0:0] mux_1327_nl;
  wire[0:0] mux_1326_nl;
  wire[0:0] or_1075_nl;
  wire[0:0] or_1073_nl;
  wire[0:0] or_1071_nl;
  wire[0:0] nand_38_nl;
  wire[0:0] mux_1325_nl;
  wire[0:0] mux_1324_nl;
  wire[0:0] or_1069_nl;
  wire[0:0] mux_1323_nl;
  wire[0:0] or_1067_nl;
  wire[0:0] nor_288_nl;
  wire[0:0] or_1066_nl;
  wire[0:0] mux_1322_nl;
  wire[0:0] mux_1321_nl;
  wire[0:0] or_1064_nl;
  wire[0:0] or_1062_nl;
  wire[0:0] mux_1320_nl;
  wire[0:0] or_1061_nl;
  wire[0:0] mux_1319_nl;
  wire[0:0] or_1059_nl;
  wire[0:0] mux_1318_nl;
  wire[0:0] or_1057_nl;
  wire[0:0] mux_1317_nl;
  wire[0:0] nor_286_nl;
  wire[0:0] nor_285_nl;
  wire[0:0] or_1050_nl;
  wire[0:0] mux_1314_nl;
  wire[0:0] or_1049_nl;
  wire[0:0] mux_1313_nl;
  wire[0:0] or_1048_nl;
  wire[0:0] mux_1312_nl;
  wire[0:0] or_1047_nl;
  wire[0:0] or_1046_nl;
  wire[0:0] mux_1379_nl;
  wire[0:0] mux_1378_nl;
  wire[0:0] mux_1377_nl;
  wire[0:0] nand_42_nl;
  wire[0:0] mux_1376_nl;
  wire[0:0] mux_1375_nl;
  wire[0:0] nor_717_nl;
  wire[0:0] nor_718_nl;
  wire[0:0] mux_1374_nl;
  wire[0:0] nor_719_nl;
  wire[0:0] nor_720_nl;
  wire[0:0] mux_1373_nl;
  wire[0:0] nand_41_nl;
  wire[0:0] mux_1372_nl;
  wire[0:0] nor_721_nl;
  wire[0:0] nor_722_nl;
  wire[0:0] mux_1371_nl;
  wire[0:0] mux_1370_nl;
  wire[0:0] or_1141_nl;
  wire[0:0] or_1139_nl;
  wire[0:0] or_1138_nl;
  wire[0:0] mux_1369_nl;
  wire[0:0] or_1137_nl;
  wire[0:0] mux_1368_nl;
  wire[0:0] mux_1367_nl;
  wire[0:0] or_1136_nl;
  wire[0:0] or_1135_nl;
  wire[0:0] mux_1366_nl;
  wire[0:0] or_1133_nl;
  wire[0:0] or_1131_nl;
  wire[0:0] mux_1365_nl;
  wire[0:0] or_1129_nl;
  wire[0:0] mux_1364_nl;
  wire[0:0] or_1128_nl;
  wire[0:0] or_1127_nl;
  wire[0:0] or_1126_nl;
  wire[0:0] mux_1363_nl;
  wire[0:0] mux_1362_nl;
  wire[0:0] mux_1361_nl;
  wire[0:0] mux_1360_nl;
  wire[0:0] mux_1359_nl;
  wire[0:0] or_1122_nl;
  wire[0:0] mux_1358_nl;
  wire[0:0] or_1121_nl;
  wire[0:0] nand_39_nl;
  wire[0:0] mux_1356_nl;
  wire[0:0] mux_1355_nl;
  wire[0:0] nor_723_nl;
  wire[0:0] nor_724_nl;
  wire[0:0] mux_1354_nl;
  wire[0:0] nor_725_nl;
  wire[0:0] nor_726_nl;
  wire[0:0] mux_1353_nl;
  wire[0:0] mux_1352_nl;
  wire[0:0] mux_1351_nl;
  wire[0:0] or_1110_nl;
  wire[0:0] mux_1350_nl;
  wire[0:0] or_1108_nl;
  wire[0:0] or_1106_nl;
  wire[0:0] or_1105_nl;
  wire[0:0] mux_1349_nl;
  wire[0:0] or_1104_nl;
  wire[0:0] or_1103_nl;
  wire[0:0] or_1102_nl;
  wire[0:0] mux_1348_nl;
  wire[0:0] mux_1347_nl;
  wire[0:0] or_1101_nl;
  wire[0:0] or_1100_nl;
  wire[0:0] or_1098_nl;
  wire[0:0] mux_1414_nl;
  wire[0:0] mux_1413_nl;
  wire[0:0] mux_1412_nl;
  wire[0:0] mux_1411_nl;
  wire[0:0] or_1205_nl;
  wire[0:0] mux_1410_nl;
  wire[0:0] or_1203_nl;
  wire[0:0] mux_1409_nl;
  wire[0:0] or_1202_nl;
  wire[0:0] or_1201_nl;
  wire[0:0] mux_1408_nl;
  wire[0:0] mux_1407_nl;
  wire[0:0] mux_1406_nl;
  wire[0:0] or_1200_nl;
  wire[0:0] or_1198_nl;
  wire[0:0] or_1196_nl;
  wire[0:0] or_1194_nl;
  wire[0:0] mux_1405_nl;
  wire[0:0] mux_1404_nl;
  wire[0:0] mux_1403_nl;
  wire[0:0] mux_1402_nl;
  wire[0:0] or_1193_nl;
  wire[0:0] or_1192_nl;
  wire[0:0] or_1191_nl;
  wire[0:0] or_1190_nl;
  wire[0:0] mux_1401_nl;
  wire[0:0] mux_1400_nl;
  wire[0:0] or_1188_nl;
  wire[0:0] mux_1399_nl;
  wire[0:0] or_1187_nl;
  wire[0:0] or_1186_nl;
  wire[0:0] or_1185_nl;
  wire[0:0] mux_1398_nl;
  wire[0:0] mux_1397_nl;
  wire[0:0] mux_1396_nl;
  wire[0:0] mux_1395_nl;
  wire[0:0] mux_1394_nl;
  wire[0:0] or_1184_nl;
  wire[0:0] or_1182_nl;
  wire[0:0] or_1180_nl;
  wire[0:0] nand_44_nl;
  wire[0:0] mux_1393_nl;
  wire[0:0] mux_1392_nl;
  wire[0:0] mux_1391_nl;
  wire[0:0] or_1178_nl;
  wire[0:0] or_1177_nl;
  wire[0:0] or_1175_nl;
  wire[0:0] or_1174_nl;
  wire[0:0] mux_1390_nl;
  wire[0:0] mux_1389_nl;
  wire[0:0] or_1172_nl;
  wire[0:0] or_1170_nl;
  wire[0:0] mux_1388_nl;
  wire[0:0] or_1169_nl;
  wire[0:0] mux_1387_nl;
  wire[0:0] or_1167_nl;
  wire[0:0] mux_1386_nl;
  wire[0:0] mux_1385_nl;
  wire[0:0] or_1160_nl;
  wire[0:0] or_1159_nl;
  wire[0:0] or_1157_nl;
  wire[0:0] or_1156_nl;
  wire[0:0] mux_1382_nl;
  wire[0:0] or_1155_nl;
  wire[0:0] mux_1381_nl;
  wire[0:0] or_1154_nl;
  wire[0:0] mux_1380_nl;
  wire[0:0] or_1153_nl;
  wire[0:0] or_1152_nl;
  wire[0:0] mux_1447_nl;
  wire[0:0] mux_1446_nl;
  wire[0:0] mux_1445_nl;
  wire[0:0] nand_48_nl;
  wire[0:0] mux_1444_nl;
  wire[0:0] mux_1443_nl;
  wire[0:0] nor_705_nl;
  wire[0:0] nor_706_nl;
  wire[0:0] mux_1442_nl;
  wire[0:0] nor_707_nl;
  wire[0:0] nor_708_nl;
  wire[0:0] mux_1441_nl;
  wire[0:0] nand_47_nl;
  wire[0:0] mux_1440_nl;
  wire[0:0] nor_709_nl;
  wire[0:0] nor_710_nl;
  wire[0:0] mux_1439_nl;
  wire[0:0] mux_1438_nl;
  wire[0:0] or_1250_nl;
  wire[0:0] or_1248_nl;
  wire[0:0] or_1247_nl;
  wire[0:0] mux_1437_nl;
  wire[0:0] or_1246_nl;
  wire[0:0] mux_1436_nl;
  wire[0:0] mux_1435_nl;
  wire[0:0] or_1245_nl;
  wire[0:0] or_1244_nl;
  wire[0:0] mux_1434_nl;
  wire[0:0] or_1242_nl;
  wire[0:0] or_1240_nl;
  wire[0:0] mux_1433_nl;
  wire[0:0] or_1238_nl;
  wire[0:0] mux_1432_nl;
  wire[0:0] or_1237_nl;
  wire[0:0] or_1236_nl;
  wire[0:0] or_1235_nl;
  wire[0:0] mux_1431_nl;
  wire[0:0] mux_1430_nl;
  wire[0:0] mux_1429_nl;
  wire[0:0] mux_1428_nl;
  wire[0:0] mux_1427_nl;
  wire[0:0] or_1231_nl;
  wire[0:0] mux_1426_nl;
  wire[0:0] or_1230_nl;
  wire[0:0] nand_45_nl;
  wire[0:0] mux_1424_nl;
  wire[0:0] mux_1423_nl;
  wire[0:0] nor_711_nl;
  wire[0:0] nor_712_nl;
  wire[0:0] mux_1422_nl;
  wire[0:0] nor_713_nl;
  wire[0:0] nor_714_nl;
  wire[0:0] mux_1421_nl;
  wire[0:0] mux_1420_nl;
  wire[0:0] mux_1419_nl;
  wire[0:0] or_1219_nl;
  wire[0:0] mux_1418_nl;
  wire[0:0] or_1217_nl;
  wire[0:0] or_1215_nl;
  wire[0:0] or_1214_nl;
  wire[0:0] mux_1417_nl;
  wire[0:0] or_1213_nl;
  wire[0:0] or_1212_nl;
  wire[0:0] or_1211_nl;
  wire[0:0] mux_1416_nl;
  wire[0:0] mux_1415_nl;
  wire[0:0] or_1210_nl;
  wire[0:0] or_1209_nl;
  wire[0:0] or_1207_nl;
  wire[0:0] mux_1482_nl;
  wire[0:0] mux_1481_nl;
  wire[0:0] mux_1480_nl;
  wire[0:0] mux_1479_nl;
  wire[0:0] or_1311_nl;
  wire[0:0] mux_1478_nl;
  wire[0:0] or_1309_nl;
  wire[0:0] mux_1477_nl;
  wire[0:0] or_1308_nl;
  wire[0:0] or_1307_nl;
  wire[0:0] mux_1476_nl;
  wire[0:0] mux_1475_nl;
  wire[0:0] mux_1474_nl;
  wire[0:0] or_1306_nl;
  wire[0:0] or_1304_nl;
  wire[0:0] or_1302_nl;
  wire[0:0] or_1300_nl;
  wire[0:0] mux_1473_nl;
  wire[0:0] mux_1472_nl;
  wire[0:0] mux_1471_nl;
  wire[0:0] mux_1470_nl;
  wire[0:0] or_1299_nl;
  wire[0:0] or_1298_nl;
  wire[0:0] or_1297_nl;
  wire[0:0] or_1296_nl;
  wire[0:0] mux_1469_nl;
  wire[0:0] mux_1468_nl;
  wire[0:0] nand_346_nl;
  wire[0:0] mux_1467_nl;
  wire[0:0] or_1293_nl;
  wire[0:0] or_1292_nl;
  wire[0:0] or_1291_nl;
  wire[0:0] mux_1466_nl;
  wire[0:0] mux_1465_nl;
  wire[0:0] mux_1464_nl;
  wire[0:0] mux_1463_nl;
  wire[0:0] mux_1462_nl;
  wire[0:0] or_1290_nl;
  wire[0:0] or_1288_nl;
  wire[0:0] or_1286_nl;
  wire[0:0] nand_50_nl;
  wire[0:0] mux_1461_nl;
  wire[0:0] mux_1460_nl;
  wire[0:0] or_1284_nl;
  wire[0:0] mux_1459_nl;
  wire[0:0] or_1282_nl;
  wire[0:0] nor_299_nl;
  wire[0:0] or_1281_nl;
  wire[0:0] mux_1458_nl;
  wire[0:0] mux_1457_nl;
  wire[0:0] or_1279_nl;
  wire[0:0] or_1277_nl;
  wire[0:0] mux_1456_nl;
  wire[0:0] or_1276_nl;
  wire[0:0] mux_1455_nl;
  wire[0:0] or_1274_nl;
  wire[0:0] mux_1454_nl;
  wire[0:0] or_1272_nl;
  wire[0:0] mux_1453_nl;
  wire[0:0] nor_297_nl;
  wire[0:0] nor_296_nl;
  wire[0:0] or_1265_nl;
  wire[0:0] mux_1450_nl;
  wire[0:0] or_1264_nl;
  wire[0:0] mux_1449_nl;
  wire[0:0] or_1263_nl;
  wire[0:0] mux_1448_nl;
  wire[0:0] or_1262_nl;
  wire[0:0] or_1261_nl;
  wire[0:0] mux_1515_nl;
  wire[0:0] mux_1514_nl;
  wire[0:0] mux_1513_nl;
  wire[0:0] nand_54_nl;
  wire[0:0] mux_1512_nl;
  wire[0:0] mux_1511_nl;
  wire[0:0] nor_693_nl;
  wire[0:0] nor_694_nl;
  wire[0:0] mux_1510_nl;
  wire[0:0] nor_695_nl;
  wire[0:0] nor_696_nl;
  wire[0:0] mux_1509_nl;
  wire[0:0] nand_53_nl;
  wire[0:0] mux_1508_nl;
  wire[0:0] nor_697_nl;
  wire[0:0] nor_698_nl;
  wire[0:0] mux_1507_nl;
  wire[0:0] mux_1506_nl;
  wire[0:0] or_1356_nl;
  wire[0:0] or_1354_nl;
  wire[0:0] or_1353_nl;
  wire[0:0] mux_1505_nl;
  wire[0:0] or_1352_nl;
  wire[0:0] mux_1504_nl;
  wire[0:0] mux_1503_nl;
  wire[0:0] or_1351_nl;
  wire[0:0] or_1350_nl;
  wire[0:0] mux_1502_nl;
  wire[0:0] or_1348_nl;
  wire[0:0] or_1346_nl;
  wire[0:0] mux_1501_nl;
  wire[0:0] or_1344_nl;
  wire[0:0] mux_1500_nl;
  wire[0:0] or_1343_nl;
  wire[0:0] or_1342_nl;
  wire[0:0] or_1341_nl;
  wire[0:0] mux_1499_nl;
  wire[0:0] mux_1498_nl;
  wire[0:0] mux_1497_nl;
  wire[0:0] mux_1496_nl;
  wire[0:0] mux_1495_nl;
  wire[0:0] or_1337_nl;
  wire[0:0] mux_1494_nl;
  wire[0:0] or_1336_nl;
  wire[0:0] nand_51_nl;
  wire[0:0] mux_1492_nl;
  wire[0:0] mux_1491_nl;
  wire[0:0] nor_699_nl;
  wire[0:0] nor_700_nl;
  wire[0:0] mux_1490_nl;
  wire[0:0] nor_701_nl;
  wire[0:0] nor_702_nl;
  wire[0:0] mux_1489_nl;
  wire[0:0] mux_1488_nl;
  wire[0:0] mux_1487_nl;
  wire[0:0] or_1325_nl;
  wire[0:0] mux_1486_nl;
  wire[0:0] or_1323_nl;
  wire[0:0] or_1321_nl;
  wire[0:0] or_1320_nl;
  wire[0:0] mux_1485_nl;
  wire[0:0] or_1319_nl;
  wire[0:0] or_1318_nl;
  wire[0:0] or_1317_nl;
  wire[0:0] mux_1484_nl;
  wire[0:0] mux_1483_nl;
  wire[0:0] or_1316_nl;
  wire[0:0] or_1315_nl;
  wire[0:0] or_1313_nl;
  wire[0:0] mux_1550_nl;
  wire[0:0] mux_1549_nl;
  wire[0:0] mux_1548_nl;
  wire[0:0] mux_1547_nl;
  wire[0:0] or_1420_nl;
  wire[0:0] mux_1546_nl;
  wire[0:0] or_1418_nl;
  wire[0:0] mux_1545_nl;
  wire[0:0] or_1417_nl;
  wire[0:0] or_1416_nl;
  wire[0:0] mux_1544_nl;
  wire[0:0] mux_1543_nl;
  wire[0:0] mux_1542_nl;
  wire[0:0] or_1415_nl;
  wire[0:0] or_1413_nl;
  wire[0:0] or_1411_nl;
  wire[0:0] or_1409_nl;
  wire[0:0] mux_1541_nl;
  wire[0:0] mux_1540_nl;
  wire[0:0] mux_1539_nl;
  wire[0:0] mux_1538_nl;
  wire[0:0] or_1408_nl;
  wire[0:0] or_1407_nl;
  wire[0:0] or_1406_nl;
  wire[0:0] or_1405_nl;
  wire[0:0] mux_1537_nl;
  wire[0:0] mux_1536_nl;
  wire[0:0] nand_340_nl;
  wire[0:0] mux_1535_nl;
  wire[0:0] or_1402_nl;
  wire[0:0] or_1401_nl;
  wire[0:0] or_1400_nl;
  wire[0:0] mux_1534_nl;
  wire[0:0] mux_1533_nl;
  wire[0:0] mux_1532_nl;
  wire[0:0] mux_1531_nl;
  wire[0:0] mux_1530_nl;
  wire[0:0] or_1399_nl;
  wire[0:0] or_1397_nl;
  wire[0:0] or_1395_nl;
  wire[0:0] nand_56_nl;
  wire[0:0] mux_1529_nl;
  wire[0:0] mux_1528_nl;
  wire[0:0] mux_1527_nl;
  wire[0:0] or_1393_nl;
  wire[0:0] or_1392_nl;
  wire[0:0] or_1390_nl;
  wire[0:0] or_1389_nl;
  wire[0:0] mux_1526_nl;
  wire[0:0] mux_1525_nl;
  wire[0:0] or_1387_nl;
  wire[0:0] or_1385_nl;
  wire[0:0] mux_1524_nl;
  wire[0:0] or_1384_nl;
  wire[0:0] mux_1523_nl;
  wire[0:0] or_1382_nl;
  wire[0:0] mux_1522_nl;
  wire[0:0] mux_1521_nl;
  wire[0:0] or_1375_nl;
  wire[0:0] or_1374_nl;
  wire[0:0] or_1372_nl;
  wire[0:0] or_1371_nl;
  wire[0:0] mux_1518_nl;
  wire[0:0] or_1370_nl;
  wire[0:0] mux_1517_nl;
  wire[0:0] or_1369_nl;
  wire[0:0] mux_1516_nl;
  wire[0:0] or_1368_nl;
  wire[0:0] or_1367_nl;
  wire[0:0] mux_1583_nl;
  wire[0:0] mux_1582_nl;
  wire[0:0] mux_1581_nl;
  wire[0:0] nand_60_nl;
  wire[0:0] mux_1580_nl;
  wire[0:0] mux_1579_nl;
  wire[0:0] nor_681_nl;
  wire[0:0] nor_682_nl;
  wire[0:0] mux_1578_nl;
  wire[0:0] and_773_nl;
  wire[0:0] and_779_nl;
  wire[0:0] mux_1577_nl;
  wire[0:0] nand_59_nl;
  wire[0:0] mux_1576_nl;
  wire[0:0] nor_685_nl;
  wire[0:0] nor_686_nl;
  wire[0:0] mux_1575_nl;
  wire[0:0] mux_1574_nl;
  wire[0:0] or_1465_nl;
  wire[0:0] or_1463_nl;
  wire[0:0] or_1462_nl;
  wire[0:0] mux_1573_nl;
  wire[0:0] or_1461_nl;
  wire[0:0] mux_1572_nl;
  wire[0:0] mux_1571_nl;
  wire[0:0] nand_331_nl;
  wire[0:0] nand_472_nl;
  wire[0:0] mux_1570_nl;
  wire[0:0] or_1457_nl;
  wire[0:0] or_1455_nl;
  wire[0:0] mux_1569_nl;
  wire[0:0] or_1453_nl;
  wire[0:0] mux_1568_nl;
  wire[0:0] or_1452_nl;
  wire[0:0] or_1451_nl;
  wire[0:0] or_1450_nl;
  wire[0:0] mux_1567_nl;
  wire[0:0] mux_1566_nl;
  wire[0:0] mux_1565_nl;
  wire[0:0] mux_1564_nl;
  wire[0:0] mux_1563_nl;
  wire[0:0] or_1446_nl;
  wire[0:0] mux_1562_nl;
  wire[0:0] or_1445_nl;
  wire[0:0] nand_57_nl;
  wire[0:0] mux_1560_nl;
  wire[0:0] mux_1559_nl;
  wire[0:0] nor_687_nl;
  wire[0:0] nor_688_nl;
  wire[0:0] mux_1558_nl;
  wire[0:0] and_789_nl;
  wire[0:0] and_790_nl;
  wire[0:0] mux_1557_nl;
  wire[0:0] mux_1556_nl;
  wire[0:0] mux_1555_nl;
  wire[0:0] or_1434_nl;
  wire[0:0] mux_1554_nl;
  wire[0:0] or_1432_nl;
  wire[0:0] or_1430_nl;
  wire[0:0] or_1429_nl;
  wire[0:0] mux_1553_nl;
  wire[0:0] or_1428_nl;
  wire[0:0] or_1427_nl;
  wire[0:0] or_1426_nl;
  wire[0:0] mux_1552_nl;
  wire[0:0] mux_1551_nl;
  wire[0:0] nand_336_nl;
  wire[0:0] nand_453_nl;
  wire[0:0] or_1422_nl;
  wire[0:0] mux_1618_nl;
  wire[0:0] mux_1617_nl;
  wire[0:0] mux_1616_nl;
  wire[0:0] mux_1615_nl;
  wire[0:0] or_1526_nl;
  wire[0:0] mux_1614_nl;
  wire[0:0] nand_317_nl;
  wire[0:0] mux_1613_nl;
  wire[0:0] or_1523_nl;
  wire[0:0] or_1522_nl;
  wire[0:0] mux_1612_nl;
  wire[0:0] mux_1611_nl;
  wire[0:0] mux_1610_nl;
  wire[0:0] or_1521_nl;
  wire[0:0] or_1519_nl;
  wire[0:0] or_1517_nl;
  wire[0:0] or_1515_nl;
  wire[0:0] mux_1609_nl;
  wire[0:0] mux_1608_nl;
  wire[0:0] mux_1607_nl;
  wire[0:0] mux_1606_nl;
  wire[0:0] nand_318_nl;
  wire[0:0] nand_319_nl;
  wire[0:0] or_1512_nl;
  wire[0:0] or_1511_nl;
  wire[0:0] mux_1605_nl;
  wire[0:0] mux_1604_nl;
  wire[0:0] nand_320_nl;
  wire[0:0] mux_1603_nl;
  wire[0:0] or_1508_nl;
  wire[0:0] or_1507_nl;
  wire[0:0] or_1506_nl;
  wire[0:0] mux_1602_nl;
  wire[0:0] mux_1601_nl;
  wire[0:0] mux_1600_nl;
  wire[0:0] mux_1599_nl;
  wire[0:0] mux_1598_nl;
  wire[0:0] or_1505_nl;
  wire[0:0] or_1503_nl;
  wire[0:0] or_1501_nl;
  wire[0:0] nand_62_nl;
  wire[0:0] mux_1597_nl;
  wire[0:0] mux_1596_nl;
  wire[0:0] nand_467_nl;
  wire[0:0] mux_1595_nl;
  wire[0:0] nand_323_nl;
  wire[0:0] and_546_nl;
  wire[0:0] nand_463_nl;
  wire[0:0] mux_1594_nl;
  wire[0:0] mux_1593_nl;
  wire[0:0] or_1494_nl;
  wire[0:0] or_1492_nl;
  wire[0:0] mux_1592_nl;
  wire[0:0] or_1491_nl;
  wire[0:0] mux_1591_nl;
  wire[0:0] or_1489_nl;
  wire[0:0] mux_1590_nl;
  wire[0:0] or_1487_nl;
  wire[0:0] mux_1589_nl;
  wire[0:0] and_547_nl;
  wire[0:0] and_548_nl;
  wire[0:0] or_1480_nl;
  wire[0:0] mux_1586_nl;
  wire[0:0] or_1479_nl;
  wire[0:0] mux_1585_nl;
  wire[0:0] or_1478_nl;
  wire[0:0] mux_1584_nl;
  wire[0:0] or_1477_nl;
  wire[0:0] or_1476_nl;
  wire[0:0] mux_1651_nl;
  wire[0:0] mux_1650_nl;
  wire[0:0] mux_1649_nl;
  wire[0:0] nand_66_nl;
  wire[0:0] mux_1648_nl;
  wire[0:0] mux_1647_nl;
  wire[0:0] nor_669_nl;
  wire[0:0] nor_670_nl;
  wire[0:0] mux_1646_nl;
  wire[0:0] nor_671_nl;
  wire[0:0] nor_672_nl;
  wire[0:0] mux_1645_nl;
  wire[0:0] nand_65_nl;
  wire[0:0] mux_1644_nl;
  wire[0:0] nor_673_nl;
  wire[0:0] nor_674_nl;
  wire[0:0] mux_1643_nl;
  wire[0:0] mux_1642_nl;
  wire[0:0] or_1571_nl;
  wire[0:0] or_1569_nl;
  wire[0:0] or_1568_nl;
  wire[0:0] mux_1641_nl;
  wire[0:0] or_1567_nl;
  wire[0:0] mux_1640_nl;
  wire[0:0] mux_1639_nl;
  wire[0:0] or_1566_nl;
  wire[0:0] or_1565_nl;
  wire[0:0] mux_1638_nl;
  wire[0:0] or_1563_nl;
  wire[0:0] or_1561_nl;
  wire[0:0] mux_1637_nl;
  wire[0:0] or_1559_nl;
  wire[0:0] mux_1636_nl;
  wire[0:0] or_1558_nl;
  wire[0:0] or_1557_nl;
  wire[0:0] or_1556_nl;
  wire[0:0] mux_1635_nl;
  wire[0:0] mux_1634_nl;
  wire[0:0] mux_1633_nl;
  wire[0:0] mux_1632_nl;
  wire[0:0] or_1554_nl;
  wire[0:0] mux_1631_nl;
  wire[0:0] mux_1630_nl;
  wire[0:0] or_1551_nl;
  wire[0:0] nand_63_nl;
  wire[0:0] mux_1628_nl;
  wire[0:0] mux_1627_nl;
  wire[0:0] nor_675_nl;
  wire[0:0] nor_676_nl;
  wire[0:0] mux_1626_nl;
  wire[0:0] nor_677_nl;
  wire[0:0] nor_678_nl;
  wire[0:0] mux_1625_nl;
  wire[0:0] mux_1624_nl;
  wire[0:0] mux_1623_nl;
  wire[0:0] or_1540_nl;
  wire[0:0] mux_1622_nl;
  wire[0:0] or_1538_nl;
  wire[0:0] or_1536_nl;
  wire[0:0] or_1535_nl;
  wire[0:0] mux_1621_nl;
  wire[0:0] or_1534_nl;
  wire[0:0] or_1533_nl;
  wire[0:0] or_1532_nl;
  wire[0:0] mux_1620_nl;
  wire[0:0] mux_1619_nl;
  wire[0:0] or_1531_nl;
  wire[0:0] or_1530_nl;
  wire[0:0] or_1528_nl;
  wire[0:0] mux_1686_nl;
  wire[0:0] mux_1685_nl;
  wire[0:0] mux_1684_nl;
  wire[0:0] mux_1683_nl;
  wire[0:0] or_1635_nl;
  wire[0:0] mux_1682_nl;
  wire[0:0] or_1633_nl;
  wire[0:0] mux_1681_nl;
  wire[0:0] or_1632_nl;
  wire[0:0] or_1631_nl;
  wire[0:0] mux_1680_nl;
  wire[0:0] mux_1679_nl;
  wire[0:0] mux_1678_nl;
  wire[0:0] or_1630_nl;
  wire[0:0] or_1628_nl;
  wire[0:0] or_1626_nl;
  wire[0:0] or_1624_nl;
  wire[0:0] mux_1677_nl;
  wire[0:0] mux_1676_nl;
  wire[0:0] mux_1675_nl;
  wire[0:0] mux_1674_nl;
  wire[0:0] or_1623_nl;
  wire[0:0] or_1622_nl;
  wire[0:0] or_1621_nl;
  wire[0:0] or_1620_nl;
  wire[0:0] mux_1673_nl;
  wire[0:0] mux_1672_nl;
  wire[0:0] or_1618_nl;
  wire[0:0] mux_1671_nl;
  wire[0:0] or_1617_nl;
  wire[0:0] or_1616_nl;
  wire[0:0] or_1615_nl;
  wire[0:0] mux_1670_nl;
  wire[0:0] mux_1669_nl;
  wire[0:0] mux_1668_nl;
  wire[0:0] mux_1667_nl;
  wire[0:0] mux_1666_nl;
  wire[0:0] or_1614_nl;
  wire[0:0] or_1612_nl;
  wire[0:0] or_1610_nl;
  wire[0:0] nand_68_nl;
  wire[0:0] mux_1665_nl;
  wire[0:0] mux_1664_nl;
  wire[0:0] mux_1663_nl;
  wire[0:0] or_1608_nl;
  wire[0:0] or_1607_nl;
  wire[0:0] or_1605_nl;
  wire[0:0] or_1604_nl;
  wire[0:0] mux_1662_nl;
  wire[0:0] mux_1661_nl;
  wire[0:0] or_1602_nl;
  wire[0:0] or_1600_nl;
  wire[0:0] mux_1660_nl;
  wire[0:0] or_1599_nl;
  wire[0:0] mux_1659_nl;
  wire[0:0] or_1597_nl;
  wire[0:0] mux_1658_nl;
  wire[0:0] mux_1657_nl;
  wire[0:0] or_1590_nl;
  wire[0:0] or_1589_nl;
  wire[0:0] or_1587_nl;
  wire[0:0] or_1586_nl;
  wire[0:0] mux_1654_nl;
  wire[0:0] or_1585_nl;
  wire[0:0] mux_1653_nl;
  wire[0:0] or_1584_nl;
  wire[0:0] mux_1652_nl;
  wire[0:0] or_1583_nl;
  wire[0:0] or_1582_nl;
  wire[0:0] mux_1719_nl;
  wire[0:0] mux_1718_nl;
  wire[0:0] mux_1717_nl;
  wire[0:0] nand_72_nl;
  wire[0:0] mux_1716_nl;
  wire[0:0] mux_1715_nl;
  wire[0:0] nor_657_nl;
  wire[0:0] nor_658_nl;
  wire[0:0] mux_1714_nl;
  wire[0:0] nor_659_nl;
  wire[0:0] nor_660_nl;
  wire[0:0] mux_1713_nl;
  wire[0:0] nand_71_nl;
  wire[0:0] mux_1712_nl;
  wire[0:0] nor_661_nl;
  wire[0:0] nor_662_nl;
  wire[0:0] mux_1711_nl;
  wire[0:0] mux_1710_nl;
  wire[0:0] or_1680_nl;
  wire[0:0] or_1678_nl;
  wire[0:0] or_1677_nl;
  wire[0:0] mux_1709_nl;
  wire[0:0] or_1676_nl;
  wire[0:0] mux_1708_nl;
  wire[0:0] mux_1707_nl;
  wire[0:0] or_1675_nl;
  wire[0:0] or_1674_nl;
  wire[0:0] mux_1706_nl;
  wire[0:0] or_1672_nl;
  wire[0:0] or_1670_nl;
  wire[0:0] mux_1705_nl;
  wire[0:0] or_1668_nl;
  wire[0:0] mux_1704_nl;
  wire[0:0] or_1667_nl;
  wire[0:0] or_1666_nl;
  wire[0:0] or_1665_nl;
  wire[0:0] mux_1703_nl;
  wire[0:0] mux_1702_nl;
  wire[0:0] mux_1701_nl;
  wire[0:0] mux_1700_nl;
  wire[0:0] or_1663_nl;
  wire[0:0] mux_1699_nl;
  wire[0:0] mux_1698_nl;
  wire[0:0] or_1660_nl;
  wire[0:0] nand_69_nl;
  wire[0:0] mux_1696_nl;
  wire[0:0] mux_1695_nl;
  wire[0:0] nor_663_nl;
  wire[0:0] nor_664_nl;
  wire[0:0] mux_1694_nl;
  wire[0:0] nor_665_nl;
  wire[0:0] nor_666_nl;
  wire[0:0] mux_1693_nl;
  wire[0:0] mux_1692_nl;
  wire[0:0] mux_1691_nl;
  wire[0:0] or_1649_nl;
  wire[0:0] mux_1690_nl;
  wire[0:0] or_1647_nl;
  wire[0:0] or_1645_nl;
  wire[0:0] or_1644_nl;
  wire[0:0] mux_1689_nl;
  wire[0:0] or_1643_nl;
  wire[0:0] or_1642_nl;
  wire[0:0] or_1641_nl;
  wire[0:0] mux_1688_nl;
  wire[0:0] mux_1687_nl;
  wire[0:0] or_1640_nl;
  wire[0:0] or_1639_nl;
  wire[0:0] or_1637_nl;
  wire[0:0] mux_1754_nl;
  wire[0:0] mux_1753_nl;
  wire[0:0] mux_1752_nl;
  wire[0:0] mux_1751_nl;
  wire[0:0] or_1741_nl;
  wire[0:0] mux_1750_nl;
  wire[0:0] or_1739_nl;
  wire[0:0] mux_1749_nl;
  wire[0:0] or_1738_nl;
  wire[0:0] or_1737_nl;
  wire[0:0] mux_1748_nl;
  wire[0:0] mux_1747_nl;
  wire[0:0] mux_1746_nl;
  wire[0:0] or_1736_nl;
  wire[0:0] or_1734_nl;
  wire[0:0] or_1732_nl;
  wire[0:0] or_1730_nl;
  wire[0:0] mux_1745_nl;
  wire[0:0] mux_1744_nl;
  wire[0:0] mux_1743_nl;
  wire[0:0] mux_1742_nl;
  wire[0:0] or_1729_nl;
  wire[0:0] or_1728_nl;
  wire[0:0] or_1727_nl;
  wire[0:0] or_1726_nl;
  wire[0:0] mux_1741_nl;
  wire[0:0] mux_1740_nl;
  wire[0:0] nand_306_nl;
  wire[0:0] mux_1739_nl;
  wire[0:0] or_1723_nl;
  wire[0:0] or_1722_nl;
  wire[0:0] or_1721_nl;
  wire[0:0] mux_1738_nl;
  wire[0:0] mux_1737_nl;
  wire[0:0] mux_1736_nl;
  wire[0:0] mux_1735_nl;
  wire[0:0] mux_1734_nl;
  wire[0:0] or_1720_nl;
  wire[0:0] or_1718_nl;
  wire[0:0] or_1716_nl;
  wire[0:0] nand_74_nl;
  wire[0:0] mux_1733_nl;
  wire[0:0] mux_1732_nl;
  wire[0:0] or_1714_nl;
  wire[0:0] mux_1731_nl;
  wire[0:0] or_1712_nl;
  wire[0:0] nor_321_nl;
  wire[0:0] or_1711_nl;
  wire[0:0] mux_1730_nl;
  wire[0:0] mux_1729_nl;
  wire[0:0] or_1709_nl;
  wire[0:0] or_1707_nl;
  wire[0:0] mux_1728_nl;
  wire[0:0] or_1706_nl;
  wire[0:0] mux_1727_nl;
  wire[0:0] or_1704_nl;
  wire[0:0] mux_1726_nl;
  wire[0:0] or_1702_nl;
  wire[0:0] mux_1725_nl;
  wire[0:0] nor_319_nl;
  wire[0:0] nor_318_nl;
  wire[0:0] or_1695_nl;
  wire[0:0] mux_1722_nl;
  wire[0:0] or_1694_nl;
  wire[0:0] mux_1721_nl;
  wire[0:0] or_1693_nl;
  wire[0:0] mux_1720_nl;
  wire[0:0] or_1692_nl;
  wire[0:0] or_1691_nl;
  wire[0:0] mux_1787_nl;
  wire[0:0] mux_1786_nl;
  wire[0:0] mux_1785_nl;
  wire[0:0] nand_78_nl;
  wire[0:0] mux_1784_nl;
  wire[0:0] mux_1783_nl;
  wire[0:0] nor_645_nl;
  wire[0:0] nor_646_nl;
  wire[0:0] mux_1782_nl;
  wire[0:0] nor_647_nl;
  wire[0:0] nor_648_nl;
  wire[0:0] mux_1781_nl;
  wire[0:0] nand_77_nl;
  wire[0:0] mux_1780_nl;
  wire[0:0] nor_649_nl;
  wire[0:0] nor_650_nl;
  wire[0:0] mux_1779_nl;
  wire[0:0] mux_1778_nl;
  wire[0:0] or_1786_nl;
  wire[0:0] or_1784_nl;
  wire[0:0] or_1783_nl;
  wire[0:0] mux_1777_nl;
  wire[0:0] or_1782_nl;
  wire[0:0] mux_1776_nl;
  wire[0:0] mux_1775_nl;
  wire[0:0] or_1781_nl;
  wire[0:0] or_1780_nl;
  wire[0:0] mux_1774_nl;
  wire[0:0] or_1778_nl;
  wire[0:0] or_1776_nl;
  wire[0:0] mux_1773_nl;
  wire[0:0] or_1774_nl;
  wire[0:0] mux_1772_nl;
  wire[0:0] or_1773_nl;
  wire[0:0] or_1772_nl;
  wire[0:0] or_1771_nl;
  wire[0:0] mux_1771_nl;
  wire[0:0] mux_1770_nl;
  wire[0:0] mux_1769_nl;
  wire[0:0] mux_1768_nl;
  wire[0:0] or_1769_nl;
  wire[0:0] mux_1767_nl;
  wire[0:0] mux_1766_nl;
  wire[0:0] or_1766_nl;
  wire[0:0] nand_75_nl;
  wire[0:0] mux_1764_nl;
  wire[0:0] mux_1763_nl;
  wire[0:0] nor_651_nl;
  wire[0:0] nor_652_nl;
  wire[0:0] mux_1762_nl;
  wire[0:0] nor_653_nl;
  wire[0:0] nor_654_nl;
  wire[0:0] mux_1761_nl;
  wire[0:0] mux_1760_nl;
  wire[0:0] mux_1759_nl;
  wire[0:0] or_1755_nl;
  wire[0:0] mux_1758_nl;
  wire[0:0] or_1753_nl;
  wire[0:0] or_1751_nl;
  wire[0:0] or_1750_nl;
  wire[0:0] mux_1757_nl;
  wire[0:0] or_1749_nl;
  wire[0:0] or_1748_nl;
  wire[0:0] or_1747_nl;
  wire[0:0] mux_1756_nl;
  wire[0:0] mux_1755_nl;
  wire[0:0] or_1746_nl;
  wire[0:0] or_1745_nl;
  wire[0:0] or_1743_nl;
  wire[0:0] mux_1822_nl;
  wire[0:0] mux_1821_nl;
  wire[0:0] mux_1820_nl;
  wire[0:0] mux_1819_nl;
  wire[0:0] or_1850_nl;
  wire[0:0] mux_1818_nl;
  wire[0:0] or_1848_nl;
  wire[0:0] mux_1817_nl;
  wire[0:0] or_1847_nl;
  wire[0:0] or_1846_nl;
  wire[0:0] mux_1816_nl;
  wire[0:0] mux_1815_nl;
  wire[0:0] mux_1814_nl;
  wire[0:0] or_1845_nl;
  wire[0:0] or_1843_nl;
  wire[0:0] or_1841_nl;
  wire[0:0] or_1839_nl;
  wire[0:0] mux_1813_nl;
  wire[0:0] mux_1812_nl;
  wire[0:0] mux_1811_nl;
  wire[0:0] mux_1810_nl;
  wire[0:0] or_1838_nl;
  wire[0:0] or_1837_nl;
  wire[0:0] or_1836_nl;
  wire[0:0] or_1835_nl;
  wire[0:0] mux_1809_nl;
  wire[0:0] mux_1808_nl;
  wire[0:0] nand_300_nl;
  wire[0:0] mux_1807_nl;
  wire[0:0] or_1832_nl;
  wire[0:0] or_1831_nl;
  wire[0:0] or_1830_nl;
  wire[0:0] mux_1806_nl;
  wire[0:0] mux_1805_nl;
  wire[0:0] mux_1804_nl;
  wire[0:0] mux_1803_nl;
  wire[0:0] mux_1802_nl;
  wire[0:0] or_1829_nl;
  wire[0:0] or_1827_nl;
  wire[0:0] or_1825_nl;
  wire[0:0] nand_80_nl;
  wire[0:0] mux_1801_nl;
  wire[0:0] mux_1800_nl;
  wire[0:0] mux_1799_nl;
  wire[0:0] or_1823_nl;
  wire[0:0] or_1822_nl;
  wire[0:0] or_1820_nl;
  wire[0:0] or_1819_nl;
  wire[0:0] mux_1798_nl;
  wire[0:0] mux_1797_nl;
  wire[0:0] or_1817_nl;
  wire[0:0] or_1815_nl;
  wire[0:0] mux_1796_nl;
  wire[0:0] or_1814_nl;
  wire[0:0] mux_1795_nl;
  wire[0:0] or_1812_nl;
  wire[0:0] mux_1794_nl;
  wire[0:0] mux_1793_nl;
  wire[0:0] or_1805_nl;
  wire[0:0] or_1804_nl;
  wire[0:0] or_1802_nl;
  wire[0:0] or_1801_nl;
  wire[0:0] mux_1790_nl;
  wire[0:0] or_1800_nl;
  wire[0:0] mux_1789_nl;
  wire[0:0] or_1799_nl;
  wire[0:0] mux_1788_nl;
  wire[0:0] or_1798_nl;
  wire[0:0] or_1797_nl;
  wire[0:0] mux_1855_nl;
  wire[0:0] mux_1854_nl;
  wire[0:0] mux_1853_nl;
  wire[0:0] nand_84_nl;
  wire[0:0] mux_1852_nl;
  wire[0:0] mux_1851_nl;
  wire[0:0] nor_633_nl;
  wire[0:0] nor_634_nl;
  wire[0:0] mux_1850_nl;
  wire[0:0] and_772_nl;
  wire[0:0] and_778_nl;
  wire[0:0] mux_1849_nl;
  wire[0:0] nand_83_nl;
  wire[0:0] mux_1848_nl;
  wire[0:0] nor_637_nl;
  wire[0:0] nor_638_nl;
  wire[0:0] mux_1847_nl;
  wire[0:0] mux_1846_nl;
  wire[0:0] or_1895_nl;
  wire[0:0] or_1893_nl;
  wire[0:0] or_1892_nl;
  wire[0:0] mux_1845_nl;
  wire[0:0] or_1891_nl;
  wire[0:0] mux_1844_nl;
  wire[0:0] mux_1843_nl;
  wire[0:0] nand_291_nl;
  wire[0:0] nand_471_nl;
  wire[0:0] mux_1842_nl;
  wire[0:0] or_1887_nl;
  wire[0:0] or_1885_nl;
  wire[0:0] mux_1841_nl;
  wire[0:0] or_1883_nl;
  wire[0:0] mux_1840_nl;
  wire[0:0] or_1882_nl;
  wire[0:0] or_1881_nl;
  wire[0:0] or_1880_nl;
  wire[0:0] mux_1839_nl;
  wire[0:0] mux_1838_nl;
  wire[0:0] mux_1837_nl;
  wire[0:0] mux_1836_nl;
  wire[0:0] or_1878_nl;
  wire[0:0] mux_1835_nl;
  wire[0:0] mux_1834_nl;
  wire[0:0] or_1875_nl;
  wire[0:0] nand_81_nl;
  wire[0:0] mux_1832_nl;
  wire[0:0] mux_1831_nl;
  wire[0:0] nor_639_nl;
  wire[0:0] nor_640_nl;
  wire[0:0] mux_1830_nl;
  wire[0:0] and_787_nl;
  wire[0:0] and_788_nl;
  wire[0:0] mux_1829_nl;
  wire[0:0] mux_1828_nl;
  wire[0:0] mux_1827_nl;
  wire[0:0] or_1864_nl;
  wire[0:0] mux_1826_nl;
  wire[0:0] or_1862_nl;
  wire[0:0] or_1860_nl;
  wire[0:0] or_1859_nl;
  wire[0:0] mux_1825_nl;
  wire[0:0] or_1858_nl;
  wire[0:0] or_1857_nl;
  wire[0:0] or_1856_nl;
  wire[0:0] mux_1824_nl;
  wire[0:0] mux_1823_nl;
  wire[0:0] nand_296_nl;
  wire[0:0] nand_452_nl;
  wire[0:0] or_1852_nl;
  wire[0:0] mux_1890_nl;
  wire[0:0] mux_1889_nl;
  wire[0:0] mux_1888_nl;
  wire[0:0] mux_1887_nl;
  wire[0:0] or_1956_nl;
  wire[0:0] mux_1886_nl;
  wire[0:0] nand_277_nl;
  wire[0:0] mux_1885_nl;
  wire[0:0] or_1953_nl;
  wire[0:0] or_1952_nl;
  wire[0:0] mux_1884_nl;
  wire[0:0] mux_1883_nl;
  wire[0:0] mux_1882_nl;
  wire[0:0] or_1951_nl;
  wire[0:0] or_1949_nl;
  wire[0:0] or_1947_nl;
  wire[0:0] or_1945_nl;
  wire[0:0] mux_1881_nl;
  wire[0:0] mux_1880_nl;
  wire[0:0] mux_1879_nl;
  wire[0:0] mux_1878_nl;
  wire[0:0] nand_278_nl;
  wire[0:0] nand_279_nl;
  wire[0:0] or_1942_nl;
  wire[0:0] or_1941_nl;
  wire[0:0] mux_1877_nl;
  wire[0:0] mux_1876_nl;
  wire[0:0] nand_280_nl;
  wire[0:0] mux_1875_nl;
  wire[0:0] or_1938_nl;
  wire[0:0] or_1937_nl;
  wire[0:0] or_1936_nl;
  wire[0:0] mux_1874_nl;
  wire[0:0] mux_1873_nl;
  wire[0:0] mux_1872_nl;
  wire[0:0] mux_1871_nl;
  wire[0:0] mux_1870_nl;
  wire[0:0] or_1935_nl;
  wire[0:0] or_1933_nl;
  wire[0:0] or_1931_nl;
  wire[0:0] nand_86_nl;
  wire[0:0] mux_1869_nl;
  wire[0:0] mux_1868_nl;
  wire[0:0] nand_466_nl;
  wire[0:0] mux_1867_nl;
  wire[0:0] nand_283_nl;
  wire[0:0] and_543_nl;
  wire[0:0] nand_462_nl;
  wire[0:0] mux_1866_nl;
  wire[0:0] mux_1865_nl;
  wire[0:0] or_1924_nl;
  wire[0:0] or_1922_nl;
  wire[0:0] mux_1864_nl;
  wire[0:0] or_1921_nl;
  wire[0:0] mux_1863_nl;
  wire[0:0] or_1919_nl;
  wire[0:0] mux_1862_nl;
  wire[0:0] or_1917_nl;
  wire[0:0] mux_1861_nl;
  wire[0:0] and_544_nl;
  wire[0:0] and_545_nl;
  wire[0:0] or_1910_nl;
  wire[0:0] mux_1858_nl;
  wire[0:0] or_1909_nl;
  wire[0:0] mux_1857_nl;
  wire[0:0] or_1908_nl;
  wire[0:0] mux_1856_nl;
  wire[0:0] or_1907_nl;
  wire[0:0] or_1906_nl;
  wire[0:0] mux_1923_nl;
  wire[0:0] mux_1922_nl;
  wire[0:0] mux_1921_nl;
  wire[0:0] nand_90_nl;
  wire[0:0] mux_1920_nl;
  wire[0:0] mux_1919_nl;
  wire[0:0] nor_621_nl;
  wire[0:0] nor_622_nl;
  wire[0:0] mux_1918_nl;
  wire[0:0] nor_623_nl;
  wire[0:0] nor_624_nl;
  wire[0:0] mux_1917_nl;
  wire[0:0] nand_89_nl;
  wire[0:0] mux_1916_nl;
  wire[0:0] nor_625_nl;
  wire[0:0] nor_626_nl;
  wire[0:0] mux_1915_nl;
  wire[0:0] mux_1914_nl;
  wire[0:0] or_2001_nl;
  wire[0:0] or_1999_nl;
  wire[0:0] or_1998_nl;
  wire[0:0] mux_1913_nl;
  wire[0:0] or_1997_nl;
  wire[0:0] mux_1912_nl;
  wire[0:0] mux_1911_nl;
  wire[0:0] or_1996_nl;
  wire[0:0] or_1995_nl;
  wire[0:0] mux_1910_nl;
  wire[0:0] or_1993_nl;
  wire[0:0] or_1991_nl;
  wire[0:0] mux_1909_nl;
  wire[0:0] or_1989_nl;
  wire[0:0] mux_1908_nl;
  wire[0:0] or_1988_nl;
  wire[0:0] or_1987_nl;
  wire[0:0] or_1986_nl;
  wire[0:0] mux_1907_nl;
  wire[0:0] mux_1906_nl;
  wire[0:0] mux_1905_nl;
  wire[0:0] mux_1904_nl;
  wire[0:0] or_1984_nl;
  wire[0:0] mux_1903_nl;
  wire[0:0] mux_1902_nl;
  wire[0:0] or_1981_nl;
  wire[0:0] nand_87_nl;
  wire[0:0] mux_1900_nl;
  wire[0:0] mux_1899_nl;
  wire[0:0] nor_627_nl;
  wire[0:0] nor_628_nl;
  wire[0:0] mux_1898_nl;
  wire[0:0] nor_629_nl;
  wire[0:0] nor_630_nl;
  wire[0:0] mux_1897_nl;
  wire[0:0] mux_1896_nl;
  wire[0:0] mux_1895_nl;
  wire[0:0] or_1970_nl;
  wire[0:0] mux_1894_nl;
  wire[0:0] or_1968_nl;
  wire[0:0] or_1966_nl;
  wire[0:0] or_1965_nl;
  wire[0:0] mux_1893_nl;
  wire[0:0] or_1964_nl;
  wire[0:0] or_1963_nl;
  wire[0:0] or_1962_nl;
  wire[0:0] mux_1892_nl;
  wire[0:0] mux_1891_nl;
  wire[0:0] or_1961_nl;
  wire[0:0] or_1960_nl;
  wire[0:0] or_1958_nl;
  wire[0:0] mux_1958_nl;
  wire[0:0] mux_1957_nl;
  wire[0:0] mux_1956_nl;
  wire[0:0] mux_1955_nl;
  wire[0:0] or_2065_nl;
  wire[0:0] mux_1954_nl;
  wire[0:0] or_2063_nl;
  wire[0:0] mux_1953_nl;
  wire[0:0] or_2062_nl;
  wire[0:0] or_2061_nl;
  wire[0:0] mux_1952_nl;
  wire[0:0] mux_1951_nl;
  wire[0:0] mux_1950_nl;
  wire[0:0] or_2060_nl;
  wire[0:0] or_2058_nl;
  wire[0:0] or_2056_nl;
  wire[0:0] or_2054_nl;
  wire[0:0] mux_1949_nl;
  wire[0:0] mux_1948_nl;
  wire[0:0] mux_1947_nl;
  wire[0:0] mux_1946_nl;
  wire[0:0] or_2053_nl;
  wire[0:0] or_2052_nl;
  wire[0:0] or_2051_nl;
  wire[0:0] or_2050_nl;
  wire[0:0] mux_1945_nl;
  wire[0:0] mux_1944_nl;
  wire[0:0] nand_271_nl;
  wire[0:0] mux_1943_nl;
  wire[0:0] or_2047_nl;
  wire[0:0] or_2046_nl;
  wire[0:0] or_2045_nl;
  wire[0:0] mux_1942_nl;
  wire[0:0] mux_1941_nl;
  wire[0:0] mux_1940_nl;
  wire[0:0] mux_1939_nl;
  wire[0:0] mux_1938_nl;
  wire[0:0] or_2044_nl;
  wire[0:0] or_2042_nl;
  wire[0:0] or_2040_nl;
  wire[0:0] nand_92_nl;
  wire[0:0] mux_1937_nl;
  wire[0:0] mux_1936_nl;
  wire[0:0] mux_1935_nl;
  wire[0:0] or_2038_nl;
  wire[0:0] or_2037_nl;
  wire[0:0] or_2035_nl;
  wire[0:0] or_2034_nl;
  wire[0:0] mux_1934_nl;
  wire[0:0] mux_1933_nl;
  wire[0:0] or_2032_nl;
  wire[0:0] or_2030_nl;
  wire[0:0] mux_1932_nl;
  wire[0:0] or_2029_nl;
  wire[0:0] mux_1931_nl;
  wire[0:0] or_2027_nl;
  wire[0:0] mux_1930_nl;
  wire[0:0] mux_1929_nl;
  wire[0:0] or_2020_nl;
  wire[0:0] or_2019_nl;
  wire[0:0] or_2017_nl;
  wire[0:0] or_2016_nl;
  wire[0:0] mux_1926_nl;
  wire[0:0] or_2015_nl;
  wire[0:0] mux_1925_nl;
  wire[0:0] or_2014_nl;
  wire[0:0] mux_1924_nl;
  wire[0:0] or_2013_nl;
  wire[0:0] or_2012_nl;
  wire[0:0] mux_1991_nl;
  wire[0:0] mux_1990_nl;
  wire[0:0] mux_1989_nl;
  wire[0:0] nand_96_nl;
  wire[0:0] mux_1988_nl;
  wire[0:0] mux_1987_nl;
  wire[0:0] nor_609_nl;
  wire[0:0] nor_610_nl;
  wire[0:0] mux_1986_nl;
  wire[0:0] and_771_nl;
  wire[0:0] and_777_nl;
  wire[0:0] mux_1985_nl;
  wire[0:0] nand_95_nl;
  wire[0:0] mux_1984_nl;
  wire[0:0] nor_613_nl;
  wire[0:0] nor_614_nl;
  wire[0:0] mux_1983_nl;
  wire[0:0] mux_1982_nl;
  wire[0:0] or_2110_nl;
  wire[0:0] or_2108_nl;
  wire[0:0] or_2107_nl;
  wire[0:0] mux_1981_nl;
  wire[0:0] or_2106_nl;
  wire[0:0] mux_1980_nl;
  wire[0:0] mux_1979_nl;
  wire[0:0] nand_262_nl;
  wire[0:0] nand_470_nl;
  wire[0:0] mux_1978_nl;
  wire[0:0] or_2102_nl;
  wire[0:0] or_2100_nl;
  wire[0:0] mux_1977_nl;
  wire[0:0] or_2098_nl;
  wire[0:0] mux_1976_nl;
  wire[0:0] or_2097_nl;
  wire[0:0] or_2096_nl;
  wire[0:0] or_2095_nl;
  wire[0:0] mux_1975_nl;
  wire[0:0] mux_1974_nl;
  wire[0:0] mux_1973_nl;
  wire[0:0] mux_1972_nl;
  wire[0:0] or_2093_nl;
  wire[0:0] mux_1971_nl;
  wire[0:0] mux_1970_nl;
  wire[0:0] or_2090_nl;
  wire[0:0] nand_93_nl;
  wire[0:0] mux_1968_nl;
  wire[0:0] mux_1967_nl;
  wire[0:0] nor_615_nl;
  wire[0:0] nor_616_nl;
  wire[0:0] mux_1966_nl;
  wire[0:0] and_785_nl;
  wire[0:0] and_786_nl;
  wire[0:0] mux_1965_nl;
  wire[0:0] mux_1964_nl;
  wire[0:0] mux_1963_nl;
  wire[0:0] or_2079_nl;
  wire[0:0] mux_1962_nl;
  wire[0:0] or_2077_nl;
  wire[0:0] or_2075_nl;
  wire[0:0] or_2074_nl;
  wire[0:0] mux_1961_nl;
  wire[0:0] or_2073_nl;
  wire[0:0] or_2072_nl;
  wire[0:0] or_2071_nl;
  wire[0:0] mux_1960_nl;
  wire[0:0] mux_1959_nl;
  wire[0:0] nand_267_nl;
  wire[0:0] nand_451_nl;
  wire[0:0] or_2067_nl;
  wire[0:0] mux_2026_nl;
  wire[0:0] mux_2025_nl;
  wire[0:0] mux_2024_nl;
  wire[0:0] mux_2023_nl;
  wire[0:0] or_2171_nl;
  wire[0:0] mux_2022_nl;
  wire[0:0] nand_248_nl;
  wire[0:0] mux_2021_nl;
  wire[0:0] or_2168_nl;
  wire[0:0] or_2167_nl;
  wire[0:0] mux_2020_nl;
  wire[0:0] mux_2019_nl;
  wire[0:0] mux_2018_nl;
  wire[0:0] or_2166_nl;
  wire[0:0] or_2164_nl;
  wire[0:0] or_2162_nl;
  wire[0:0] or_2160_nl;
  wire[0:0] mux_2017_nl;
  wire[0:0] mux_2016_nl;
  wire[0:0] mux_2015_nl;
  wire[0:0] mux_2014_nl;
  wire[0:0] nand_249_nl;
  wire[0:0] nand_250_nl;
  wire[0:0] or_2157_nl;
  wire[0:0] or_2156_nl;
  wire[0:0] mux_2013_nl;
  wire[0:0] mux_2012_nl;
  wire[0:0] nand_251_nl;
  wire[0:0] mux_2011_nl;
  wire[0:0] or_2153_nl;
  wire[0:0] or_2152_nl;
  wire[0:0] or_2151_nl;
  wire[0:0] mux_2010_nl;
  wire[0:0] mux_2009_nl;
  wire[0:0] mux_2008_nl;
  wire[0:0] mux_2007_nl;
  wire[0:0] mux_2006_nl;
  wire[0:0] or_2150_nl;
  wire[0:0] or_2148_nl;
  wire[0:0] or_2146_nl;
  wire[0:0] nand_98_nl;
  wire[0:0] mux_2005_nl;
  wire[0:0] mux_2004_nl;
  wire[0:0] nand_465_nl;
  wire[0:0] mux_2003_nl;
  wire[0:0] nand_254_nl;
  wire[0:0] and_540_nl;
  wire[0:0] nand_461_nl;
  wire[0:0] mux_2002_nl;
  wire[0:0] mux_2001_nl;
  wire[0:0] or_2139_nl;
  wire[0:0] or_2137_nl;
  wire[0:0] mux_2000_nl;
  wire[0:0] or_2136_nl;
  wire[0:0] mux_1999_nl;
  wire[0:0] or_2134_nl;
  wire[0:0] mux_1998_nl;
  wire[0:0] or_2132_nl;
  wire[0:0] mux_1997_nl;
  wire[0:0] and_541_nl;
  wire[0:0] and_542_nl;
  wire[0:0] or_2125_nl;
  wire[0:0] mux_1994_nl;
  wire[0:0] or_2124_nl;
  wire[0:0] mux_1993_nl;
  wire[0:0] or_2123_nl;
  wire[0:0] mux_1992_nl;
  wire[0:0] or_2122_nl;
  wire[0:0] or_2121_nl;
  wire[0:0] mux_2059_nl;
  wire[0:0] mux_2058_nl;
  wire[0:0] mux_2057_nl;
  wire[0:0] nand_102_nl;
  wire[0:0] mux_2056_nl;
  wire[0:0] mux_2055_nl;
  wire[0:0] nor_597_nl;
  wire[0:0] nor_598_nl;
  wire[0:0] mux_2054_nl;
  wire[0:0] and_770_nl;
  wire[0:0] and_776_nl;
  wire[0:0] mux_2053_nl;
  wire[0:0] nand_101_nl;
  wire[0:0] mux_2052_nl;
  wire[0:0] nor_601_nl;
  wire[0:0] nor_602_nl;
  wire[0:0] mux_2051_nl;
  wire[0:0] mux_2050_nl;
  wire[0:0] or_2216_nl;
  wire[0:0] or_2214_nl;
  wire[0:0] or_2213_nl;
  wire[0:0] mux_2049_nl;
  wire[0:0] or_2212_nl;
  wire[0:0] mux_2048_nl;
  wire[0:0] mux_2047_nl;
  wire[0:0] nand_239_nl;
  wire[0:0] nand_469_nl;
  wire[0:0] mux_2046_nl;
  wire[0:0] or_2208_nl;
  wire[0:0] or_2206_nl;
  wire[0:0] mux_2045_nl;
  wire[0:0] or_2204_nl;
  wire[0:0] mux_2044_nl;
  wire[0:0] or_2203_nl;
  wire[0:0] or_2202_nl;
  wire[0:0] or_2201_nl;
  wire[0:0] mux_2043_nl;
  wire[0:0] mux_2042_nl;
  wire[0:0] mux_2041_nl;
  wire[0:0] mux_2040_nl;
  wire[0:0] or_2199_nl;
  wire[0:0] mux_2039_nl;
  wire[0:0] mux_2038_nl;
  wire[0:0] or_2196_nl;
  wire[0:0] nand_99_nl;
  wire[0:0] mux_2036_nl;
  wire[0:0] mux_2035_nl;
  wire[0:0] nor_603_nl;
  wire[0:0] nor_604_nl;
  wire[0:0] mux_2034_nl;
  wire[0:0] and_783_nl;
  wire[0:0] and_784_nl;
  wire[0:0] mux_2033_nl;
  wire[0:0] mux_2032_nl;
  wire[0:0] mux_2031_nl;
  wire[0:0] or_2185_nl;
  wire[0:0] mux_2030_nl;
  wire[0:0] or_2183_nl;
  wire[0:0] or_2181_nl;
  wire[0:0] or_2180_nl;
  wire[0:0] mux_2029_nl;
  wire[0:0] or_2179_nl;
  wire[0:0] or_2178_nl;
  wire[0:0] or_2177_nl;
  wire[0:0] mux_2028_nl;
  wire[0:0] mux_2027_nl;
  wire[0:0] nand_244_nl;
  wire[0:0] nand_450_nl;
  wire[0:0] or_2173_nl;
  wire[0:0] mux_2094_nl;
  wire[0:0] mux_2093_nl;
  wire[0:0] mux_2092_nl;
  wire[0:0] mux_2091_nl;
  wire[0:0] or_2280_nl;
  wire[0:0] mux_2090_nl;
  wire[0:0] nand_222_nl;
  wire[0:0] mux_2089_nl;
  wire[0:0] or_2277_nl;
  wire[0:0] or_2276_nl;
  wire[0:0] mux_2088_nl;
  wire[0:0] mux_2087_nl;
  wire[0:0] mux_2086_nl;
  wire[0:0] or_2275_nl;
  wire[0:0] or_2273_nl;
  wire[0:0] or_2271_nl;
  wire[0:0] or_2269_nl;
  wire[0:0] mux_2085_nl;
  wire[0:0] mux_2084_nl;
  wire[0:0] mux_2083_nl;
  wire[0:0] mux_2082_nl;
  wire[0:0] nand_223_nl;
  wire[0:0] nand_224_nl;
  wire[0:0] or_2266_nl;
  wire[0:0] or_2265_nl;
  wire[0:0] mux_2081_nl;
  wire[0:0] mux_2080_nl;
  wire[0:0] nand_225_nl;
  wire[0:0] mux_2079_nl;
  wire[0:0] or_2262_nl;
  wire[0:0] or_2261_nl;
  wire[0:0] or_2260_nl;
  wire[0:0] mux_2078_nl;
  wire[0:0] mux_2077_nl;
  wire[0:0] mux_2076_nl;
  wire[0:0] mux_2075_nl;
  wire[0:0] mux_2074_nl;
  wire[0:0] or_2259_nl;
  wire[0:0] or_2257_nl;
  wire[0:0] or_2255_nl;
  wire[0:0] nand_104_nl;
  wire[0:0] mux_2073_nl;
  wire[0:0] mux_2072_nl;
  wire[0:0] mux_2071_nl;
  wire[0:0] nand_227_nl;
  wire[0:0] nand_464_nl;
  wire[0:0] nand_229_nl;
  wire[0:0] nand_460_nl;
  wire[0:0] mux_2070_nl;
  wire[0:0] mux_2069_nl;
  wire[0:0] or_2247_nl;
  wire[0:0] or_2245_nl;
  wire[0:0] mux_2068_nl;
  wire[0:0] or_2244_nl;
  wire[0:0] mux_2067_nl;
  wire[0:0] or_2242_nl;
  wire[0:0] mux_2066_nl;
  wire[0:0] mux_2065_nl;
  wire[0:0] nand_233_nl;
  wire[0:0] or_2234_nl;
  wire[0:0] nand_234_nl;
  wire[0:0] or_2231_nl;
  wire[0:0] mux_2062_nl;
  wire[0:0] or_2230_nl;
  wire[0:0] mux_2061_nl;
  wire[0:0] or_2229_nl;
  wire[0:0] mux_2060_nl;
  wire[0:0] or_2228_nl;
  wire[0:0] or_2227_nl;
  wire[0:0] mux_2127_nl;
  wire[0:0] mux_2126_nl;
  wire[0:0] mux_2125_nl;
  wire[0:0] nand_108_nl;
  wire[0:0] mux_2124_nl;
  wire[0:0] mux_2123_nl;
  wire[0:0] and_536_nl;
  wire[0:0] and_537_nl;
  wire[0:0] mux_2122_nl;
  wire[0:0] and_769_nl;
  wire[0:0] and_775_nl;
  wire[0:0] mux_2121_nl;
  wire[0:0] nand_107_nl;
  wire[0:0] mux_2120_nl;
  wire[0:0] nor_591_nl;
  wire[0:0] nor_592_nl;
  wire[0:0] mux_2119_nl;
  wire[0:0] mux_2118_nl;
  wire[0:0] or_2325_nl;
  wire[0:0] or_2323_nl;
  wire[0:0] or_2322_nl;
  wire[0:0] mux_2117_nl;
  wire[0:0] or_2321_nl;
  wire[0:0] mux_2116_nl;
  wire[0:0] mux_2115_nl;
  wire[0:0] nand_208_nl;
  wire[0:0] nand_468_nl;
  wire[0:0] mux_2114_nl;
  wire[0:0] or_2317_nl;
  wire[0:0] or_2315_nl;
  wire[0:0] mux_2113_nl;
  wire[0:0] or_2313_nl;
  wire[0:0] mux_2112_nl;
  wire[0:0] or_2312_nl;
  wire[0:0] or_2311_nl;
  wire[0:0] or_2310_nl;
  wire[0:0] mux_2111_nl;
  wire[0:0] mux_2110_nl;
  wire[0:0] mux_2109_nl;
  wire[0:0] mux_2108_nl;
  wire[0:0] or_2308_nl;
  wire[0:0] mux_2107_nl;
  wire[0:0] mux_2106_nl;
  wire[0:0] or_2305_nl;
  wire[0:0] nand_105_nl;
  wire[0:0] mux_2104_nl;
  wire[0:0] mux_2103_nl;
  wire[0:0] and_538_nl;
  wire[0:0] and_539_nl;
  wire[0:0] mux_2102_nl;
  wire[0:0] and_781_nl;
  wire[0:0] and_782_nl;
  wire[0:0] mux_2101_nl;
  wire[0:0] mux_2100_nl;
  wire[0:0] mux_2099_nl;
  wire[0:0] or_2294_nl;
  wire[0:0] mux_2098_nl;
  wire[0:0] or_2292_nl;
  wire[0:0] nand_215_nl;
  wire[0:0] or_2289_nl;
  wire[0:0] mux_2097_nl;
  wire[0:0] or_2288_nl;
  wire[0:0] or_2287_nl;
  wire[0:0] or_2286_nl;
  wire[0:0] mux_2096_nl;
  wire[0:0] mux_2095_nl;
  wire[0:0] nand_216_nl;
  wire[0:0] nand_449_nl;
  wire[0:0] or_2282_nl;
  wire[0:0] mux_2159_nl;
  wire[0:0] mux_2158_nl;
  wire[0:0] mux_2157_nl;
  wire[0:0] and_530_nl;
  wire[0:0] mux_2156_nl;
  wire[0:0] and_531_nl;
  wire[0:0] mux_2155_nl;
  wire[0:0] nor_570_nl;
  wire[0:0] nor_571_nl;
  wire[0:0] and_532_nl;
  wire[0:0] nor_572_nl;
  wire[0:0] mux_2154_nl;
  wire[0:0] mux_2153_nl;
  wire[0:0] nor_573_nl;
  wire[0:0] mux_2152_nl;
  wire[0:0] mux_2151_nl;
  wire[0:0] or_2835_nl;
  wire[0:0] nand_188_nl;
  wire[0:0] or_2377_nl;
  wire[0:0] mux_2150_nl;
  wire[0:0] mux_2149_nl;
  wire[0:0] and_533_nl;
  wire[0:0] mux_2148_nl;
  wire[0:0] and_766_nl;
  wire[0:0] and_767_nl;
  wire[0:0] nor_576_nl;
  wire[0:0] nor_577_nl;
  wire[0:0] mux_2147_nl;
  wire[0:0] nand_459_nl;
  wire[0:0] mux_2146_nl;
  wire[0:0] or_2365_nl;
  wire[0:0] mux_2145_nl;
  wire[0:0] nand_190_nl;
  wire[0:0] nand_191_nl;
  wire[0:0] mux_2144_nl;
  wire[0:0] mux_2143_nl;
  wire[0:0] mux_2142_nl;
  wire[0:0] nor_578_nl;
  wire[0:0] nor_579_nl;
  wire[0:0] mux_2141_nl;
  wire[0:0] mux_2140_nl;
  wire[0:0] nand_192_nl;
  wire[0:0] nand_193_nl;
  wire[0:0] or_2357_nl;
  wire[0:0] mux_2139_nl;
  wire[0:0] mux_2138_nl;
  wire[0:0] mux_2137_nl;
  wire[0:0] mux_2136_nl;
  wire[0:0] nor_580_nl;
  wire[0:0] nor_581_nl;
  wire[0:0] and_768_nl;
  wire[0:0] and_534_nl;
  wire[0:0] mux_2135_nl;
  wire[0:0] mux_2134_nl;
  wire[0:0] mux_2133_nl;
  wire[0:0] nand_448_nl;
  wire[0:0] nand_422_nl;
  wire[0:0] nand_197_nl;
  wire[0:0] or_2347_nl;
  wire[0:0] mux_2132_nl;
  wire[0:0] nor_583_nl;
  wire[0:0] mux_2131_nl;
  wire[0:0] nor_584_nl;
  wire[0:0] mux_2130_nl;
  wire[0:0] and_774_nl;
  wire[0:0] mux_2129_nl;
  wire[0:0] and_780_nl;
  wire[0:0] mux_2128_nl;
  wire[0:0] and_535_nl;
  wire[0:0] and_791_nl;
  wire[0:0] and_792_nl;
  wire[0:0] mux_2800_nl;
  wire[0:0] or_2913_nl;
  wire[0:0] mux_2799_nl;
  wire[0:0] or_2912_nl;
  wire[0:0] nand_481_nl;
  wire[0:0] mux_nl;
  wire[0:0] or_2999_nl;
  wire[0:0] or_2918_nl;
  wire[0:0] or_2917_nl;
  wire[0:0] mux_2834_nl;
  wire[0:0] mux_2833_nl;
  wire[0:0] nand_484_nl;
  wire[0:0] mux_2832_nl;
  wire[0:0] or_2958_nl;
  wire[0:0] mux_2828_nl;
  wire[0:0] or_2953_nl;
  wire[0:0] mux_2827_nl;
  wire[0:0] mux_2826_nl;
  wire[0:0] or_2952_nl;
  wire[0:0] or_2951_nl;
  wire[0:0] mux_2825_nl;
  wire[0:0] or_2950_nl;
  wire[0:0] or_2949_nl;
  wire[0:0] mux_2824_nl;
  wire[0:0] nand_479_nl;
  wire[0:0] mux_2823_nl;
  wire[0:0] mux_2822_nl;
  wire[0:0] or_2944_nl;
  wire[0:0] or_2943_nl;
  wire[0:0] or_2942_nl;
  wire[0:0] mux_2862_nl;
  wire[0:0] nand_477_nl;
  wire[0:0] mux_2861_nl;
  wire[0:0] mux_2860_nl;
  wire[0:0] or_2996_nl;
  wire[0:0] mux_2856_nl;
  wire[0:0] mux_2855_nl;
  wire[0:0] mux_2854_nl;
  wire[0:0] mux_2853_nl;
  wire[0:0] nand_476_nl;
  wire[0:0] or_2989_nl;
  wire[0:0] or_2987_nl;
  wire[0:0] or_2986_nl;
  wire[0:0] mux_2851_nl;
  wire[0:0] or_2984_nl;
  wire[0:0] nand_475_nl;
  wire[0:0] mux_2850_nl;
  wire[0:0] nor_1007_nl;
  wire[0:0] nor_1008_nl;
  wire[63:0] COMP_LOOP_mux_291_nl;
  wire[63:0] COMP_LOOP_mux1h_842_nl;
  wire[0:0] mux_2897_nl;
  wire[0:0] mux_2898_nl;
  wire[0:0] mux_2899_nl;
  wire[0:0] or_3024_nl;
  wire[0:0] mux_2900_nl;
  wire[0:0] or_3025_nl;
  wire[0:0] mux_2901_nl;
  wire[0:0] nand_491_nl;
  wire[0:0] mux_2902_nl;
  wire[0:0] or_3026_nl;
  wire[9:0] COMP_LOOP_mux_292_nl;
  wire[9:0] COMP_LOOP_mux_293_nl;
  wire[65:0] acc_1_nl;
  wire[66:0] nl_acc_1_nl;
  wire[0:0] operator_64_false_operator_64_false_or_58_nl;
  wire[0:0] operator_64_false_or_130_nl;
  wire[0:0] operator_64_false_operator_64_false_mux_58_nl;
  wire[0:0] operator_64_false_or_131_nl;
  wire[0:0] operator_64_false_operator_64_false_mux_59_nl;
  wire[0:0] operator_64_false_or_132_nl;
  wire[0:0] operator_64_false_operator_64_false_mux_60_nl;
  wire[0:0] operator_64_false_or_133_nl;
  wire[0:0] operator_64_false_operator_64_false_mux_61_nl;
  wire[0:0] operator_64_false_or_134_nl;
  wire[0:0] operator_64_false_operator_64_false_mux_62_nl;
  wire[0:0] operator_64_false_or_135_nl;
  wire[0:0] operator_64_false_operator_64_false_mux_63_nl;
  wire[0:0] operator_64_false_or_136_nl;
  wire[0:0] operator_64_false_operator_64_false_mux_64_nl;
  wire[0:0] operator_64_false_or_137_nl;
  wire[0:0] operator_64_false_operator_64_false_mux_65_nl;
  wire[0:0] operator_64_false_or_138_nl;
  wire[0:0] operator_64_false_operator_64_false_mux_66_nl;
  wire[0:0] operator_64_false_or_139_nl;
  wire[0:0] operator_64_false_operator_64_false_mux_67_nl;
  wire[0:0] operator_64_false_or_140_nl;
  wire[0:0] operator_64_false_operator_64_false_mux_68_nl;
  wire[0:0] operator_64_false_or_141_nl;
  wire[0:0] operator_64_false_operator_64_false_mux_69_nl;
  wire[0:0] operator_64_false_or_142_nl;
  wire[0:0] operator_64_false_operator_64_false_mux_70_nl;
  wire[0:0] operator_64_false_or_143_nl;
  wire[0:0] operator_64_false_operator_64_false_mux_71_nl;
  wire[0:0] operator_64_false_or_144_nl;
  wire[0:0] operator_64_false_operator_64_false_mux_72_nl;
  wire[0:0] operator_64_false_or_145_nl;
  wire[0:0] operator_64_false_operator_64_false_mux_73_nl;
  wire[0:0] operator_64_false_or_146_nl;
  wire[0:0] operator_64_false_operator_64_false_mux_74_nl;
  wire[0:0] operator_64_false_or_147_nl;
  wire[0:0] operator_64_false_operator_64_false_mux_75_nl;
  wire[0:0] operator_64_false_or_148_nl;
  wire[0:0] operator_64_false_operator_64_false_mux_76_nl;
  wire[0:0] operator_64_false_or_149_nl;
  wire[0:0] operator_64_false_operator_64_false_mux_77_nl;
  wire[0:0] operator_64_false_or_150_nl;
  wire[0:0] operator_64_false_operator_64_false_mux_78_nl;
  wire[0:0] operator_64_false_or_151_nl;
  wire[0:0] operator_64_false_operator_64_false_mux_79_nl;
  wire[0:0] operator_64_false_or_152_nl;
  wire[0:0] operator_64_false_operator_64_false_mux_80_nl;
  wire[0:0] operator_64_false_or_153_nl;
  wire[0:0] operator_64_false_operator_64_false_mux_81_nl;
  wire[0:0] operator_64_false_or_154_nl;
  wire[0:0] operator_64_false_operator_64_false_mux_82_nl;
  wire[0:0] operator_64_false_or_155_nl;
  wire[0:0] operator_64_false_operator_64_false_mux_83_nl;
  wire[0:0] operator_64_false_or_156_nl;
  wire[0:0] operator_64_false_operator_64_false_mux_84_nl;
  wire[0:0] operator_64_false_or_157_nl;
  wire[0:0] operator_64_false_operator_64_false_mux_85_nl;
  wire[0:0] operator_64_false_or_158_nl;
  wire[0:0] operator_64_false_operator_64_false_mux_86_nl;
  wire[0:0] operator_64_false_or_159_nl;
  wire[0:0] operator_64_false_operator_64_false_mux_87_nl;
  wire[0:0] operator_64_false_or_160_nl;
  wire[0:0] operator_64_false_operator_64_false_mux_88_nl;
  wire[0:0] operator_64_false_or_161_nl;
  wire[0:0] operator_64_false_operator_64_false_mux_89_nl;
  wire[0:0] operator_64_false_or_162_nl;
  wire[0:0] operator_64_false_operator_64_false_mux_90_nl;
  wire[0:0] operator_64_false_or_163_nl;
  wire[0:0] operator_64_false_operator_64_false_mux_91_nl;
  wire[0:0] operator_64_false_or_164_nl;
  wire[0:0] operator_64_false_operator_64_false_mux_92_nl;
  wire[0:0] operator_64_false_or_165_nl;
  wire[0:0] operator_64_false_operator_64_false_mux_93_nl;
  wire[0:0] operator_64_false_or_166_nl;
  wire[0:0] operator_64_false_operator_64_false_mux_94_nl;
  wire[0:0] operator_64_false_or_167_nl;
  wire[0:0] operator_64_false_operator_64_false_mux_95_nl;
  wire[0:0] operator_64_false_or_168_nl;
  wire[0:0] operator_64_false_operator_64_false_mux_96_nl;
  wire[0:0] operator_64_false_or_169_nl;
  wire[0:0] operator_64_false_operator_64_false_mux_97_nl;
  wire[0:0] operator_64_false_or_170_nl;
  wire[0:0] operator_64_false_operator_64_false_mux_98_nl;
  wire[0:0] operator_64_false_or_171_nl;
  wire[0:0] operator_64_false_operator_64_false_mux_99_nl;
  wire[0:0] operator_64_false_or_172_nl;
  wire[0:0] operator_64_false_operator_64_false_mux_100_nl;
  wire[0:0] operator_64_false_or_173_nl;
  wire[0:0] operator_64_false_operator_64_false_mux_101_nl;
  wire[0:0] operator_64_false_or_174_nl;
  wire[0:0] operator_64_false_operator_64_false_mux_102_nl;
  wire[0:0] operator_64_false_or_175_nl;
  wire[0:0] operator_64_false_operator_64_false_mux_103_nl;
  wire[0:0] operator_64_false_or_176_nl;
  wire[0:0] operator_64_false_operator_64_false_mux_104_nl;
  wire[0:0] operator_64_false_or_177_nl;
  wire[0:0] operator_64_false_operator_64_false_mux_105_nl;
  wire[0:0] operator_64_false_or_178_nl;
  wire[0:0] operator_64_false_operator_64_false_mux_106_nl;
  wire[0:0] operator_64_false_or_179_nl;
  wire[0:0] operator_64_false_operator_64_false_mux_107_nl;
  wire[0:0] operator_64_false_or_180_nl;
  wire[0:0] operator_64_false_operator_64_false_mux_108_nl;
  wire[0:0] operator_64_false_or_181_nl;
  wire[0:0] operator_64_false_operator_64_false_mux_109_nl;
  wire[0:0] operator_64_false_or_182_nl;
  wire[0:0] operator_64_false_operator_64_false_mux_110_nl;
  wire[0:0] operator_64_false_or_183_nl;
  wire[0:0] operator_64_false_operator_64_false_mux_111_nl;
  wire[0:0] operator_64_false_or_184_nl;
  wire[0:0] operator_64_false_operator_64_false_mux_112_nl;
  wire[1:0] operator_64_false_or_185_nl;
  wire[1:0] operator_64_false_operator_64_false_nor_111_nl;
  wire[1:0] operator_64_false_mux1h_62_nl;
  wire[0:0] operator_64_false_or_186_nl;
  wire[6:0] operator_64_false_mux1h_63_nl;
  wire[0:0] operator_64_false_or_187_nl;
  wire[0:0] operator_64_false_or_188_nl;
  wire[0:0] operator_64_false_operator_64_false_or_59_nl;
  wire[1:0] operator_64_false_or_189_nl;
  wire[1:0] operator_64_false_and_65_nl;
  wire[1:0] operator_64_false_operator_64_false_mux_113_nl;
  wire[0:0] operator_64_false_nor_121_nl;
  wire[2:0] operator_64_false_or_190_nl;
  wire[2:0] operator_64_false_and_66_nl;
  wire[2:0] operator_64_false_mux1h_64_nl;
  wire[0:0] operator_64_false_or_191_nl;
  wire[0:0] operator_64_false_or_192_nl;
  wire[0:0] operator_64_false_nor_122_nl;
  wire[0:0] operator_64_false_or_193_nl;
  wire[0:0] operator_64_false_operator_64_false_mux_114_nl;
  wire[0:0] operator_64_false_or_194_nl;
  wire[0:0] operator_64_false_operator_64_false_mux_115_nl;
  wire[0:0] operator_64_false_operator_64_false_or_60_nl;
  wire[0:0] operator_64_false_operator_64_false_or_61_nl;
  wire[64:0] acc_2_nl;
  wire[65:0] nl_acc_2_nl;
  wire[63:0] operator_64_false_mux1h_3_nl;
  wire[0:0] operator_64_false_or_7_nl;
  wire[0:0] operator_64_false_operator_64_false_nand_1_nl;
  wire[63:0] operator_64_false_or_9_nl;
  wire[63:0] operator_64_false_mux1h_4_nl;
  wire[0:0] operator_64_false_or_10_nl;
  wire[0:0] operator_64_false_or_11_nl;
  wire[12:0] acc_3_nl;
  wire[13:0] nl_acc_3_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_3_nl;
  wire[3:0] COMP_LOOP_COMP_LOOP_or_4_nl;
  wire[3:0] COMP_LOOP_and_451_nl;
  wire[0:0] not_7303_nl;
  wire[0:0] COMP_LOOP_or_41_nl;
  wire[5:0] COMP_LOOP_or_42_nl;
  wire[5:0] COMP_LOOP_mux1h_843_nl;
  wire[0:0] COMP_LOOP_or_43_nl;
  wire[2:0] COMP_LOOP_COMP_LOOP_and_992_nl;
  wire[0:0] COMP_LOOP_nor_626_nl;
  wire[1:0] COMP_LOOP_COMP_LOOP_and_993_nl;
  wire[1:0] COMP_LOOP_mux_294_nl;
  wire[0:0] COMP_LOOP_nor_627_nl;
  wire[2:0] COMP_LOOP_and_452_nl;
  wire[2:0] COMP_LOOP_mux1h_844_nl;
  wire[0:0] not_7304_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_5_nl;
  wire[0:0] COMP_LOOP_mux1h_845_nl;
  wire[0:0] COMP_LOOP_mux1h_846_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_994_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_995_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_996_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_997_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_998_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_999_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1000_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1001_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1002_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1003_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1004_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1005_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1006_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1007_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1008_nl;
  wire[0:0] COMP_LOOP_mux1h_847_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1009_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1010_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1011_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1012_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1013_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1014_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1015_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1016_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1017_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1018_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1019_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1020_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1021_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1022_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1023_nl;
  wire[0:0] COMP_LOOP_mux1h_848_nl;
  wire[0:0] COMP_LOOP_mux1h_849_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1024_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1025_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1026_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1027_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1028_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1029_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1030_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1031_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1032_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1033_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1034_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1035_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1036_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1037_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1038_nl;
  wire[0:0] COMP_LOOP_mux1h_850_nl;
  wire[0:0] COMP_LOOP_mux1h_851_nl;
  wire[0:0] COMP_LOOP_mux1h_852_nl;
  wire[0:0] COMP_LOOP_mux1h_853_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1039_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1040_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1041_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1042_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1043_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1044_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1045_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1046_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1047_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1048_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1049_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1050_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1051_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1052_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1053_nl;
  wire[0:0] COMP_LOOP_mux1h_854_nl;
  wire[0:0] COMP_LOOP_mux1h_855_nl;
  wire[0:0] COMP_LOOP_mux1h_856_nl;
  wire[0:0] COMP_LOOP_mux1h_857_nl;
  wire[0:0] COMP_LOOP_mux1h_858_nl;
  wire[0:0] COMP_LOOP_mux1h_859_nl;
  wire[0:0] COMP_LOOP_mux1h_860_nl;

  // Interconnect Declarations for Component Instantiations 
  wire[0:0] mux_2265_nl;
  wire[0:0] mux_2264_nl;
  wire[0:0] mux_2263_nl;
  wire[0:0] nor_556_nl;
  wire[0:0] mux_2262_nl;
  wire[0:0] or_2429_nl;
  wire[0:0] mux_2261_nl;
  wire[0:0] or_2427_nl;
  wire[0:0] or_2426_nl;
  wire[0:0] and_522_nl;
  wire[0:0] mux_2260_nl;
  wire[0:0] nand_457_nl;
  wire[0:0] mux_2259_nl;
  wire[0:0] and_523_nl;
  wire[0:0] mux_2258_nl;
  wire[0:0] or_2422_nl;
  wire[0:0] and_524_nl;
  wire[0:0] mux_2257_nl;
  wire[0:0] or_2418_nl;
  wire[0:0] mux_2256_nl;
  wire[0:0] nor_557_nl;
  wire[0:0] mux_2255_nl;
  wire[0:0] mux_2254_nl;
  wire[0:0] nor_559_nl;
  wire[0:0] mux_2253_nl;
  wire[0:0] or_2409_nl;
  wire [63:0] nl_COMP_LOOP_1_modulo_dev_cmp_base_rsc_dat;
  assign or_2429_nl = (fsm_output[2:0]!=3'b001) | nand_445_cse;
  assign or_2427_nl = (~ (fsm_output[0])) | (~ (fsm_output[2])) | (fsm_output[8])
      | (fsm_output[5]);
  assign or_2426_nl = (fsm_output[0]) | (fsm_output[2]) | nand_445_cse;
  assign mux_2261_nl = MUX_s_1_2_2(or_2427_nl, or_2426_nl, fsm_output[1]);
  assign mux_2262_nl = MUX_s_1_2_2(or_2429_nl, mux_2261_nl, fsm_output[9]);
  assign nor_556_nl = ~((fsm_output[4]) | mux_2262_nl);
  assign nand_457_nl = ~((fsm_output[1]) & (fsm_output[0]) & (fsm_output[2]) & (~
      (fsm_output[8])) & (fsm_output[5]));
  assign mux_2260_nl = MUX_s_1_2_2(or_tmp_2355, nand_457_nl, fsm_output[9]);
  assign and_522_nl = (fsm_output[4]) & (~ mux_2260_nl);
  assign mux_2263_nl = MUX_s_1_2_2(nor_556_nl, and_522_nl, fsm_output[6]);
  assign or_2422_nl = (fsm_output[1]) | (~ (fsm_output[0])) | (~ (fsm_output[2]))
      | (fsm_output[8]) | (~ (fsm_output[5]));
  assign mux_2258_nl = MUX_s_1_2_2(or_2422_nl, or_tmp_2355, fsm_output[9]);
  assign and_523_nl = (fsm_output[4]) & (~ mux_2258_nl);
  assign or_2418_nl = (~ (fsm_output[1])) | (fsm_output[0]) | (fsm_output[2]) | (~
      (fsm_output[8])) | (fsm_output[5]);
  assign mux_2257_nl = MUX_s_1_2_2(or_2418_nl, or_tmp_2352, fsm_output[9]);
  assign and_524_nl = (fsm_output[4]) & (~ mux_2257_nl);
  assign mux_2259_nl = MUX_s_1_2_2(and_523_nl, and_524_nl, fsm_output[6]);
  assign mux_2264_nl = MUX_s_1_2_2(mux_2263_nl, mux_2259_nl, fsm_output[3]);
  assign mux_2255_nl = MUX_s_1_2_2(or_tmp_2352, or_tmp_2348, fsm_output[9]);
  assign nor_557_nl = ~((fsm_output[6]) | (~ (fsm_output[4])) | mux_2255_nl);
  assign or_2409_nl = (fsm_output[1]) | (~ (fsm_output[0])) | (fsm_output[2]) | (fsm_output[8])
      | (~ (fsm_output[5]));
  assign mux_2253_nl = MUX_s_1_2_2(or_tmp_2348, or_2409_nl, fsm_output[9]);
  assign nor_559_nl = ~((fsm_output[4]) | mux_2253_nl);
  assign mux_2254_nl = MUX_s_1_2_2(nor_558_cse, nor_559_nl, fsm_output[6]);
  assign mux_2256_nl = MUX_s_1_2_2(nor_557_nl, mux_2254_nl, fsm_output[3]);
  assign mux_2265_nl = MUX_s_1_2_2(mux_2264_nl, mux_2256_nl, fsm_output[7]);
  assign nl_COMP_LOOP_1_modulo_dev_cmp_base_rsc_dat = MUX_v_64_2_2(z_out_3, COMP_LOOP_10_modExp_dev_1_while_mul_mut,
      mux_2265_nl);
  wire [63:0] nl_COMP_LOOP_1_modulo_dev_cmp_m_rsc_dat;
  assign nl_COMP_LOOP_1_modulo_dev_cmp_m_rsc_dat = p_sva;
  wire[0:0] mux_2291_nl;
  wire[0:0] mux_2290_nl;
  wire[0:0] mux_2289_nl;
  wire[0:0] mux_2288_nl;
  wire[0:0] mux_2287_nl;
  wire[0:0] or_2453_nl;
  wire[0:0] mux_2286_nl;
  wire[0:0] nand_119_nl;
  wire[0:0] mux_2285_nl;
  wire[0:0] or_2452_nl;
  wire[0:0] mux_2284_nl;
  wire[0:0] mux_2283_nl;
  wire[0:0] mux_2282_nl;
  wire[0:0] or_2451_nl;
  wire[0:0] or_2450_nl;
  wire[0:0] mux_2281_nl;
  wire[0:0] mux_2280_nl;
  wire[0:0] mux_2279_nl;
  wire[0:0] mux_2278_nl;
  wire[0:0] mux_2276_nl;
  wire[0:0] or_2449_nl;
  wire[0:0] mux_2275_nl;
  wire[0:0] or_2448_nl;
  wire[0:0] mux_2273_nl;
  wire[0:0] or_2444_nl;
  wire[0:0] mux_2272_nl;
  wire[0:0] or_2443_nl;
  wire[0:0] or_2441_nl;
  wire[0:0] mux_2271_nl;
  wire[0:0] or_2439_nl;
  wire[0:0] mux_2270_nl;
  wire[0:0] mux_2269_nl;
  wire[0:0] or_2435_nl;
  wire [0:0] nl_COMP_LOOP_1_modulo_dev_cmp_ccs_ccore_start_rsc_dat;
  assign or_2453_nl = (fsm_output[7]) | (~ (fsm_output[4])) | (~ (fsm_output[2]))
      | (fsm_output[8]) | (fsm_output[5]);
  assign mux_2287_nl = MUX_s_1_2_2(or_2453_nl, or_2573_cse, fsm_output[1]);
  assign nand_119_nl = ~((fsm_output[4]) & (~ mux_2252_cse));
  assign mux_2286_nl = MUX_s_1_2_2(nand_119_nl, mux_tmp_2226, fsm_output[1]);
  assign mux_2288_nl = MUX_s_1_2_2(mux_2287_nl, mux_2286_nl, fsm_output[9]);
  assign or_2452_nl = (fsm_output[1]) | (~ (fsm_output[7])) | (fsm_output[4]) | (fsm_output[2])
      | (fsm_output[8]) | (fsm_output[5]);
  assign mux_2285_nl = MUX_s_1_2_2(or_tmp_2381, or_2452_nl, fsm_output[9]);
  assign mux_2289_nl = MUX_s_1_2_2(mux_2288_nl, mux_2285_nl, fsm_output[6]);
  assign or_2451_nl = nor_368_cse | mux_2252_cse;
  assign mux_2282_nl = MUX_s_1_2_2(or_2451_nl, mux_tmp_2216, fsm_output[1]);
  assign or_2450_nl = (~ (fsm_output[1])) | (fsm_output[7]) | (fsm_output[4]) | (~
      (fsm_output[2])) | (fsm_output[8]) | (fsm_output[5]);
  assign mux_2283_nl = MUX_s_1_2_2(mux_2282_nl, or_2450_nl, fsm_output[9]);
  assign mux_2284_nl = MUX_s_1_2_2(mux_tmp_2223, mux_2283_nl, fsm_output[6]);
  assign mux_2290_nl = MUX_s_1_2_2(mux_2289_nl, mux_2284_nl, fsm_output[3]);
  assign or_2449_nl = (~ (fsm_output[4])) | (fsm_output[2]) | (~ (fsm_output[8]))
      | (fsm_output[5]);
  assign mux_2276_nl = MUX_s_1_2_2(or_2449_nl, mux_tmp_2215, fsm_output[7]);
  assign mux_2278_nl = MUX_s_1_2_2(mux_tmp_2226, mux_2276_nl, fsm_output[1]);
  assign or_2448_nl = (fsm_output[7]) | (~ (fsm_output[2])) | (fsm_output[8]) | (fsm_output[5]);
  assign mux_2275_nl = MUX_s_1_2_2(or_2448_nl, or_2573_cse, fsm_output[1]);
  assign mux_2279_nl = MUX_s_1_2_2(mux_2278_nl, mux_2275_nl, fsm_output[9]);
  assign mux_2280_nl = MUX_s_1_2_2(mux_2279_nl, mux_tmp_2223, fsm_output[6]);
  assign or_2443_nl = (fsm_output[7]) | (~ (fsm_output[4])) | (~ (fsm_output[2]))
      | (fsm_output[8]) | (~ (fsm_output[5]));
  assign or_2441_nl = nor_368_cse | (~ (fsm_output[2])) | (fsm_output[8]) | (~ (fsm_output[5]));
  assign mux_2272_nl = MUX_s_1_2_2(or_2443_nl, or_2441_nl, fsm_output[1]);
  assign or_2444_nl = (fsm_output[9]) | mux_2272_nl;
  assign or_2439_nl = (fsm_output[1]) | (fsm_output[7]) | (fsm_output[4]) | (~ (fsm_output[2]))
      | (fsm_output[8]) | (fsm_output[5]);
  assign or_2435_nl = (fsm_output[2]) | (fsm_output[8]) | (~ (fsm_output[5]));
  assign mux_2269_nl = MUX_s_1_2_2(or_tmp_2373, or_2435_nl, fsm_output[7]);
  assign mux_2270_nl = MUX_s_1_2_2(mux_2269_nl, mux_tmp_2216, fsm_output[1]);
  assign mux_2271_nl = MUX_s_1_2_2(or_2439_nl, mux_2270_nl, fsm_output[9]);
  assign mux_2273_nl = MUX_s_1_2_2(or_2444_nl, mux_2271_nl, fsm_output[6]);
  assign mux_2281_nl = MUX_s_1_2_2(mux_2280_nl, mux_2273_nl, fsm_output[3]);
  assign mux_2291_nl = MUX_s_1_2_2(mux_2290_nl, mux_2281_nl, fsm_output[0]);
  assign nl_COMP_LOOP_1_modulo_dev_cmp_ccs_ccore_start_rsc_dat = ~ mux_2291_nl;
  wire [3:0] nl_STAGE_MAIN_LOOP_lshift_rg_s;
  assign nl_STAGE_MAIN_LOOP_lshift_rg_s = COMP_LOOP_slc_acc_3_12_1_slc[3:0];
  wire [0:0] nl_inPlaceNTT_DIF_core_wait_dp_inst_ensig_cgo_iro;
  assign nl_inPlaceNTT_DIF_core_wait_dp_inst_ensig_cgo_iro = ~ mux_2240_itm;
  wire [0:0] nl_inPlaceNTT_DIF_core_core_fsm_inst_STAGE_MAIN_LOOP_C_3_tr0;
  assign nl_inPlaceNTT_DIF_core_core_fsm_inst_STAGE_MAIN_LOOP_C_3_tr0 = ~ (z_out_2[64]);
  wire [0:0] nl_inPlaceNTT_DIF_core_core_fsm_inst_STAGE_VEC_LOOP_C_0_tr0;
  assign nl_inPlaceNTT_DIF_core_core_fsm_inst_STAGE_VEC_LOOP_C_0_tr0 = ~ (z_out_2[63]);
  wire [0:0] nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_16_tr0;
  assign nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_16_tr0 = ~ operator_64_false_1_slc_operator_64_false_1_acc_5_itm;
  wire [0:0] nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_45_tr0;
  assign nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_45_tr0 = ~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm;
  wire [0:0] nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_90_tr0;
  assign nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_90_tr0 = ~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm;
  wire [0:0] nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_135_tr0;
  assign nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_135_tr0 = ~ operator_64_false_slc_operator_64_false_acc_1_60_itm;
  wire [0:0] nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_180_tr0;
  assign nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_180_tr0 = ~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm;
  wire [0:0] nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_225_tr0;
  assign nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_225_tr0 = ~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm;
  wire [0:0] nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_270_tr0;
  assign nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_270_tr0 = ~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm;
  wire [0:0] nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_315_tr0;
  assign nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_315_tr0 = ~ operator_64_false_slc_operator_64_false_acc_1_60_itm;
  wire [0:0] nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_360_tr0;
  assign nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_360_tr0 = ~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm;
  wire [0:0] nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_405_tr0;
  assign nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_405_tr0 = ~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm;
  wire [0:0] nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_450_tr0;
  assign nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_450_tr0 = ~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm;
  wire [0:0] nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_495_tr0;
  assign nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_495_tr0 = ~ operator_64_false_slc_operator_64_false_acc_1_60_itm;
  wire [0:0] nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_540_tr0;
  assign nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_540_tr0 = ~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm;
  wire [0:0] nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_585_tr0;
  assign nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_585_tr0 = ~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm;
  wire [0:0] nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_630_tr0;
  assign nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_630_tr0 = ~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm;
  wire [0:0] nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_675_tr0;
  assign nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_675_tr0 = ~ operator_64_false_slc_operator_64_false_acc_1_60_itm;
  wire [0:0] nl_inPlaceNTT_DIF_core_core_fsm_inst_STAGE_VEC_LOOP_C_1_tr0;
  assign nl_inPlaceNTT_DIF_core_core_fsm_inst_STAGE_VEC_LOOP_C_1_tr0 = z_out_1[10];
  wire [0:0] nl_inPlaceNTT_DIF_core_core_fsm_inst_STAGE_MAIN_LOOP_C_4_tr0;
  assign nl_inPlaceNTT_DIF_core_core_fsm_inst_STAGE_MAIN_LOOP_C_4_tr0 = z_out_2[4];
  ccs_in_v1 #(.rscid(32'sd5),
  .width(32'sd64)) p_rsci (
      .dat(p_rsc_dat),
      .idat(p_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd6),
  .width(32'sd64)) r_rsci (
      .dat(r_rsc_dat),
      .idat(r_rsci_idat)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_15_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_15_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_14_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_14_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_13_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_13_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_12_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_12_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_11_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_11_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_10_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_10_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_9_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_9_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_8_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_8_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_7_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_7_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_6_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_6_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_5_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_5_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_4_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_4_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_3_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_3_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_2_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_2_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_1_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_1_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_0_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_0_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) p_rsc_triosy_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(p_rsc_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) r_rsc_triosy_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(r_rsc_triosy_lz)
    );
  modulo_dev  COMP_LOOP_1_modulo_dev_cmp (
      .base_rsc_dat(nl_COMP_LOOP_1_modulo_dev_cmp_base_rsc_dat[63:0]),
      .m_rsc_dat(nl_COMP_LOOP_1_modulo_dev_cmp_m_rsc_dat[63:0]),
      .return_rsc_z(COMP_LOOP_1_modulo_dev_cmp_return_rsc_z),
      .ccs_ccore_start_rsc_dat(nl_COMP_LOOP_1_modulo_dev_cmp_ccs_ccore_start_rsc_dat[0:0]),
      .ccs_ccore_clk(clk),
      .ccs_ccore_srst(rst),
      .ccs_ccore_en(COMP_LOOP_1_modulo_dev_cmp_ccs_ccore_en)
    );
  mgc_rem #(.width_a(32'sd64),
  .width_b(32'sd64),
  .signd(32'sd0)) modExp_dev_while_rem_cmp (
      .a(modExp_dev_while_rem_cmp_a),
      .b(reg_COMP_LOOP_1_modulo_dev_cmp_m_rsc_dat_cse),
      .z(modExp_dev_while_rem_cmp_z)
    );
  mgc_div #(.width_a(32'sd64),
  .width_b(32'sd10),
  .signd(32'sd0)) STAGE_MAIN_LOOP_div_cmp (
      .a(STAGE_MAIN_LOOP_div_cmp_a),
      .b(STAGE_MAIN_LOOP_div_cmp_b),
      .z(STAGE_MAIN_LOOP_div_cmp_z)
    );
  mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd10)) STAGE_MAIN_LOOP_lshift_rg (
      .a(1'b1),
      .s(nl_STAGE_MAIN_LOOP_lshift_rg_s[3:0]),
      .z(STAGE_MAIN_LOOP_lshift_psp_1_sva_mx0w0)
    );
  inPlaceNTT_DIF_core_wait_dp inPlaceNTT_DIF_core_wait_dp_inst (
      .ensig_cgo_iro(nl_inPlaceNTT_DIF_core_wait_dp_inst_ensig_cgo_iro[0:0]),
      .ensig_cgo(reg_ensig_cgo_cse),
      .COMP_LOOP_1_modulo_dev_cmp_ccs_ccore_en(COMP_LOOP_1_modulo_dev_cmp_ccs_ccore_en)
    );
  inPlaceNTT_DIF_core_core_fsm inPlaceNTT_DIF_core_core_fsm_inst (
      .clk(clk),
      .rst(rst),
      .fsm_output(fsm_output),
      .STAGE_MAIN_LOOP_C_3_tr0(nl_inPlaceNTT_DIF_core_core_fsm_inst_STAGE_MAIN_LOOP_C_3_tr0[0:0]),
      .modExp_dev_while_C_11_tr0(COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm),
      .STAGE_VEC_LOOP_C_0_tr0(nl_inPlaceNTT_DIF_core_core_fsm_inst_STAGE_VEC_LOOP_C_0_tr0[0:0]),
      .COMP_LOOP_C_16_tr0(nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_16_tr0[0:0]),
      .COMP_LOOP_1_modExp_dev_1_while_C_11_tr0(COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm),
      .COMP_LOOP_C_45_tr0(nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_45_tr0[0:0]),
      .COMP_LOOP_2_modExp_dev_1_while_C_11_tr0(COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm),
      .COMP_LOOP_C_90_tr0(nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_90_tr0[0:0]),
      .COMP_LOOP_3_modExp_dev_1_while_C_11_tr0(COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm),
      .COMP_LOOP_C_135_tr0(nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_135_tr0[0:0]),
      .COMP_LOOP_4_modExp_dev_1_while_C_11_tr0(COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm),
      .COMP_LOOP_C_180_tr0(nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_180_tr0[0:0]),
      .COMP_LOOP_5_modExp_dev_1_while_C_11_tr0(COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm),
      .COMP_LOOP_C_225_tr0(nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_225_tr0[0:0]),
      .COMP_LOOP_6_modExp_dev_1_while_C_11_tr0(COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm),
      .COMP_LOOP_C_270_tr0(nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_270_tr0[0:0]),
      .COMP_LOOP_7_modExp_dev_1_while_C_11_tr0(COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm),
      .COMP_LOOP_C_315_tr0(nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_315_tr0[0:0]),
      .COMP_LOOP_8_modExp_dev_1_while_C_11_tr0(COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm),
      .COMP_LOOP_C_360_tr0(nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_360_tr0[0:0]),
      .COMP_LOOP_9_modExp_dev_1_while_C_11_tr0(COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm),
      .COMP_LOOP_C_405_tr0(nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_405_tr0[0:0]),
      .COMP_LOOP_10_modExp_dev_1_while_C_11_tr0(COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm),
      .COMP_LOOP_C_450_tr0(nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_450_tr0[0:0]),
      .COMP_LOOP_11_modExp_dev_1_while_C_11_tr0(COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm),
      .COMP_LOOP_C_495_tr0(nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_495_tr0[0:0]),
      .COMP_LOOP_12_modExp_dev_1_while_C_11_tr0(COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm),
      .COMP_LOOP_C_540_tr0(nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_540_tr0[0:0]),
      .COMP_LOOP_13_modExp_dev_1_while_C_11_tr0(COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm),
      .COMP_LOOP_C_585_tr0(nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_585_tr0[0:0]),
      .COMP_LOOP_14_modExp_dev_1_while_C_11_tr0(COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm),
      .COMP_LOOP_C_630_tr0(nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_630_tr0[0:0]),
      .COMP_LOOP_15_modExp_dev_1_while_C_11_tr0(COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm),
      .COMP_LOOP_C_675_tr0(nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_675_tr0[0:0]),
      .COMP_LOOP_16_modExp_dev_1_while_C_11_tr0(COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm),
      .COMP_LOOP_C_720_tr0(COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm),
      .STAGE_VEC_LOOP_C_1_tr0(nl_inPlaceNTT_DIF_core_core_fsm_inst_STAGE_VEC_LOOP_C_1_tr0[0:0]),
      .STAGE_MAIN_LOOP_C_4_tr0(nl_inPlaceNTT_DIF_core_core_fsm_inst_STAGE_MAIN_LOOP_C_4_tr0[0:0])
    );
  assign nand_437_cse = ~(COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm
      & (fsm_output[5]) & (fsm_output[6]) & (~ (fsm_output[3])) & (fsm_output[2]));
  assign mux_1112_cse = MUX_s_1_2_2(or_tmp_669, nand_tmp_19, COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm);
  assign mux_2235_nl = MUX_s_1_2_2(mux_2232_itm, (~ mux_tmp_2129), fsm_output[4]);
  assign mux_2233_nl = MUX_s_1_2_2(mux_2232_itm, (~ mux_tmp_2114), fsm_output[4]);
  assign mux_2231_nl = MUX_s_1_2_2(mux_tmp_2131, mux_tmp_2118, fsm_output[4]);
  assign mux_2234_nl = MUX_s_1_2_2(mux_2233_nl, mux_2231_nl, fsm_output[0]);
  assign mux_2236_nl = MUX_s_1_2_2(mux_2235_nl, mux_2234_nl, fsm_output[1]);
  assign mux_2227_nl = MUX_s_1_2_2(or_2733_cse, (~ or_tmp_2324), fsm_output[9]);
  assign mux_2228_nl = MUX_s_1_2_2(mux_2227_nl, (fsm_output[8]), fsm_output[4]);
  assign mux_2226_nl = MUX_s_1_2_2(mux_tmp_2161, nor_tmp_357, fsm_output[4]);
  assign mux_2229_nl = MUX_s_1_2_2(mux_2228_nl, mux_2226_nl, fsm_output[0]);
  assign mux_2224_nl = MUX_s_1_2_2(mux_tmp_2112, and_679_cse, fsm_output[4]);
  assign mux_2225_nl = MUX_s_1_2_2(mux_2224_nl, mux_tmp_2139, fsm_output[0]);
  assign mux_2230_nl = MUX_s_1_2_2(mux_2229_nl, mux_2225_nl, fsm_output[1]);
  assign mux_2237_nl = MUX_s_1_2_2(mux_2236_nl, mux_2230_nl, fsm_output[5]);
  assign mux_2223_nl = MUX_s_1_2_2(mux_tmp_2142, mux_tmp_2139, fsm_output[5]);
  assign mux_2238_nl = MUX_s_1_2_2(mux_2237_nl, mux_2223_nl, fsm_output[6]);
  assign mux_2221_nl = MUX_s_1_2_2((~ mux_tmp_2135), mux_tmp_2139, fsm_output[5]);
  assign mux_2216_nl = MUX_s_1_2_2(or_2733_cse, (fsm_output[7]), fsm_output[9]);
  assign mux_2217_nl = MUX_s_1_2_2(mux_tmp_2110, mux_2216_nl, fsm_output[4]);
  assign mux_2218_nl = MUX_s_1_2_2(mux_tmp_2142, mux_2217_nl, fsm_output[0]);
  assign mux_2213_nl = MUX_s_1_2_2((~ (fsm_output[7])), (fsm_output[8]), fsm_output[9]);
  assign mux_2214_nl = MUX_s_1_2_2(mux_2213_nl, mux_tmp_2161, fsm_output[4]);
  assign mux_2211_nl = MUX_s_1_2_2(or_tmp_2324, mux_tmp_2112, fsm_output[4]);
  assign mux_2215_nl = MUX_s_1_2_2(mux_2214_nl, mux_2211_nl, fsm_output[0]);
  assign mux_2219_nl = MUX_s_1_2_2(mux_2218_nl, mux_2215_nl, fsm_output[1]);
  assign or_2841_nl = (~ (fsm_output[4])) | (fsm_output[9]);
  assign mux_2208_nl = MUX_s_1_2_2((~ or_tmp_2322), (fsm_output[8]), or_2841_nl);
  assign mux_2209_nl = MUX_s_1_2_2(mux_tmp_2124, mux_2208_nl, fsm_output[0]);
  assign mux_2206_nl = MUX_s_1_2_2(nor_tmp_357, mux_tmp_2110, fsm_output[4]);
  assign mux_2207_nl = MUX_s_1_2_2(mux_2206_nl, mux_tmp_2111, fsm_output[0]);
  assign mux_2210_nl = MUX_s_1_2_2(mux_2209_nl, mux_2207_nl, fsm_output[1]);
  assign mux_2220_nl = MUX_s_1_2_2(mux_2219_nl, mux_2210_nl, fsm_output[5]);
  assign mux_2222_nl = MUX_s_1_2_2(mux_2221_nl, mux_2220_nl, fsm_output[6]);
  assign mux_2239_nl = MUX_s_1_2_2(mux_2238_nl, mux_2222_nl, fsm_output[3]);
  assign or_2392_nl = nor_569_cse | (fsm_output[8]);
  assign mux_2200_nl = MUX_s_1_2_2((~ or_tmp_2322), or_2392_nl, fsm_output[4]);
  assign mux_2198_nl = MUX_s_1_2_2(and_679_cse, (~ (fsm_output[7])), fsm_output[9]);
  assign mux_2199_nl = MUX_s_1_2_2(mux_2198_nl, or_tmp_2324, fsm_output[4]);
  assign mux_2201_nl = MUX_s_1_2_2(mux_2200_nl, mux_2199_nl, fsm_output[0]);
  assign mux_2195_nl = MUX_s_1_2_2((fsm_output[7]), mux_tmp_2112, fsm_output[9]);
  assign mux_2196_nl = MUX_s_1_2_2(mux_2195_nl, or_tmp_2324, fsm_output[4]);
  assign mux_2197_nl = MUX_s_1_2_2(mux_2196_nl, mux_tmp_2135, fsm_output[0]);
  assign mux_2202_nl = MUX_s_1_2_2(mux_2201_nl, mux_2197_nl, fsm_output[1]);
  assign mux_2203_nl = MUX_s_1_2_2((~ mux_2202_nl), mux_tmp_2139, fsm_output[5]);
  assign mux_2191_nl = MUX_s_1_2_2(mux_tmp_2139, mux_tmp_2132, fsm_output[0]);
  assign mux_2189_nl = MUX_s_1_2_2(mux_tmp_2130, mux_tmp_2127, fsm_output[0]);
  assign mux_2192_nl = MUX_s_1_2_2(mux_2191_nl, mux_2189_nl, fsm_output[1]);
  assign mux_2194_nl = MUX_s_1_2_2(mux_tmp_2142, mux_2192_nl, fsm_output[5]);
  assign mux_2204_nl = MUX_s_1_2_2(mux_2203_nl, mux_2194_nl, fsm_output[6]);
  assign mux_2184_nl = MUX_s_1_2_2(mux_tmp_2132, mux_tmp_2130, fsm_output[0]);
  assign mux_2179_nl = MUX_s_1_2_2(mux_tmp_2127, mux_tmp_2124, fsm_output[0]);
  assign mux_2185_nl = MUX_s_1_2_2(mux_2184_nl, mux_2179_nl, fsm_output[1]);
  assign mux_2187_nl = MUX_s_1_2_2((~ mux_tmp_2135), mux_2185_nl, fsm_output[5]);
  assign mux_2170_nl = MUX_s_1_2_2(mux_tmp_2118, mux_tmp_2113, fsm_output[4]);
  assign mux_2167_nl = MUX_s_1_2_2((~ or_tmp_2324), or_tmp_2322, fsm_output[9]);
  assign mux_2168_nl = MUX_s_1_2_2(mux_2167_nl, mux_tmp_2113, fsm_output[4]);
  assign mux_2171_nl = MUX_s_1_2_2(mux_2170_nl, mux_2168_nl, fsm_output[0]);
  assign mux_2166_nl = MUX_s_1_2_2(mux_tmp_2114, mux_tmp_2113, fsm_output[4]);
  assign mux_2172_nl = MUX_s_1_2_2(mux_2171_nl, mux_2166_nl, fsm_output[1]);
  assign mux_2173_nl = MUX_s_1_2_2(mux_2172_nl, mux_tmp_2111, fsm_output[5]);
  assign mux_2188_nl = MUX_s_1_2_2(mux_2187_nl, mux_2173_nl, fsm_output[6]);
  assign mux_2205_nl = MUX_s_1_2_2(mux_2204_nl, mux_2188_nl, fsm_output[3]);
  assign mux_2240_itm = MUX_s_1_2_2(mux_2239_nl, mux_2205_nl, fsm_output[2]);
  assign nor_558_cse = ~((fsm_output[4]) | (fsm_output[9]) | (~ (fsm_output[1]))
      | (~ (fsm_output[0])) | (~ (fsm_output[2])) | (fsm_output[8]) | (~ (fsm_output[5])));
  assign nor_368_cse = ~((fsm_output[7]) | (~ (fsm_output[4])));
  assign and_516_cse = (fsm_output[2:1]==2'b11);
  assign and_515_cse = (fsm_output[1:0]==2'b11);
  assign or_602_cse = (fsm_output[4:3]!=2'b00);
  assign or_2500_cse = (fsm_output[1:0]!=2'b00);
  assign mux_1016_nl = MUX_s_1_2_2((fsm_output[6]), or_307_cse, fsm_output[5]);
  assign mux_1031_cse = MUX_s_1_2_2(mux_1016_nl, or_420_cse, fsm_output[4]);
  assign nand_169_cse = ~((fsm_output[2]) & (fsm_output[5]) & (fsm_output[8]));
  assign or_2573_cse = (fsm_output[4]) | (~ (fsm_output[7])) | (~ (fsm_output[2]))
      | (fsm_output[5]) | (fsm_output[8]);
  assign or_598_cse = (fsm_output[3:2]!=2'b00);
  assign nor_813_cse = ~((fsm_output[9:7]!=3'b000));
  assign and_330_rgt = and_dcpl_294 & and_dcpl_93;
  assign mux_79_cse = MUX_s_1_2_2(and_711_cse, or_165_cse, fsm_output[2]);
  assign nand_490_cse = ~((fsm_output[9:8]==2'b11));
  assign nor_1039_cse = ~((fsm_output[5]) | (fsm_output[6]) | (fsm_output[3]));
  assign or_111_cse = (fsm_output[7:6]!=2'b00);
  assign or_2700_cse = (fsm_output[2:1]!=2'b00);
  assign and_711_cse = (fsm_output[3]) & (fsm_output[6]);
  assign or_165_cse = (fsm_output[3]) | (fsm_output[6]);
  assign and_475_cse = (fsm_output[5]) & (fsm_output[6]) & (fsm_output[8]);
  assign nor_510_cse = ~((fsm_output[5]) | (fsm_output[6]) | (fsm_output[8]));
  assign and_697_cse = (fsm_output[0]) & (fsm_output[2]);
  assign nand_445_cse = ~((fsm_output[5]) & (fsm_output[8]));
  assign and_679_cse = (fsm_output[8:7]==2'b11);
  assign and_756_cse = (fsm_output[8:6]==3'b111);
  assign nor_936_cse = ~((fsm_output[8:6]!=3'b000));
  assign or_307_cse = (fsm_output[2]) | (fsm_output[3]) | (fsm_output[6]);
  assign or_2733_cse = (fsm_output[8:7]!=2'b00);
  assign and_459_cse = (fsm_output[7]) & (fsm_output[9]);
  assign or_420_cse = (fsm_output[6:5]!=2'b00);
  assign and_623_cse = (fsm_output[5:4]==2'b11);
  assign and_613_cse = (fsm_output[6:5]==2'b11);
  assign nor_497_cse = ~((fsm_output[5]) | (fsm_output[6]) | (fsm_output[7]) | (fsm_output[9]));
  assign and_581_cse = (fsm_output[4]) & (fsm_output[0]);
  assign nor_832_cse = ~((fsm_output[4]) | (fsm_output[0]));
  assign nor_1040_cse = ~((fsm_output[0]) | (~ (fsm_output[9])));
  assign or_3018_cse = (~ (fsm_output[0])) | (fsm_output[9]);
  assign nor_569_cse = ~((fsm_output[9]) | (fsm_output[7]));
  assign nl_COMP_LOOP_1_operator_64_false_acc_tmp = STAGE_VEC_LOOP_j_sva_9_0 + conv_u2u_9_10({COMP_LOOP_k_9_4_sva_4_0
      , 4'b0000}) + conv_u2u_9_10(STAGE_MAIN_LOOP_lshift_psp_1_sva[9:1]);
  assign COMP_LOOP_1_operator_64_false_acc_tmp = nl_COMP_LOOP_1_operator_64_false_acc_tmp[9:0];
  assign nl_COMP_LOOP_acc_8_psp_sva_1 = (STAGE_VEC_LOOP_j_sva_9_0[9:2]) + conv_u2u_7_8({COMP_LOOP_k_9_4_sva_4_0
      , 2'b01});
  assign COMP_LOOP_acc_8_psp_sva_1 = nl_COMP_LOOP_acc_8_psp_sva_1[7:0];
  assign nl_COMP_LOOP_acc_cse_4_sva_1 = STAGE_VEC_LOOP_j_sva_9_0 + conv_u2u_9_10({COMP_LOOP_k_9_4_sva_4_0
      , 4'b0011});
  assign COMP_LOOP_acc_cse_4_sva_1 = nl_COMP_LOOP_acc_cse_4_sva_1[9:0];
  assign nl_COMP_LOOP_acc_cse_2_sva_1 = STAGE_VEC_LOOP_j_sva_9_0 + conv_u2u_9_10({COMP_LOOP_k_9_4_sva_4_0
      , 4'b0001});
  assign COMP_LOOP_acc_cse_2_sva_1 = nl_COMP_LOOP_acc_cse_2_sva_1[9:0];
  assign nl_operator_64_false_acc_cse_2_sva_mx0w0 = STAGE_VEC_LOOP_j_sva_9_0 + conv_u2u_9_10({COMP_LOOP_k_9_4_sva_4_0
      , 4'b0001}) + conv_u2u_9_10(STAGE_MAIN_LOOP_lshift_psp_1_sva[9:1]);
  assign operator_64_false_acc_cse_2_sva_mx0w0 = nl_operator_64_false_acc_cse_2_sva_mx0w0[9:0];
  assign nl_operator_64_false_acc_cse_3_sva_mx0w0 = STAGE_VEC_LOOP_j_sva_9_0 + conv_u2u_9_10({COMP_LOOP_k_9_4_sva_4_0
      , 4'b0010}) + conv_u2u_9_10(STAGE_MAIN_LOOP_lshift_psp_1_sva[9:1]);
  assign operator_64_false_acc_cse_3_sva_mx0w0 = nl_operator_64_false_acc_cse_3_sva_mx0w0[9:0];
  assign nl_operator_64_false_acc_cse_4_sva_mx0w0 = STAGE_VEC_LOOP_j_sva_9_0 + conv_u2u_9_10({COMP_LOOP_k_9_4_sva_4_0
      , 4'b0011}) + conv_u2u_9_10(STAGE_MAIN_LOOP_lshift_psp_1_sva[9:1]);
  assign operator_64_false_acc_cse_4_sva_mx0w0 = nl_operator_64_false_acc_cse_4_sva_mx0w0[9:0];
  assign nl_operator_64_false_acc_cse_5_sva_mx0w0 = STAGE_VEC_LOOP_j_sva_9_0 + conv_u2u_9_10({COMP_LOOP_k_9_4_sva_4_0
      , 4'b0100}) + conv_u2u_9_10(STAGE_MAIN_LOOP_lshift_psp_1_sva[9:1]);
  assign operator_64_false_acc_cse_5_sva_mx0w0 = nl_operator_64_false_acc_cse_5_sva_mx0w0[9:0];
  assign nl_operator_64_false_acc_cse_6_sva_mx0w0 = STAGE_VEC_LOOP_j_sva_9_0 + conv_u2u_9_10({COMP_LOOP_k_9_4_sva_4_0
      , 4'b0101}) + conv_u2u_9_10(STAGE_MAIN_LOOP_lshift_psp_1_sva[9:1]);
  assign operator_64_false_acc_cse_6_sva_mx0w0 = nl_operator_64_false_acc_cse_6_sva_mx0w0[9:0];
  assign nl_operator_64_false_acc_cse_7_sva_mx0w0 = STAGE_VEC_LOOP_j_sva_9_0 + conv_u2u_9_10({COMP_LOOP_k_9_4_sva_4_0
      , 4'b0110}) + conv_u2u_9_10(STAGE_MAIN_LOOP_lshift_psp_1_sva[9:1]);
  assign operator_64_false_acc_cse_7_sva_mx0w0 = nl_operator_64_false_acc_cse_7_sva_mx0w0[9:0];
  assign nl_operator_64_false_acc_cse_8_sva_mx0w0 = STAGE_VEC_LOOP_j_sva_9_0 + conv_u2u_9_10({COMP_LOOP_k_9_4_sva_4_0
      , 4'b0111}) + conv_u2u_9_10(STAGE_MAIN_LOOP_lshift_psp_1_sva[9:1]);
  assign operator_64_false_acc_cse_8_sva_mx0w0 = nl_operator_64_false_acc_cse_8_sva_mx0w0[9:0];
  assign nl_operator_64_false_acc_cse_9_sva_mx0w0 = STAGE_VEC_LOOP_j_sva_9_0 + conv_u2u_9_10({COMP_LOOP_k_9_4_sva_4_0
      , 4'b1000}) + conv_u2u_9_10(STAGE_MAIN_LOOP_lshift_psp_1_sva[9:1]);
  assign operator_64_false_acc_cse_9_sva_mx0w0 = nl_operator_64_false_acc_cse_9_sva_mx0w0[9:0];
  assign nl_operator_64_false_acc_cse_10_sva_mx0w0 = STAGE_VEC_LOOP_j_sva_9_0 + conv_u2u_9_10({COMP_LOOP_k_9_4_sva_4_0
      , 4'b1001}) + conv_u2u_9_10(STAGE_MAIN_LOOP_lshift_psp_1_sva[9:1]);
  assign operator_64_false_acc_cse_10_sva_mx0w0 = nl_operator_64_false_acc_cse_10_sva_mx0w0[9:0];
  assign nl_operator_64_false_acc_cse_11_sva_mx0w0 = STAGE_VEC_LOOP_j_sva_9_0 + conv_u2u_9_10({COMP_LOOP_k_9_4_sva_4_0
      , 4'b1010}) + conv_u2u_9_10(STAGE_MAIN_LOOP_lshift_psp_1_sva[9:1]);
  assign operator_64_false_acc_cse_11_sva_mx0w0 = nl_operator_64_false_acc_cse_11_sva_mx0w0[9:0];
  assign nl_operator_64_false_acc_cse_12_sva_mx0w0 = STAGE_VEC_LOOP_j_sva_9_0 + conv_u2u_9_10({COMP_LOOP_k_9_4_sva_4_0
      , 4'b1011}) + conv_u2u_9_10(STAGE_MAIN_LOOP_lshift_psp_1_sva[9:1]);
  assign operator_64_false_acc_cse_12_sva_mx0w0 = nl_operator_64_false_acc_cse_12_sva_mx0w0[9:0];
  assign nl_operator_64_false_acc_cse_13_sva_mx0w0 = STAGE_VEC_LOOP_j_sva_9_0 + conv_u2u_9_10({COMP_LOOP_k_9_4_sva_4_0
      , 4'b1100}) + conv_u2u_9_10(STAGE_MAIN_LOOP_lshift_psp_1_sva[9:1]);
  assign operator_64_false_acc_cse_13_sva_mx0w0 = nl_operator_64_false_acc_cse_13_sva_mx0w0[9:0];
  assign nl_operator_64_false_acc_cse_14_sva_mx0w0 = STAGE_VEC_LOOP_j_sva_9_0 + conv_u2u_9_10({COMP_LOOP_k_9_4_sva_4_0
      , 4'b1101}) + conv_u2u_9_10(STAGE_MAIN_LOOP_lshift_psp_1_sva[9:1]);
  assign operator_64_false_acc_cse_14_sva_mx0w0 = nl_operator_64_false_acc_cse_14_sva_mx0w0[9:0];
  assign nl_operator_64_false_acc_cse_15_sva_mx0w0 = STAGE_VEC_LOOP_j_sva_9_0 + conv_u2u_9_10({COMP_LOOP_k_9_4_sva_4_0
      , 4'b1110}) + conv_u2u_9_10(STAGE_MAIN_LOOP_lshift_psp_1_sva[9:1]);
  assign operator_64_false_acc_cse_15_sva_mx0w0 = nl_operator_64_false_acc_cse_15_sva_mx0w0[9:0];
  assign nl_operator_64_false_acc_cse_sva_mx0w0 = STAGE_VEC_LOOP_j_sva_9_0 + conv_u2u_9_10({COMP_LOOP_k_9_4_sva_4_0
      , 4'b1111}) + conv_u2u_9_10(STAGE_MAIN_LOOP_lshift_psp_1_sva[9:1]);
  assign operator_64_false_acc_cse_sva_mx0w0 = nl_operator_64_false_acc_cse_sva_mx0w0[9:0];
  assign or_tmp = (fsm_output[6:2]!=5'b00000);
  assign nor_tmp_1 = (fsm_output[2]) & (fsm_output[3]) & (fsm_output[6]);
  assign nor_tmp_3 = (fsm_output[9]) & (fsm_output[6]);
  assign and_dcpl = ~((fsm_output[9:8]!=2'b00));
  assign and_dcpl_5 = and_711_cse & (~ (fsm_output[2]));
  assign or_tmp_33 = (fsm_output[3]) | (~ (fsm_output[6]));
  assign or_424_nl = (fsm_output[2]) | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_tmp_79 = MUX_s_1_2_2(or_420_cse, or_424_nl, fsm_output[4]);
  assign nand_442_cse = ~((fsm_output[3:2]==2'b11));
  assign mux_156_cse = MUX_s_1_2_2((~ (fsm_output[6])), (fsm_output[6]), fsm_output[5]);
  assign or_204_cse = (fsm_output[2]) | (fsm_output[6]);
  assign nor_tmp_87 = (fsm_output[8:5]==4'b1111);
  assign mux_tmp_302 = MUX_s_1_2_2(nor_936_cse, and_756_cse, fsm_output[5]);
  assign or_tmp_235 = (fsm_output[8:5]!=4'b0000);
  assign mux_494_cse = MUX_s_1_2_2((~ (fsm_output[9])), (fsm_output[9]), fsm_output[7]);
  assign nor_tmp_130 = (fsm_output[9:8]==2'b11);
  assign and_tmp_11 = (fsm_output[9]) & or_2733_cse;
  assign or_444_nl = (fsm_output[0]) | (fsm_output[6]);
  assign or_533_nl = (~ (fsm_output[0])) | (fsm_output[6]);
  assign mux_792_cse = MUX_s_1_2_2(or_444_nl, or_533_nl, fsm_output[9]);
  assign and_dcpl_44 = (fsm_output[9:8]==2'b01);
  assign and_dcpl_70 = (fsm_output[9:8]==2'b10);
  assign or_2836_nl = (fsm_output[2]) | (fsm_output[5]) | (fsm_output[7]) | (fsm_output[8])
      | (fsm_output[9]);
  assign nand_389_nl = ~((fsm_output[2]) & (fsm_output[5]) & (fsm_output[7]) & (fsm_output[8])
      & (fsm_output[9]));
  assign mux_1048_nl = MUX_s_1_2_2(or_2836_nl, nand_389_nl, or_2500_cse);
  assign nand_390_nl = ~((fsm_output[5]) & (fsm_output[7]) & (fsm_output[8]) & (fsm_output[9]));
  assign mux_1049_nl = MUX_s_1_2_2(mux_1048_nl, nand_390_nl, or_602_cse);
  assign nand_391_nl = ~((fsm_output[9:7]==3'b111));
  assign not_tmp_266 = MUX_s_1_2_2(mux_1049_nl, nand_391_nl, fsm_output[6]);
  assign and_dcpl_91 = (fsm_output[4]) & (~ (fsm_output[0]));
  assign and_dcpl_92 = and_dcpl_91 & (~ (fsm_output[7]));
  assign and_dcpl_93 = and_dcpl_92 & and_dcpl;
  assign and_dcpl_94 = (fsm_output[1]) & (~ (fsm_output[5]));
  assign and_dcpl_95 = ~((fsm_output[3]) | (fsm_output[6]));
  assign and_dcpl_96 = and_dcpl_95 & (~ (fsm_output[2]));
  assign and_dcpl_97 = and_dcpl_96 & and_dcpl_94;
  assign and_dcpl_98 = and_dcpl_97 & and_dcpl_93;
  assign or_tmp_546 = (fsm_output[5]) | (~ (fsm_output[1]));
  assign and_dcpl_105 = nor_832_cse & (~ (fsm_output[7]));
  assign and_dcpl_106 = and_dcpl_105 & and_dcpl;
  assign and_dcpl_109 = and_dcpl_5 & and_dcpl_94;
  assign xor_dcpl = (fsm_output[4]) ^ (fsm_output[0]);
  assign and_dcpl_113 = and_dcpl_5 & xor_dcpl;
  assign nor_809_nl = ~((fsm_output[4]) | (fsm_output[1]) | (~ (fsm_output[2])));
  assign nor_810_nl = ~((~ (fsm_output[4])) | (~ (fsm_output[1])) | (fsm_output[2]));
  assign not_tmp_280 = MUX_s_1_2_2(nor_809_nl, nor_810_nl, fsm_output[0]);
  assign and_dcpl_125 = (fsm_output[2]) & (~ (fsm_output[1])) & (fsm_output[7]) &
      and_dcpl;
  assign and_dcpl_131 = and_623_cse & (fsm_output[7]);
  assign and_dcpl_135 = (fsm_output[3:2]==2'b01);
  assign and_dcpl_143 = (fsm_output[1]) & (fsm_output[5]);
  assign and_dcpl_146 = (fsm_output[3]) & (~ (fsm_output[6]));
  assign and_dcpl_147 = and_dcpl_146 & (fsm_output[2]);
  assign and_dcpl_158 = (~ (fsm_output[1])) & (fsm_output[5]);
  assign and_dcpl_159 = and_dcpl_158 & (~ (fsm_output[4]));
  assign and_741_nl = (fsm_output[0]) & (fsm_output[3]) & (fsm_output[6]);
  assign nor_797_nl = ~((fsm_output[0]) | (fsm_output[6]) | (fsm_output[3]));
  assign not_tmp_292 = MUX_s_1_2_2(and_741_nl, nor_797_nl, fsm_output[7]);
  assign and_dcpl_176 = (fsm_output[2:1]==2'b01);
  assign and_dcpl_192 = ~((fsm_output[1]) | (fsm_output[5]));
  assign and_dcpl_199 = and_dcpl_95 & (fsm_output[2]);
  assign or_tmp_591 = (fsm_output[6]) | (~ (fsm_output[3]));
  assign and_dcpl_225 = and_dcpl_158 & (~ (fsm_output[7])) & nor_tmp_130;
  assign not_tmp_311 = ~((fsm_output[3]) & (fsm_output[6]) & (fsm_output[5]));
  assign not_tmp_312 = ~((fsm_output[6:5]==2'b11));
  assign nor_775_nl = ~((operator_64_false_acc_cse_6_sva[3:0]!=4'b0000) | (fsm_output[3:2]!=2'b01)
      | not_tmp_312);
  assign nor_776_nl = ~((COMP_LOOP_acc_9_psp_sva[2:0]!=3'b000) | (STAGE_VEC_LOOP_j_sva_9_0[0])
      | (fsm_output[3:2]!=2'b01) | not_tmp_312);
  assign mux_1085_nl = MUX_s_1_2_2(nor_775_nl, nor_776_nl, fsm_output[4]);
  assign nand_tmp_16 = ~((fsm_output[8]) & mux_1085_nl);
  assign or_694_cse = (fsm_output[4]) | (STAGE_VEC_LOOP_j_sva_9_0[2:0]!=3'b000) |
      (fsm_output[2]) | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign or_tmp_669 = (fsm_output[6:5]!=2'b01) | nand_442_cse;
  assign or_735_nl = (fsm_output[3:2]!=2'b01);
  assign mux_1111_nl = MUX_s_1_2_2(nand_442_cse, or_735_nl, fsm_output[6]);
  assign nand_tmp_19 = ~((fsm_output[5]) & (~ mux_1111_nl));
  assign not_tmp_322 = ~((fsm_output[6]) & (fsm_output[3]) & (fsm_output[2]));
  assign nor_763_nl = ~((operator_64_false_acc_cse_6_sva[3:0]!=4'b0001) | (fsm_output[3:2]!=2'b01)
      | not_tmp_312);
  assign nor_764_nl = ~((COMP_LOOP_acc_9_psp_sva[2:0]!=3'b000) | (~ (STAGE_VEC_LOOP_j_sva_9_0[0]))
      | (fsm_output[3:2]!=2'b01) | not_tmp_312);
  assign mux_1153_nl = MUX_s_1_2_2(nor_763_nl, nor_764_nl, fsm_output[4]);
  assign nand_tmp_22 = ~((fsm_output[8]) & mux_1153_nl);
  assign or_803_cse = (fsm_output[4]) | (STAGE_VEC_LOOP_j_sva_9_0[2:0]!=3'b001) |
      (fsm_output[2]) | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign nor_751_nl = ~((operator_64_false_acc_cse_6_sva[3:0]!=4'b0010) | (fsm_output[3:2]!=2'b01)
      | not_tmp_312);
  assign nor_752_nl = ~((COMP_LOOP_acc_9_psp_sva[2:0]!=3'b001) | (STAGE_VEC_LOOP_j_sva_9_0[0])
      | (fsm_output[3:2]!=2'b01) | not_tmp_312);
  assign mux_1221_nl = MUX_s_1_2_2(nor_751_nl, nor_752_nl, fsm_output[4]);
  assign nand_tmp_28 = ~((fsm_output[8]) & mux_1221_nl);
  assign or_909_cse = (fsm_output[4]) | (STAGE_VEC_LOOP_j_sva_9_0[2:0]!=3'b010) |
      (fsm_output[2]) | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign nor_739_nl = ~((operator_64_false_acc_cse_6_sva[3:0]!=4'b0011) | (fsm_output[3:2]!=2'b01)
      | not_tmp_312);
  assign nor_740_nl = ~((COMP_LOOP_acc_9_psp_sva[2:0]!=3'b001) | (~ (STAGE_VEC_LOOP_j_sva_9_0[0]))
      | (fsm_output[3:2]!=2'b01) | not_tmp_312);
  assign mux_1289_nl = MUX_s_1_2_2(nor_739_nl, nor_740_nl, fsm_output[4]);
  assign nand_tmp_34 = ~((fsm_output[8]) & mux_1289_nl);
  assign or_1018_cse = (fsm_output[4]) | (STAGE_VEC_LOOP_j_sva_9_0[2:0]!=3'b011)
      | (fsm_output[2]) | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign nor_727_nl = ~((operator_64_false_acc_cse_6_sva[3:0]!=4'b0100) | (fsm_output[3:2]!=2'b01)
      | not_tmp_312);
  assign nor_728_nl = ~((COMP_LOOP_acc_9_psp_sva[2:0]!=3'b010) | (STAGE_VEC_LOOP_j_sva_9_0[0])
      | (fsm_output[3:2]!=2'b01) | not_tmp_312);
  assign mux_1357_nl = MUX_s_1_2_2(nor_727_nl, nor_728_nl, fsm_output[4]);
  assign nand_tmp_40 = ~((fsm_output[8]) & mux_1357_nl);
  assign or_1124_cse = (fsm_output[4]) | (STAGE_VEC_LOOP_j_sva_9_0[2:0]!=3'b100)
      | (fsm_output[2]) | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign nor_715_nl = ~((operator_64_false_acc_cse_6_sva[3:0]!=4'b0101) | (fsm_output[3:2]!=2'b01)
      | not_tmp_312);
  assign nor_716_nl = ~((COMP_LOOP_acc_9_psp_sva[2:0]!=3'b010) | (~ (STAGE_VEC_LOOP_j_sva_9_0[0]))
      | (fsm_output[3:2]!=2'b01) | not_tmp_312);
  assign mux_1425_nl = MUX_s_1_2_2(nor_715_nl, nor_716_nl, fsm_output[4]);
  assign nand_tmp_46 = ~((fsm_output[8]) & mux_1425_nl);
  assign or_1233_cse = (fsm_output[4]) | (STAGE_VEC_LOOP_j_sva_9_0[2:0]!=3'b101)
      | (fsm_output[2]) | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign nor_703_nl = ~((operator_64_false_acc_cse_6_sva[3:0]!=4'b0110) | (fsm_output[3:2]!=2'b01)
      | not_tmp_312);
  assign nor_704_nl = ~((COMP_LOOP_acc_9_psp_sva[2:0]!=3'b011) | (STAGE_VEC_LOOP_j_sva_9_0[0])
      | (fsm_output[3:2]!=2'b01) | not_tmp_312);
  assign mux_1493_nl = MUX_s_1_2_2(nor_703_nl, nor_704_nl, fsm_output[4]);
  assign nand_tmp_52 = ~((fsm_output[8]) & mux_1493_nl);
  assign or_1339_cse = (fsm_output[4]) | (STAGE_VEC_LOOP_j_sva_9_0[2:0]!=3'b110)
      | (fsm_output[2]) | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign nor_691_nl = ~((operator_64_false_acc_cse_6_sva[3:0]!=4'b0111) | (fsm_output[3:2]!=2'b01)
      | not_tmp_312);
  assign nor_692_nl = ~((COMP_LOOP_acc_9_psp_sva[2:0]!=3'b011) | (~ (STAGE_VEC_LOOP_j_sva_9_0[0]))
      | (fsm_output[3:2]!=2'b01) | not_tmp_312);
  assign mux_1561_nl = MUX_s_1_2_2(nor_691_nl, nor_692_nl, fsm_output[4]);
  assign nand_tmp_58 = ~((fsm_output[8]) & mux_1561_nl);
  assign or_1448_cse = (fsm_output[4]) | (STAGE_VEC_LOOP_j_sva_9_0[2:0]!=3'b111)
      | (fsm_output[2]) | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign nor_679_nl = ~((operator_64_false_acc_cse_6_sva[3:0]!=4'b1000) | (fsm_output[3:2]!=2'b01)
      | not_tmp_312);
  assign nor_680_nl = ~((COMP_LOOP_acc_9_psp_sva[2:0]!=3'b100) | (STAGE_VEC_LOOP_j_sva_9_0[0])
      | (fsm_output[3:2]!=2'b01) | not_tmp_312);
  assign mux_1629_nl = MUX_s_1_2_2(nor_679_nl, nor_680_nl, fsm_output[4]);
  assign nand_tmp_64 = ~((fsm_output[8]) & mux_1629_nl);
  assign nor_667_nl = ~((operator_64_false_acc_cse_6_sva[3:0]!=4'b1001) | (fsm_output[3:2]!=2'b01)
      | not_tmp_312);
  assign nor_668_nl = ~((COMP_LOOP_acc_9_psp_sva[2:0]!=3'b100) | (~ (STAGE_VEC_LOOP_j_sva_9_0[0]))
      | (fsm_output[3:2]!=2'b01) | not_tmp_312);
  assign mux_1697_nl = MUX_s_1_2_2(nor_667_nl, nor_668_nl, fsm_output[4]);
  assign nand_tmp_70 = ~((fsm_output[8]) & mux_1697_nl);
  assign nor_655_nl = ~((operator_64_false_acc_cse_6_sva[3:0]!=4'b1010) | (fsm_output[3:2]!=2'b01)
      | not_tmp_312);
  assign nor_656_nl = ~((COMP_LOOP_acc_9_psp_sva[2:0]!=3'b101) | (STAGE_VEC_LOOP_j_sva_9_0[0])
      | (fsm_output[3:2]!=2'b01) | not_tmp_312);
  assign mux_1765_nl = MUX_s_1_2_2(nor_655_nl, nor_656_nl, fsm_output[4]);
  assign nand_tmp_76 = ~((fsm_output[8]) & mux_1765_nl);
  assign nor_643_nl = ~((operator_64_false_acc_cse_6_sva[3:0]!=4'b1011) | (fsm_output[3:2]!=2'b01)
      | not_tmp_312);
  assign nor_644_nl = ~((COMP_LOOP_acc_9_psp_sva[2:0]!=3'b101) | (~ (STAGE_VEC_LOOP_j_sva_9_0[0]))
      | (fsm_output[3:2]!=2'b01) | not_tmp_312);
  assign mux_1833_nl = MUX_s_1_2_2(nor_643_nl, nor_644_nl, fsm_output[4]);
  assign nand_tmp_82 = ~((fsm_output[8]) & mux_1833_nl);
  assign nor_631_nl = ~((operator_64_false_acc_cse_6_sva[3:0]!=4'b1100) | (fsm_output[3:2]!=2'b01)
      | not_tmp_312);
  assign nor_632_nl = ~((COMP_LOOP_acc_9_psp_sva[2:0]!=3'b110) | (STAGE_VEC_LOOP_j_sva_9_0[0])
      | (fsm_output[3:2]!=2'b01) | not_tmp_312);
  assign mux_1901_nl = MUX_s_1_2_2(nor_631_nl, nor_632_nl, fsm_output[4]);
  assign nand_tmp_88 = ~((fsm_output[8]) & mux_1901_nl);
  assign nor_619_nl = ~((operator_64_false_acc_cse_6_sva[3:0]!=4'b1101) | (fsm_output[3:2]!=2'b01)
      | not_tmp_312);
  assign nor_620_nl = ~((COMP_LOOP_acc_9_psp_sva[2:0]!=3'b110) | (~ (STAGE_VEC_LOOP_j_sva_9_0[0]))
      | (fsm_output[3:2]!=2'b01) | not_tmp_312);
  assign mux_1969_nl = MUX_s_1_2_2(nor_619_nl, nor_620_nl, fsm_output[4]);
  assign nand_tmp_94 = ~((fsm_output[8]) & mux_1969_nl);
  assign nor_607_nl = ~((operator_64_false_acc_cse_6_sva[3:0]!=4'b1110) | (fsm_output[3:2]!=2'b01)
      | not_tmp_312);
  assign nor_608_nl = ~((COMP_LOOP_acc_9_psp_sva[2:0]!=3'b111) | (STAGE_VEC_LOOP_j_sva_9_0[0])
      | (fsm_output[3:2]!=2'b01) | not_tmp_312);
  assign mux_2037_nl = MUX_s_1_2_2(nor_607_nl, nor_608_nl, fsm_output[4]);
  assign nand_tmp_100 = ~((fsm_output[8]) & mux_2037_nl);
  assign nor_595_nl = ~((~((operator_64_false_acc_cse_6_sva[3:0]==4'b1111) & (fsm_output[3:2]==2'b01)))
      | not_tmp_312);
  assign nor_596_nl = ~((~((COMP_LOOP_acc_9_psp_sva[2:0]==3'b111) & (STAGE_VEC_LOOP_j_sva_9_0[0])
      & (fsm_output[3:2]==2'b01))) | not_tmp_312);
  assign mux_2105_nl = MUX_s_1_2_2(nor_595_nl, nor_596_nl, fsm_output[4]);
  assign nand_tmp_106 = ~((fsm_output[8]) & mux_2105_nl);
  assign or_tmp_2322 = (fsm_output[8:7]!=2'b10);
  assign mux_tmp_2110 = MUX_s_1_2_2((~ or_tmp_2322), (fsm_output[8]), fsm_output[9]);
  assign mux_tmp_2111 = MUX_s_1_2_2(and_679_cse, mux_tmp_2110, fsm_output[4]);
  assign mux_tmp_2112 = MUX_s_1_2_2((~ (fsm_output[8])), (fsm_output[8]), fsm_output[7]);
  assign mux_tmp_2113 = MUX_s_1_2_2((~ or_2733_cse), mux_tmp_2112, fsm_output[9]);
  assign or_tmp_2324 = (fsm_output[8:7]!=2'b01);
  assign mux_tmp_2114 = MUX_s_1_2_2((~ or_tmp_2324), (fsm_output[7]), fsm_output[9]);
  assign mux_tmp_2118 = MUX_s_1_2_2((~ (fsm_output[8])), or_tmp_2324, fsm_output[9]);
  assign or_2390_nl = (fsm_output[9]) | (~ or_tmp_2322);
  assign mux_2174_nl = MUX_s_1_2_2((~ or_tmp_2322), or_2733_cse, fsm_output[9]);
  assign mux_tmp_2124 = MUX_s_1_2_2(or_2390_nl, mux_2174_nl, fsm_output[4]);
  assign mux_2177_nl = MUX_s_1_2_2((~ and_679_cse), mux_tmp_2112, fsm_output[9]);
  assign mux_2176_nl = MUX_s_1_2_2((~ mux_tmp_2112), (fsm_output[7]), fsm_output[9]);
  assign mux_tmp_2127 = MUX_s_1_2_2(mux_2177_nl, mux_2176_nl, fsm_output[4]);
  assign mux_tmp_2129 = MUX_s_1_2_2((fsm_output[7]), or_tmp_2322, fsm_output[9]);
  assign mux_tmp_2130 = MUX_s_1_2_2(mux_tmp_2113, mux_tmp_2129, fsm_output[4]);
  assign mux_tmp_2131 = MUX_s_1_2_2(or_tmp_2322, and_679_cse, fsm_output[9]);
  assign mux_tmp_2132 = MUX_s_1_2_2(mux_tmp_2113, mux_tmp_2131, fsm_output[4]);
  assign mux_tmp_2135 = MUX_s_1_2_2(mux_tmp_2129, or_tmp_2324, fsm_output[4]);
  assign mux_tmp_2139 = MUX_s_1_2_2(mux_tmp_2113, and_679_cse, fsm_output[4]);
  assign mux_tmp_2142 = MUX_s_1_2_2(mux_tmp_2110, mux_tmp_2114, fsm_output[4]);
  assign nor_tmp_357 = ((fsm_output[9]) | (fsm_output[7])) & (fsm_output[8]);
  assign mux_tmp_2161 = MUX_s_1_2_2(mux_tmp_2112, or_2733_cse, fsm_output[9]);
  assign mux_2232_itm = MUX_s_1_2_2(mux_tmp_2112, and_679_cse, fsm_output[9]);
  assign and_dcpl_239 = and_dcpl_199 & and_dcpl_192;
  assign and_dcpl_240 = and_dcpl_239 & and_dcpl_93;
  assign or_2412_nl = (fsm_output[8]) | (~ (fsm_output[5]));
  assign or_2411_nl = (~ (fsm_output[8])) | (fsm_output[5]);
  assign mux_2252_cse = MUX_s_1_2_2(or_2412_nl, or_2411_nl, fsm_output[2]);
  assign or_tmp_2348 = (fsm_output[1:0]!=2'b00) | mux_2252_cse;
  assign or_tmp_2352 = (~ (fsm_output[1])) | (~ (fsm_output[0])) | (fsm_output[2])
      | (~ (fsm_output[8])) | (fsm_output[5]);
  assign or_tmp_2355 = (~ (fsm_output[1])) | (fsm_output[0]) | (~ (fsm_output[2]))
      | (fsm_output[8]) | (~ (fsm_output[5]));
  assign and_dcpl_241 = (~ (fsm_output[4])) & (fsm_output[0]);
  assign and_dcpl_242 = and_dcpl_241 & (~ (fsm_output[7]));
  assign and_dcpl_243 = and_dcpl_242 & and_dcpl;
  assign and_dcpl_244 = nor_tmp_1 & and_dcpl_192;
  assign and_dcpl_245 = and_dcpl_244 & and_dcpl_243;
  assign and_dcpl_246 = nor_832_cse & (fsm_output[7]);
  assign and_dcpl_248 = and_dcpl_199 & and_dcpl_94;
  assign and_dcpl_249 = and_dcpl_248 & and_dcpl_246 & and_dcpl;
  assign and_dcpl_251 = and_581_cse & (fsm_output[7]);
  assign and_dcpl_252 = and_dcpl_251 & and_dcpl;
  assign and_dcpl_253 = and_dcpl_147 & and_dcpl_143;
  assign and_dcpl_254 = and_dcpl_253 & and_dcpl_252;
  assign and_dcpl_255 = and_dcpl_91 & (fsm_output[7]);
  assign and_dcpl_256 = and_dcpl_255 & and_dcpl;
  assign and_dcpl_257 = and_dcpl_5 & and_dcpl_158;
  assign and_dcpl_258 = and_dcpl_257 & and_dcpl_256;
  assign and_dcpl_259 = and_581_cse & (~ (fsm_output[7]));
  assign and_dcpl_260 = and_dcpl_259 & and_dcpl_44;
  assign and_dcpl_261 = and_dcpl_96 & and_dcpl_158;
  assign and_dcpl_262 = and_dcpl_261 & and_dcpl_260;
  assign and_dcpl_263 = and_dcpl_105 & and_dcpl_44;
  assign and_dcpl_264 = and_dcpl_5 & and_dcpl_143;
  assign and_dcpl_265 = and_dcpl_264 & and_dcpl_263;
  assign and_dcpl_266 = and_dcpl_241 & (fsm_output[7]);
  assign and_dcpl_267 = and_dcpl_266 & and_dcpl_44;
  assign and_dcpl_268 = and_dcpl_96 & and_dcpl_143;
  assign and_dcpl_269 = and_dcpl_268 & and_dcpl_267;
  assign and_dcpl_270 = and_dcpl_255 & and_dcpl_44;
  assign and_dcpl_271 = and_dcpl_244 & and_dcpl_270;
  assign and_dcpl_273 = and_dcpl_239 & and_dcpl_259 & and_dcpl_70;
  assign and_dcpl_275 = nor_tmp_1 & and_dcpl_94;
  assign and_dcpl_276 = and_dcpl_275 & and_dcpl_105 & and_dcpl_70;
  assign and_dcpl_278 = and_dcpl_248 & and_dcpl_266 & and_dcpl_70;
  assign and_dcpl_279 = and_dcpl_246 & and_dcpl_70;
  assign and_dcpl_280 = (~ (fsm_output[3])) & (fsm_output[6]);
  assign and_dcpl_282 = and_dcpl_280 & (~ (fsm_output[2])) & and_dcpl_192;
  assign and_dcpl_283 = and_dcpl_282 & and_dcpl_279;
  assign and_dcpl_284 = and_dcpl_251 & and_dcpl_70;
  assign and_dcpl_285 = and_dcpl_257 & and_dcpl_284;
  assign and_dcpl_286 = and_dcpl_92 & nor_tmp_130;
  assign and_dcpl_287 = and_dcpl_268 & and_dcpl_286;
  assign and_dcpl_288 = and_dcpl_242 & nor_tmp_130;
  assign and_dcpl_289 = and_dcpl_264 & and_dcpl_288;
  assign or_tmp_2368 = (fsm_output[2]) | nand_445_cse;
  assign or_2634_nl = (~ (fsm_output[8])) | (fsm_output[2]) | (fsm_output[5]);
  assign mux_tmp_2215 = MUX_s_1_2_2(or_tmp_2368, or_2634_nl, fsm_output[4]);
  assign or_2431_nl = (~ (fsm_output[4])) | (fsm_output[2]) | (fsm_output[8]) | (fsm_output[5]);
  assign mux_tmp_2216 = MUX_s_1_2_2(mux_tmp_2215, or_2431_nl, fsm_output[7]);
  assign or_tmp_2373 = (fsm_output[4]) | mux_2252_cse;
  assign or_tmp_2381 = (~ (fsm_output[1])) | (fsm_output[7]) | (~ (fsm_output[4]))
      | (~ (fsm_output[2])) | (fsm_output[8]) | (~ (fsm_output[5]));
  assign nand_180_nl = ~((fsm_output[1]) & (fsm_output[7]) & (fsm_output[4]) & (fsm_output[2])
      & (fsm_output[8]) & (fsm_output[5]));
  assign mux_tmp_2223 = MUX_s_1_2_2(nand_180_nl, or_tmp_2381, fsm_output[9]);
  assign mux_tmp_2226 = MUX_s_1_2_2(or_tmp_2368, or_tmp_2373, fsm_output[7]);
  assign and_dcpl_290 = and_dcpl_239 & and_dcpl_243;
  assign or_tmp_2391 = (~ (fsm_output[2])) | (fsm_output[8]) | (fsm_output[7]);
  assign or_tmp_2393 = (fsm_output[2]) | (fsm_output[8]) | (~ (fsm_output[7]));
  assign or_tmp_2395 = (fsm_output[5]) | (fsm_output[8]) | (~ (fsm_output[7]));
  assign or_2464_nl = (~((fsm_output[2:0]!=3'b000))) | (fsm_output[8:7]!=2'b10);
  assign or_2462_nl = ((fsm_output[2:0]==3'b111)) | (fsm_output[8:7]!=2'b00);
  assign mux_tmp_2244 = MUX_s_1_2_2(or_2464_nl, or_2462_nl, fsm_output[5]);
  assign or_tmp_2401 = (~ (fsm_output[2])) | (fsm_output[8]) | (~ (fsm_output[7]));
  assign or_tmp_2402 = (fsm_output[2]) | (~ (fsm_output[8])) | (fsm_output[7]);
  assign mux_tmp_2247 = MUX_s_1_2_2(or_tmp_2402, or_tmp_2401, and_515_cse);
  assign nor_554_cse = ~((fsm_output[2:1]!=2'b00));
  assign or_tmp_2406 = nor_554_cse | (fsm_output[8:7]!=2'b10);
  assign mux_tmp_2250 = MUX_s_1_2_2(or_tmp_2393, or_tmp_2391, or_2500_cse);
  assign not_tmp_572 = ~((fsm_output[8:7]==2'b11));
  assign or_tmp_2409 = (or_2500_cse & (fsm_output[2])) | not_tmp_572;
  assign nor_552_nl = ~((fsm_output[0]) | (~ (fsm_output[2])));
  assign mux_2326_cse = MUX_s_1_2_2(nor_552_nl, and_697_cse, fsm_output[9]);
  assign nand_176_cse = ~((fsm_output[3]) & (fsm_output[6]) & mux_2326_cse);
  assign or_2486_nl = (fsm_output[5]) | nand_176_cse;
  assign or_2484_nl = (~ (fsm_output[5])) | (~ (fsm_output[3])) | (~ (fsm_output[6]))
      | (fsm_output[9]) | (~ (fsm_output[0])) | (fsm_output[2]);
  assign mux_tmp_2276 = MUX_s_1_2_2(or_2486_nl, or_2484_nl, fsm_output[8]);
  assign nor_550_nl = ~((fsm_output[0]) | (fsm_output[2]));
  assign nor_551_nl = ~((~ (fsm_output[0])) | (fsm_output[2]));
  assign mux_2332_cse = MUX_s_1_2_2(nor_550_nl, nor_551_nl, fsm_output[9]);
  assign or_2497_nl = (~ (fsm_output[5])) | (fsm_output[3]) | (fsm_output[6]) | (~
      (fsm_output[9])) | (fsm_output[0]) | (~ (fsm_output[2]));
  assign nand_120_nl = ~((fsm_output[6]) & mux_2332_cse);
  assign or_2492_nl = (fsm_output[6]) | (~ (fsm_output[9])) | (fsm_output[0]) | (fsm_output[2]);
  assign mux_2333_nl = MUX_s_1_2_2(nand_120_nl, or_2492_nl, fsm_output[3]);
  assign or_2495_nl = (fsm_output[5]) | mux_2333_nl;
  assign mux_2334_nl = MUX_s_1_2_2(or_2497_nl, or_2495_nl, fsm_output[8]);
  assign or_2498_nl = (fsm_output[7]) | mux_2334_nl;
  assign or_2491_nl = (fsm_output[8]) | (fsm_output[5]) | (fsm_output[3]) | (fsm_output[6])
      | (fsm_output[9]) | (~ and_697_cse);
  assign mux_2331_nl = MUX_s_1_2_2(mux_tmp_2276, or_2491_nl, fsm_output[7]);
  assign mux_2335_nl = MUX_s_1_2_2(or_2498_nl, mux_2331_nl, fsm_output[4]);
  assign or_2489_nl = (~ (fsm_output[5])) | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[9])
      | (~ (fsm_output[0])) | (fsm_output[2]);
  assign or_2488_nl = (fsm_output[5]) | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[9])
      | (~ and_697_cse);
  assign mux_2328_nl = MUX_s_1_2_2(or_2489_nl, or_2488_nl, fsm_output[8]);
  assign mux_2329_nl = MUX_s_1_2_2(mux_2328_nl, mux_tmp_2276, fsm_output[7]);
  assign nand_175_nl = ~((fsm_output[8]) & (fsm_output[5]) & (fsm_output[3]) & (fsm_output[6])
      & (fsm_output[9]) & (~ (fsm_output[0])) & (~ (fsm_output[2])));
  assign or_2482_nl = (fsm_output[5]) | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[9]))
      | (fsm_output[0]) | (~ (fsm_output[2]));
  assign or_2480_nl = (~ (fsm_output[5])) | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[9])
      | (fsm_output[0]) | (fsm_output[2]);
  assign mux_2324_nl = MUX_s_1_2_2(or_2482_nl, or_2480_nl, fsm_output[8]);
  assign mux_2325_nl = MUX_s_1_2_2(nand_175_nl, mux_2324_nl, fsm_output[7]);
  assign mux_2330_nl = MUX_s_1_2_2(mux_2329_nl, mux_2325_nl, fsm_output[4]);
  assign mux_2336_itm = MUX_s_1_2_2(mux_2335_nl, mux_2330_nl, fsm_output[1]);
  assign and_dcpl_293 = and_dcpl_97 & (~ (fsm_output[4])) & (~ (fsm_output[7])) &
      and_dcpl;
  assign and_dcpl_294 = and_dcpl_96 & and_dcpl_192;
  assign and_dcpl_295 = and_dcpl_294 & and_dcpl_243;
  assign or_tmp_2439 = and_516_cse | (fsm_output[6]) | (fsm_output[3]);
  assign and_tmp_24 = (fsm_output[8:7]==2'b11) & mux_1031_cse;
  assign nor_tmp_388 = (fsm_output[0]) & (fsm_output[6]);
  assign or_tmp_2447 = (~ (fsm_output[2])) | (fsm_output[5]) | (~ (fsm_output[9]))
      | (fsm_output[0]) | (~ (fsm_output[6]));
  assign or_tmp_2451 = (~ (fsm_output[2])) | (fsm_output[5]) | mux_792_cse;
  assign nor_541_nl = ~((fsm_output[3]) | (~ (fsm_output[8])) | (fsm_output[2]) |
      (fsm_output[5]) | (~ (fsm_output[9])) | (fsm_output[0]) | (~ (fsm_output[6])));
  assign nor_542_nl = ~((~ (fsm_output[3])) | (fsm_output[8]) | (~ (fsm_output[2]))
      | (fsm_output[5]) | (fsm_output[9]) | (~ nor_tmp_388));
  assign mux_2357_nl = MUX_s_1_2_2(nor_541_nl, nor_542_nl, fsm_output[7]);
  assign nor_825_nl = ~((fsm_output[0]) | (~ (fsm_output[6])));
  assign mux_2354_nl = MUX_s_1_2_2(nor_825_nl, nor_tmp_388, fsm_output[9]);
  assign or_2521_nl = (fsm_output[2]) | (~((fsm_output[5]) & mux_2354_nl));
  assign mux_2355_nl = MUX_s_1_2_2(or_tmp_2447, or_2521_nl, fsm_output[8]);
  assign and_506_nl = (fsm_output[3]) & (~ mux_2355_nl);
  assign or_2518_nl = (fsm_output[2]) | (~ (fsm_output[5])) | (fsm_output[9]) | (~
      (fsm_output[0])) | (fsm_output[6]);
  assign mux_2353_nl = MUX_s_1_2_2(or_tmp_2451, or_2518_nl, fsm_output[8]);
  assign nor_544_nl = ~((fsm_output[3]) | mux_2353_nl);
  assign mux_2356_nl = MUX_s_1_2_2(and_506_nl, nor_544_nl, fsm_output[7]);
  assign mux_2358_nl = MUX_s_1_2_2(mux_2357_nl, mux_2356_nl, fsm_output[4]);
  assign or_2831_nl = (fsm_output[2]) | (~ (fsm_output[5])) | mux_792_cse;
  assign mux_2350_nl = MUX_s_1_2_2(or_2831_nl, or_tmp_2451, fsm_output[8]);
  assign nor_545_nl = ~((fsm_output[3]) | mux_2350_nl);
  assign or_2510_nl = (fsm_output[2]) | (~ (fsm_output[5])) | (fsm_output[9]) | (fsm_output[0])
      | (~ (fsm_output[6]));
  assign mux_2348_nl = MUX_s_1_2_2(or_tmp_2447, or_2510_nl, fsm_output[8]);
  assign and_507_nl = (fsm_output[3]) & (~ mux_2348_nl);
  assign mux_2351_nl = MUX_s_1_2_2(nor_545_nl, and_507_nl, fsm_output[7]);
  assign nor_546_nl = ~((fsm_output[2]) | (fsm_output[5]) | (fsm_output[9]) | (~
      nor_tmp_388));
  assign nor_547_nl = ~((~ (fsm_output[2])) | (~ (fsm_output[5])) | (fsm_output[9])
      | (~ (fsm_output[0])) | (fsm_output[6]));
  assign mux_2347_nl = MUX_s_1_2_2(nor_546_nl, nor_547_nl, fsm_output[8]);
  assign and_508_nl = (~((fsm_output[7]) | (~ (fsm_output[3])))) & mux_2347_nl;
  assign mux_2352_nl = MUX_s_1_2_2(mux_2351_nl, and_508_nl, fsm_output[4]);
  assign not_tmp_597 = MUX_s_1_2_2(mux_2358_nl, mux_2352_nl, fsm_output[1]);
  assign or_2549_cse = (~ (fsm_output[0])) | (fsm_output[9]) | (fsm_output[5]) |
      (~ (fsm_output[8])) | (fsm_output[2]);
  assign or_2555_nl = (fsm_output[9]) | (~ (fsm_output[5])) | (fsm_output[8]) | (~
      (fsm_output[2]));
  assign nand_420_nl = ~((fsm_output[9]) & (fsm_output[5]) & (~ (fsm_output[8]))
      & (fsm_output[2]));
  assign mux_2374_cse = MUX_s_1_2_2(or_2555_nl, nand_420_nl, fsm_output[0]);
  assign or_2612_nl = (fsm_output[5]) | (fsm_output[1]) | (fsm_output[2]) | (fsm_output[6])
      | (fsm_output[3]);
  assign mux_tmp_2377 = MUX_s_1_2_2(or_420_cse, or_2612_nl, fsm_output[4]);
  assign or_tmp_2548 = (fsm_output[5:4]!=2'b00) | or_tmp_2439;
  assign or_tmp_2549 = (fsm_output[1]) | (fsm_output[2]) | (fsm_output[6]) | (fsm_output[3]);
  assign mux_tmp_2380 = MUX_s_1_2_2(and_dcpl_96, or_tmp_2549, fsm_output[5]);
  assign nor_tmp_399 = or_2700_cse & (fsm_output[6]) & (fsm_output[3]);
  assign mux_tmp_2381 = MUX_s_1_2_2((~ nor_tmp_1), nor_tmp_399, fsm_output[5]);
  assign mux_tmp_2382 = MUX_s_1_2_2(mux_tmp_2381, mux_tmp_2380, fsm_output[4]);
  assign not_tmp_617 = ~((fsm_output[1]) & (fsm_output[2]) & (fsm_output[6]) & (fsm_output[3]));
  assign mux_2439_nl = MUX_s_1_2_2(or_tmp_2439, (~ or_tmp_2549), fsm_output[5]);
  assign mux_2438_nl = MUX_s_1_2_2((~ nor_tmp_399), and_711_cse, fsm_output[5]);
  assign mux_tmp_2389 = MUX_s_1_2_2(mux_2439_nl, mux_2438_nl, fsm_output[4]);
  assign or_tmp_2551 = (fsm_output[5]) | and_dcpl_96;
  assign or_tmp_2552 = (fsm_output[5]) | (~ or_tmp_2439);
  assign mux_tmp_2400 = MUX_s_1_2_2(and_711_cse, or_165_cse, and_516_cse);
  assign nor_tmp_403 = (and_516_cse | (fsm_output[6])) & (fsm_output[3]);
  assign and_dcpl_307 = and_dcpl_266 & and_dcpl;
  assign and_dcpl_311 = and_dcpl_280 & (fsm_output[2]) & and_dcpl_143;
  assign and_dcpl_313 = and_dcpl_92 & and_dcpl_44;
  assign and_dcpl_317 = and_dcpl_246 & and_dcpl_44;
  assign and_dcpl_319 = and_dcpl_251 & and_dcpl_44;
  assign and_dcpl_321 = and_dcpl_92 & and_dcpl_70;
  assign and_dcpl_323 = and_dcpl_242 & and_dcpl_70;
  assign and_dcpl_329 = and_dcpl_259 & nor_tmp_130;
  assign and_dcpl_331 = and_dcpl_105 & nor_tmp_130;
  assign and_dcpl_345 = and_dcpl_248 & and_dcpl_246 & nor_tmp_130;
  assign and_dcpl_346 = and_dcpl_259 & and_dcpl;
  assign mux_tmp_2449 = MUX_s_1_2_2((fsm_output[6]), or_tmp_2549, fsm_output[5]);
  assign mux_tmp_2450 = MUX_s_1_2_2(mux_tmp_2449, or_420_cse, fsm_output[4]);
  assign or_dcpl_72 = or_307_cse | or_tmp_546 | (~ (fsm_output[4])) | (fsm_output[0])
      | (fsm_output[7]) | (fsm_output[8]) | (fsm_output[9]);
  assign mux_tmp_2457 = MUX_s_1_2_2(and_dcpl_95, and_711_cse, fsm_output[2]);
  assign mux_tmp_2458 = MUX_s_1_2_2((~ (fsm_output[3])), (fsm_output[3]), fsm_output[6]);
  assign mux_tmp_2459 = MUX_s_1_2_2(and_dcpl_95, mux_tmp_2458, fsm_output[2]);
  assign mux_2511_nl = MUX_s_1_2_2(mux_tmp_2459, mux_tmp_2457, fsm_output[1]);
  assign or_tmp_2585 = (fsm_output[5]) | mux_2511_nl;
  assign mux_2507_nl = MUX_s_1_2_2(and_dcpl_96, and_711_cse, fsm_output[5]);
  assign mux_tmp_2461 = MUX_s_1_2_2((~ or_tmp_2585), mux_2507_nl, fsm_output[4]);
  assign mux_tmp_2462 = MUX_s_1_2_2(and_dcpl_96, nor_tmp_399, fsm_output[5]);
  assign mux_tmp_2467 = MUX_s_1_2_2(mux_tmp_2458, and_711_cse, fsm_output[2]);
  assign mux_tmp_2468 = MUX_s_1_2_2(mux_tmp_2457, mux_tmp_2467, fsm_output[1]);
  assign or_tmp_2587 = (fsm_output[5]) | mux_tmp_2468;
  assign mux_tmp_2469 = MUX_s_1_2_2(not_tmp_617, or_tmp_2549, fsm_output[5]);
  assign mux_tmp_2470 = MUX_s_1_2_2(mux_tmp_2469, or_tmp_2587, fsm_output[4]);
  assign or_tmp_2588 = (fsm_output[5]) | (~ nor_tmp_1);
  assign mux_2524_nl = MUX_s_1_2_2(mux_tmp_2458, and_711_cse, or_2700_cse);
  assign nand_137_nl = ~((fsm_output[5]) & (~ mux_2524_nl));
  assign mux_tmp_2474 = MUX_s_1_2_2(nand_137_nl, or_tmp_2588, fsm_output[4]);
  assign and_494_nl = or_204_cse & (fsm_output[3]);
  assign mux_2531_nl = MUX_s_1_2_2(mux_tmp_2467, and_494_nl, fsm_output[1]);
  assign nand_tmp_140 = ~((fsm_output[5]) & (~ mux_2531_nl));
  assign nor_tmp_417 = (fsm_output[5]) & (fsm_output[6]) & (fsm_output[8]) & (fsm_output[9]);
  assign nor_516_nl = ~((fsm_output[6]) | (fsm_output[8]) | (fsm_output[9]));
  assign and_489_nl = (fsm_output[6]) & (fsm_output[8]) & (fsm_output[9]);
  assign mux_tmp_2529 = MUX_s_1_2_2(nor_516_nl, and_489_nl, fsm_output[5]);
  assign not_tmp_662 = ~((fsm_output[5]) | (fsm_output[6]) | (fsm_output[8]) | (fsm_output[9]));
  assign mux_2583_nl = MUX_s_1_2_2(not_tmp_662, mux_tmp_2529, or_2700_cse);
  assign mux_2584_nl = MUX_s_1_2_2(not_tmp_662, mux_2583_nl, fsm_output[3]);
  assign mux_2581_nl = MUX_s_1_2_2(mux_tmp_2529, nor_tmp_417, and_515_cse);
  assign mux_2582_nl = MUX_s_1_2_2(mux_2581_nl, nor_tmp_417, or_598_cse);
  assign mux_2585_nl = MUX_s_1_2_2(mux_2584_nl, mux_2582_nl, fsm_output[4]);
  assign mux_2586_itm = MUX_s_1_2_2(mux_2585_nl, nor_tmp_130, fsm_output[7]);
  assign mux_tmp_2538 = MUX_s_1_2_2(mux_tmp_79, mux_tmp_2377, fsm_output[0]);
  assign not_tmp_664 = ~((fsm_output[7]) | mux_tmp_2538);
  assign mux_2607_nl = MUX_s_1_2_2((~ (fsm_output[6])), or_tmp_33, and_516_cse);
  assign mux_2608_nl = MUX_s_1_2_2(mux_2607_nl, (fsm_output[6]), fsm_output[5]);
  assign or_2877_nl = (fsm_output[2]) | (fsm_output[5]);
  assign mux_2606_nl = MUX_s_1_2_2(or_tmp_591, (fsm_output[6]), or_2877_nl);
  assign mux_2609_nl = MUX_s_1_2_2(mux_2608_nl, mux_2606_nl, fsm_output[4]);
  assign mux_2603_nl = MUX_s_1_2_2((~ (fsm_output[6])), or_tmp_33, fsm_output[2]);
  assign mux_2604_nl = MUX_s_1_2_2(mux_2603_nl, (fsm_output[6]), fsm_output[5]);
  assign or_2604_nl = (fsm_output[5]) | (fsm_output[1]) | (fsm_output[2]);
  assign mux_2602_nl = MUX_s_1_2_2(or_tmp_591, (fsm_output[6]), or_2604_nl);
  assign mux_2605_nl = MUX_s_1_2_2(mux_2604_nl, mux_2602_nl, fsm_output[4]);
  assign mux_2610_nl = MUX_s_1_2_2(mux_2609_nl, mux_2605_nl, fsm_output[0]);
  assign and_dcpl_354 = (~ mux_2610_nl) & nor_813_cse;
  assign mux_2613_nl = MUX_s_1_2_2(mux_tmp_2538, (~ or_tmp_2548), fsm_output[7]);
  assign and_dcpl_357 = mux_2613_nl & and_dcpl;
  assign and_483_nl = (fsm_output[0]) & (fsm_output[4]) & (fsm_output[5]) & (fsm_output[1])
      & (fsm_output[2]);
  assign mux_2617_nl = MUX_s_1_2_2((fsm_output[6]), or_165_cse, and_483_nl);
  assign mux_2618_nl = MUX_s_1_2_2(mux_tmp_2538, (~ mux_2617_nl), fsm_output[7]);
  assign and_dcpl_359 = mux_2618_nl & and_dcpl;
  assign nor_tmp_427 = (fsm_output[6:3]==4'b1111);
  assign mux_2622_nl = MUX_s_1_2_2(mux_tmp_2538, (~ nor_tmp_427), fsm_output[7]);
  assign and_dcpl_361 = mux_2622_nl & and_dcpl;
  assign nor_871_nl = ~((fsm_output[8]) | (fsm_output[6]));
  assign and_684_nl = (fsm_output[8]) & (fsm_output[6]);
  assign mux_tmp_2574 = MUX_s_1_2_2(nor_871_nl, and_684_nl, fsm_output[5]);
  assign or_tmp_2638 = and_623_cse | (fsm_output[6]);
  assign mux_tmp_2583 = MUX_s_1_2_2((fsm_output[6]), or_tmp_2549, and_623_cse);
  assign mux_2635_nl = MUX_s_1_2_2(mux_tmp_2583, or_tmp_2638, fsm_output[0]);
  assign or_2712_nl = (fsm_output[7]) | mux_2635_nl;
  assign mux_2636_nl = MUX_s_1_2_2(not_tmp_664, or_2712_nl, fsm_output[8]);
  assign and_dcpl_364 = ~(mux_2636_nl | (fsm_output[9]));
  assign or_2719_nl = (fsm_output[3:2]!=2'b00) | and_515_cse | (fsm_output[6:5]!=2'b00);
  assign mux_2643_nl = MUX_s_1_2_2(or_420_cse, or_2719_nl, fsm_output[4]);
  assign nor_940_nl = ~((fsm_output[7]) | mux_2643_nl);
  assign and_395_nl = (fsm_output[3]) & or_2700_cse & (fsm_output[6:5]==2'b11);
  assign mux_2642_nl = MUX_s_1_2_2(and_395_nl, and_613_cse, fsm_output[4]);
  assign or_2900_nl = (fsm_output[7]) | mux_2642_nl;
  assign mux_2644_nl = MUX_s_1_2_2(nor_940_nl, or_2900_nl, fsm_output[8]);
  assign and_dcpl_367 = ~(mux_2644_nl | (fsm_output[9]));
  assign mux_2650_nl = MUX_s_1_2_2(mux_1031_cse, mux_tmp_2450, fsm_output[0]);
  assign and_400_nl = (fsm_output[7]) & mux_2650_nl;
  assign mux_2651_nl = MUX_s_1_2_2(not_tmp_664, and_400_nl, fsm_output[8]);
  assign and_dcpl_370 = ~(mux_2651_nl | (fsm_output[9]));
  assign not_tmp_696 = ~((fsm_output[8:5]!=4'b0000));
  assign not_tmp_698 = ~((fsm_output[8:7]!=2'b00) | mux_tmp_2538);
  assign mux_2659_nl = MUX_s_1_2_2(nor_tmp_1, (fsm_output[6]), fsm_output[5]);
  assign mux_2660_nl = MUX_s_1_2_2(and_613_cse, mux_2659_nl, fsm_output[4]);
  assign and_403_nl = (fsm_output[7]) & mux_2660_nl;
  assign mux_2661_nl = MUX_s_1_2_2(not_tmp_664, and_403_nl, fsm_output[8]);
  assign and_dcpl_372 = ~(mux_2661_nl | (fsm_output[9]));
  assign mux_tmp_2612 = MUX_s_1_2_2((~ (fsm_output[9])), (fsm_output[9]), fsm_output[6]);
  assign not_tmp_703 = ~((fsm_output[6]) | (fsm_output[9]));
  assign mux_2664_nl = MUX_s_1_2_2(not_tmp_703, mux_tmp_2612, fsm_output[3]);
  assign mux_tmp_2614 = MUX_s_1_2_2(mux_2664_nl, nor_tmp_3, fsm_output[4]);
  assign or_2740_nl = (fsm_output[3:2]!=2'b00) | and_515_cse | (fsm_output[8:5]!=4'b0000);
  assign mux_2674_nl = MUX_s_1_2_2(or_tmp_235, or_2740_nl, fsm_output[4]);
  assign or_2735_nl = (fsm_output[0]) | (fsm_output[1]) | (fsm_output[5]) | (fsm_output[6])
      | (fsm_output[7]) | (fsm_output[8]);
  assign mux_2672_nl = MUX_s_1_2_2(or_tmp_235, or_2735_nl, fsm_output[2]);
  assign or_2737_nl = (fsm_output[3]) | mux_2672_nl;
  assign mux_2673_nl = MUX_s_1_2_2(or_tmp_235, or_2737_nl, fsm_output[4]);
  assign not_tmp_706 = MUX_s_1_2_2(mux_2674_nl, (~ mux_2673_nl), fsm_output[9]);
  assign or_tmp_2668 = (fsm_output[8:6]!=3'b000);
  assign and_tmp_32 = (fsm_output[9]) & or_tmp_2668;
  assign mux_tmp_2625 = MUX_s_1_2_2(and_tmp_11, and_tmp_32, fsm_output[3]);
  assign mux_tmp_2626 = MUX_s_1_2_2((~ or_tmp_2668), or_2733_cse, fsm_output[9]);
  assign or_2747_nl = (fsm_output[3:2]!=2'b00) | and_515_cse | (fsm_output[9]);
  assign mux_2685_nl = MUX_s_1_2_2((fsm_output[9]), or_2747_nl, fsm_output[4]);
  assign and_461_nl = (fsm_output[2]) & (fsm_output[3]) & (fsm_output[1]) & (fsm_output[9]);
  assign mux_2684_nl = MUX_s_1_2_2(and_461_nl, (fsm_output[9]), fsm_output[4]);
  assign mux_2686_nl = MUX_s_1_2_2((~ mux_2685_nl), mux_2684_nl, fsm_output[6]);
  assign mux_2687_nl = MUX_s_1_2_2(mux_2686_nl, nor_tmp_3, fsm_output[5]);
  assign mux_2688_itm = MUX_s_1_2_2(mux_2687_nl, (fsm_output[9]), or_2733_cse);
  assign mux_2698_nl = MUX_s_1_2_2(mux_494_cse, and_459_cse, fsm_output[2]);
  assign mux_2699_nl = MUX_s_1_2_2(nor_569_cse, mux_2698_nl, fsm_output[4]);
  assign mux_2696_nl = MUX_s_1_2_2(nor_569_cse, mux_494_cse, fsm_output[2]);
  assign mux_2697_nl = MUX_s_1_2_2(mux_2696_nl, and_459_cse, fsm_output[4]);
  assign mux_2700_nl = MUX_s_1_2_2(mux_2699_nl, mux_2697_nl, and_515_cse);
  assign mux_2695_nl = MUX_s_1_2_2(mux_494_cse, and_459_cse, fsm_output[4]);
  assign mux_2701_nl = MUX_s_1_2_2(mux_2700_nl, mux_2695_nl, fsm_output[3]);
  assign mux_2702_nl = MUX_s_1_2_2(mux_2701_nl, and_459_cse, or_420_cse);
  assign mux_2703_itm = MUX_s_1_2_2(mux_2702_nl, (fsm_output[9]), fsm_output[8]);
  assign nor_tmp_459 = (fsm_output[6]) & (fsm_output[7]) & (fsm_output[9]);
  assign mux_tmp_2653 = MUX_s_1_2_2(nor_569_cse, and_459_cse, fsm_output[6]);
  assign nor_tmp_463 = (fsm_output[5]) & (fsm_output[6]) & (fsm_output[7]) & (fsm_output[9]);
  assign or_2762_nl = (fsm_output[8]) | ((fsm_output[7:6]==2'b11));
  assign mux_2715_itm = MUX_s_1_2_2(not_tmp_698, or_2762_nl, fsm_output[9]);
  assign nor_tmp_467 = (fsm_output[5]) & (fsm_output[8]) & (fsm_output[9]);
  assign mux_tmp_2666 = MUX_s_1_2_2(and_dcpl, nor_tmp_130, fsm_output[5]);
  assign not_tmp_729 = ~((fsm_output[5]) | (fsm_output[8]) | (fsm_output[9]));
  assign nor_494_nl = ~(and_515_cse | (fsm_output[5]) | (fsm_output[6]) | (fsm_output[7])
      | (fsm_output[9]));
  assign and_444_nl = or_2500_cse & (fsm_output[5]) & (fsm_output[6]) & (fsm_output[7])
      & (fsm_output[9]);
  assign mux_2724_nl = MUX_s_1_2_2(nor_494_nl, and_444_nl, fsm_output[3]);
  assign and_445_nl = (fsm_output[3]) & (fsm_output[5]) & (fsm_output[6]) & (fsm_output[7])
      & (fsm_output[9]);
  assign mux_2725_nl = MUX_s_1_2_2(mux_2724_nl, and_445_nl, fsm_output[2]);
  assign mux_2726_nl = MUX_s_1_2_2(nor_497_cse, mux_2725_nl, fsm_output[4]);
  assign mux_2727_itm = MUX_s_1_2_2(mux_2726_nl, (fsm_output[9]), fsm_output[8]);
  assign and_412_nl = (fsm_output[8]) & ((fsm_output[7]) | mux_tmp_2583);
  assign mux_2734_itm = MUX_s_1_2_2(not_tmp_698, and_412_nl, fsm_output[9]);
  assign mux_2739_nl = MUX_s_1_2_2(not_tmp_662, mux_tmp_2529, fsm_output[3]);
  assign mux_tmp_2689 = MUX_s_1_2_2(mux_2739_nl, nor_tmp_417, fsm_output[4]);
  assign mux_2741_nl = MUX_s_1_2_2(mux_tmp_2529, nor_tmp_417, fsm_output[3]);
  assign mux_2742_nl = MUX_s_1_2_2(not_tmp_662, mux_2741_nl, fsm_output[4]);
  assign mux_2743_nl = MUX_s_1_2_2(mux_2742_nl, mux_tmp_2689, and_515_cse);
  assign mux_2744_nl = MUX_s_1_2_2(mux_2743_nl, mux_tmp_2689, fsm_output[2]);
  assign mux_2745_itm = MUX_s_1_2_2(mux_2744_nl, nor_tmp_130, fsm_output[7]);
  assign and_694_cse = (fsm_output[2]) & (fsm_output[6]);
  assign mux_2762_nl = MUX_s_1_2_2((~ (fsm_output[3])), (fsm_output[3]), and_694_cse);
  assign mux_2763_nl = MUX_s_1_2_2(mux_2762_nl, mux_tmp_2459, fsm_output[1]);
  assign nor_490_nl = ~((fsm_output[5]) | mux_2763_nl);
  assign mux_tmp_2713 = MUX_s_1_2_2(nor_490_nl, mux_tmp_2462, fsm_output[4]);
  assign mux_tmp_2714 = MUX_s_1_2_2(and_dcpl_96, nor_tmp_1, fsm_output[5]);
  assign mux_tmp_2720 = MUX_s_1_2_2(mux_tmp_2459, mux_tmp_2467, fsm_output[1]);
  assign or_tmp_2733 = (fsm_output[5]) | mux_tmp_2720;
  assign or_tmp_2734 = (~ (fsm_output[5])) | (fsm_output[1]) | (fsm_output[2]) |
      (fsm_output[6]) | (fsm_output[3]);
  assign mux_tmp_2721 = MUX_s_1_2_2(or_tmp_2734, or_tmp_2733, fsm_output[4]);
  assign or_tmp_2735 = (fsm_output[5]) | mux_tmp_2459;
  assign or_tmp_2736 = (fsm_output[5]) | not_tmp_617;
  assign nand_145_nl = ~((fsm_output[5]) & (~ mux_tmp_2467));
  assign mux_tmp_2724 = MUX_s_1_2_2(nand_145_nl, or_tmp_2736, fsm_output[4]);
  assign mux_2782_nl = MUX_s_1_2_2((~ (fsm_output[3])), (fsm_output[3]), or_204_cse);
  assign mux_2783_nl = MUX_s_1_2_2(mux_tmp_2467, mux_2782_nl, fsm_output[1]);
  assign nand_tmp_148 = ~((fsm_output[5]) & (~ mux_2783_nl));
  assign mux_2793_nl = MUX_s_1_2_2(nand_tmp_148, or_tmp_2588, fsm_output[4]);
  assign mux_2794_nl = MUX_s_1_2_2(mux_tmp_2724, mux_2793_nl, fsm_output[0]);
  assign mux_2791_nl = MUX_s_1_2_2(or_tmp_2736, or_tmp_2733, fsm_output[4]);
  assign mux_2792_nl = MUX_s_1_2_2(mux_tmp_2721, mux_2791_nl, fsm_output[0]);
  assign mux_2795_nl = MUX_s_1_2_2(mux_2794_nl, mux_2792_nl, fsm_output[7]);
  assign mux_2787_nl = MUX_s_1_2_2((~ or_tmp_2549), nor_tmp_399, fsm_output[5]);
  assign mux_2788_nl = MUX_s_1_2_2((~ or_tmp_2735), mux_2787_nl, fsm_output[4]);
  assign mux_2789_nl = MUX_s_1_2_2(mux_tmp_2713, mux_2788_nl, fsm_output[0]);
  assign mux_2784_nl = MUX_s_1_2_2(or_tmp_2439, (~ nor_tmp_1), fsm_output[5]);
  assign mux_2785_nl = MUX_s_1_2_2(mux_2784_nl, nand_tmp_148, fsm_output[4]);
  assign mux_2780_nl = MUX_s_1_2_2(mux_tmp_2467, mux_79_cse, fsm_output[1]);
  assign nand_147_nl = ~((fsm_output[5]) & (~ mux_2780_nl));
  assign mux_2781_nl = MUX_s_1_2_2((~ mux_tmp_2714), nand_147_nl, fsm_output[4]);
  assign mux_2786_nl = MUX_s_1_2_2(mux_2785_nl, mux_2781_nl, fsm_output[0]);
  assign mux_2790_nl = MUX_s_1_2_2((~ mux_2789_nl), mux_2786_nl, fsm_output[7]);
  assign mux_2796_nl = MUX_s_1_2_2(mux_2795_nl, mux_2790_nl, fsm_output[8]);
  assign nand_146_nl = ~((fsm_output[5]) & (~ mux_tmp_2720));
  assign mux_2776_nl = MUX_s_1_2_2(nand_146_nl, or_tmp_2736, fsm_output[4]);
  assign mux_2777_nl = MUX_s_1_2_2(mux_2776_nl, mux_tmp_2724, fsm_output[0]);
  assign mux_2773_nl = MUX_s_1_2_2(or_tmp_2734, or_tmp_2735, fsm_output[4]);
  assign mux_2774_nl = MUX_s_1_2_2(mux_2773_nl, mux_tmp_2721, fsm_output[0]);
  assign mux_2778_nl = MUX_s_1_2_2(mux_2777_nl, mux_2774_nl, fsm_output[7]);
  assign mux_2767_nl = MUX_s_1_2_2((~ mux_79_cse), mux_tmp_2459, fsm_output[1]);
  assign nor_489_nl = ~((fsm_output[5]) | mux_2767_nl);
  assign mux_2768_nl = MUX_s_1_2_2(nor_489_nl, mux_tmp_2714, fsm_output[4]);
  assign mux_2769_nl = MUX_s_1_2_2(mux_2768_nl, mux_tmp_2713, fsm_output[0]);
  assign mux_2770_nl = MUX_s_1_2_2((~ mux_2769_nl), or_tmp_2548, fsm_output[7]);
  assign mux_2779_nl = MUX_s_1_2_2(mux_2778_nl, mux_2770_nl, fsm_output[8]);
  assign mux_2797_itm = MUX_s_1_2_2(mux_2796_nl, mux_2779_nl, fsm_output[9]);
  assign and_504_nl = (fsm_output[3]) & (fsm_output[6]) & (~ (fsm_output[0])) & (fsm_output[9])
      & (~ mux_2252_cse);
  assign or_2547_nl = (fsm_output[9]) | mux_2252_cse;
  assign nand_126_nl = ~((fsm_output[9]) & (~ mux_2252_cse));
  assign mux_2369_nl = MUX_s_1_2_2(or_2547_nl, nand_126_nl, fsm_output[0]);
  assign nor_534_nl = ~((fsm_output[3]) | (fsm_output[6]) | mux_2369_nl);
  assign mux_2370_nl = MUX_s_1_2_2(and_504_nl, nor_534_nl, fsm_output[7]);
  assign nor_535_nl = ~((~ (fsm_output[0])) | (fsm_output[9]) | nand_169_cse);
  assign nor_536_nl = ~((~ (fsm_output[0])) | (fsm_output[9]) | (fsm_output[2]) |
      (fsm_output[8]) | (fsm_output[5]));
  assign mux_2367_nl = MUX_s_1_2_2(nor_535_nl, nor_536_nl, fsm_output[6]);
  assign and_505_nl = (fsm_output[7]) & (fsm_output[3]) & mux_2367_nl;
  assign mux_2371_nl = MUX_s_1_2_2(mux_2370_nl, and_505_nl, fsm_output[4]);
  assign or_2539_nl = (~ (fsm_output[6])) | (~ (fsm_output[0])) | (fsm_output[9])
      | (~ (fsm_output[2])) | (fsm_output[8]) | (~ (fsm_output[5]));
  assign mux_2364_nl = MUX_s_1_2_2(mux_2374_cse, or_2549_cse, fsm_output[6]);
  assign mux_2365_nl = MUX_s_1_2_2(or_2539_nl, mux_2364_nl, fsm_output[3]);
  assign nor_537_nl = ~((fsm_output[7]) | mux_2365_nl);
  assign or_2531_nl = (fsm_output[9]) | (fsm_output[2]) | (~ (fsm_output[8])) | (fsm_output[5]);
  assign or_2530_nl = (~ (fsm_output[9])) | (fsm_output[2]) | (~ (fsm_output[8]))
      | (fsm_output[5]);
  assign mux_2361_nl = MUX_s_1_2_2(or_2531_nl, or_2530_nl, fsm_output[0]);
  assign nor_538_nl = ~((fsm_output[3]) | (fsm_output[6]) | mux_2361_nl);
  assign nor_539_nl = ~((~ (fsm_output[6])) | (fsm_output[0]) | (fsm_output[9]) |
      nand_169_cse);
  assign nor_540_nl = ~((~ (fsm_output[6])) | (fsm_output[0]) | (~ (fsm_output[9]))
      | (fsm_output[2]) | (fsm_output[8]) | (fsm_output[5]));
  assign mux_2360_nl = MUX_s_1_2_2(nor_539_nl, nor_540_nl, fsm_output[3]);
  assign mux_2362_nl = MUX_s_1_2_2(nor_538_nl, mux_2360_nl, fsm_output[7]);
  assign mux_2366_nl = MUX_s_1_2_2(nor_537_nl, mux_2362_nl, fsm_output[4]);
  assign COMP_LOOP_10_modExp_dev_1_while_mul_mut_mx0c4 = MUX_s_1_2_2(mux_2371_nl,
      mux_2366_nl, fsm_output[1]);
  assign or_2571_nl = (~ (fsm_output[5])) | (~ (fsm_output[8])) | (fsm_output[2]);
  assign or_2625_nl = (fsm_output[8]) | (~ (fsm_output[2])) | (fsm_output[5]);
  assign mux_2382_nl = MUX_s_1_2_2(or_2571_nl, or_2625_nl, fsm_output[9]);
  assign nand_172_nl = ~((fsm_output[9]) & (fsm_output[5]) & (fsm_output[8]) & (~
      (fsm_output[2])));
  assign mux_2383_nl = MUX_s_1_2_2(mux_2382_nl, nand_172_nl, fsm_output[0]);
  assign nor_525_nl = ~((fsm_output[4]) | (fsm_output[1]) | mux_2383_nl);
  assign nor_526_nl = ~((~ (fsm_output[0])) | (fsm_output[9]) | (~ (fsm_output[5]))
      | (fsm_output[8]) | (~ (fsm_output[2])));
  assign nor_527_nl = ~((fsm_output[0]) | (~ (fsm_output[9])) | (~ (fsm_output[5]))
      | (fsm_output[8]) | (~ (fsm_output[2])));
  assign mux_2381_nl = MUX_s_1_2_2(nor_526_nl, nor_527_nl, fsm_output[1]);
  assign and_501_nl = (fsm_output[4]) & mux_2381_nl;
  assign mux_2384_nl = MUX_s_1_2_2(nor_525_nl, and_501_nl, fsm_output[6]);
  assign nor_528_nl = ~((~ (fsm_output[4])) | (fsm_output[1]) | mux_2374_cse);
  assign or_2560_nl = (fsm_output[0]) | (~ (fsm_output[9])) | (fsm_output[5]) | (~
      (fsm_output[8])) | (fsm_output[2]);
  assign mux_2379_nl = MUX_s_1_2_2(or_2549_cse, or_2560_nl, fsm_output[1]);
  assign and_502_nl = (fsm_output[4]) & (~ mux_2379_nl);
  assign mux_2380_nl = MUX_s_1_2_2(nor_528_nl, and_502_nl, fsm_output[6]);
  assign mux_2385_nl = MUX_s_1_2_2(mux_2384_nl, mux_2380_nl, fsm_output[3]);
  assign nor_529_nl = ~((fsm_output[9]) | (fsm_output[5]) | (~ (fsm_output[8])) |
      (fsm_output[2]));
  assign nor_530_nl = ~((~ (fsm_output[9])) | (fsm_output[5]) | (~ (fsm_output[8]))
      | (fsm_output[2]));
  assign mux_2376_nl = MUX_s_1_2_2(nor_529_nl, nor_530_nl, fsm_output[0]);
  assign and_503_nl = (fsm_output[4]) & (fsm_output[1]) & mux_2376_nl;
  assign mux_2377_nl = MUX_s_1_2_2(and_503_nl, nor_558_cse, fsm_output[6]);
  assign nor_532_nl = ~((fsm_output[4]) | (~ (fsm_output[1])) | mux_2374_cse);
  assign or_2550_nl = (fsm_output[0]) | (~ (fsm_output[9])) | (~ (fsm_output[5]))
      | (fsm_output[8]) | (fsm_output[2]);
  assign mux_2373_nl = MUX_s_1_2_2(or_2550_nl, or_2549_cse, fsm_output[1]);
  assign nor_533_nl = ~((fsm_output[4]) | mux_2373_nl);
  assign mux_2375_nl = MUX_s_1_2_2(nor_532_nl, nor_533_nl, fsm_output[6]);
  assign mux_2378_nl = MUX_s_1_2_2(mux_2377_nl, mux_2375_nl, fsm_output[3]);
  assign COMP_LOOP_10_modExp_dev_1_while_mul_mut_mx0c5 = MUX_s_1_2_2(mux_2385_nl,
      mux_2378_nl, fsm_output[7]);
  assign STAGE_VEC_LOOP_j_sva_9_0_mx0c1 = and_dcpl_268 & and_dcpl_266 & nor_tmp_130;
  assign COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c3 =
      and_dcpl_253 & and_dcpl_243;
  assign COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c4 =
      and_dcpl_257 & and_dcpl_106;
  assign COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c5 =
      and_dcpl_109 & and_dcpl_256;
  assign COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c6 =
      and_dcpl_97 & and_dcpl_260;
  assign COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c7 =
      and_dcpl_244 & and_dcpl_263;
  assign COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c8 =
      and_dcpl_253 & and_dcpl_270;
  assign COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c9 =
      and_dcpl_311 & and_dcpl_319;
  assign COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c10 =
      and_dcpl_261 & and_dcpl_321;
  assign COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c11 =
      and_dcpl_268 & and_dcpl_279;
  assign COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c12 =
      and_dcpl_109 & and_dcpl_284;
  assign COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c13 =
      and_dcpl_239 & and_dcpl_286;
  assign or_2664_nl = (fsm_output[5]) | (~ nor_tmp_399);
  assign mux_2541_nl = MUX_s_1_2_2(nand_tmp_140, or_2664_nl, fsm_output[4]);
  assign mux_2542_nl = MUX_s_1_2_2(mux_tmp_2474, mux_2541_nl, fsm_output[0]);
  assign mux_2539_nl = MUX_s_1_2_2(or_tmp_2588, or_tmp_2587, fsm_output[4]);
  assign mux_2540_nl = MUX_s_1_2_2(mux_tmp_2470, mux_2539_nl, fsm_output[0]);
  assign mux_2543_nl = MUX_s_1_2_2(mux_2542_nl, mux_2540_nl, fsm_output[7]);
  assign mux_2535_nl = MUX_s_1_2_2((~ or_tmp_2549), nor_tmp_403, fsm_output[5]);
  assign mux_2536_nl = MUX_s_1_2_2((~ or_tmp_2585), mux_2535_nl, fsm_output[4]);
  assign mux_2537_nl = MUX_s_1_2_2(mux_tmp_2461, mux_2536_nl, fsm_output[0]);
  assign mux_2532_nl = MUX_s_1_2_2(or_tmp_2439, (~ nor_tmp_399), fsm_output[5]);
  assign mux_2533_nl = MUX_s_1_2_2(mux_2532_nl, nand_tmp_140, fsm_output[4]);
  assign nand_139_nl = ~((fsm_output[5]) & (~ mux_tmp_2400));
  assign mux_2530_nl = MUX_s_1_2_2((~ mux_tmp_2462), nand_139_nl, fsm_output[4]);
  assign mux_2534_nl = MUX_s_1_2_2(mux_2533_nl, mux_2530_nl, fsm_output[0]);
  assign mux_2538_nl = MUX_s_1_2_2((~ mux_2537_nl), mux_2534_nl, fsm_output[7]);
  assign mux_2544_nl = MUX_s_1_2_2(mux_2543_nl, mux_2538_nl, fsm_output[8]);
  assign nand_138_nl = ~((fsm_output[5]) & (~ mux_tmp_2468));
  assign mux_2526_nl = MUX_s_1_2_2(nand_138_nl, or_tmp_2588, fsm_output[4]);
  assign mux_2527_nl = MUX_s_1_2_2(mux_2526_nl, mux_tmp_2474, fsm_output[0]);
  assign mux_2522_nl = MUX_s_1_2_2(mux_tmp_2469, or_tmp_2585, fsm_output[4]);
  assign mux_2523_nl = MUX_s_1_2_2(mux_2522_nl, mux_tmp_2470, fsm_output[0]);
  assign mux_2528_nl = MUX_s_1_2_2(mux_2527_nl, mux_2523_nl, fsm_output[7]);
  assign mux_2514_nl = MUX_s_1_2_2(and_dcpl_95, mux_tmp_2458, and_516_cse);
  assign nor_520_nl = ~((fsm_output[5]) | mux_2514_nl);
  assign mux_2515_nl = MUX_s_1_2_2(nor_520_nl, mux_tmp_2462, fsm_output[4]);
  assign mux_2516_nl = MUX_s_1_2_2(mux_2515_nl, mux_tmp_2461, fsm_output[0]);
  assign mux_2517_nl = MUX_s_1_2_2((~ mux_2516_nl), or_tmp_2548, fsm_output[7]);
  assign mux_2529_nl = MUX_s_1_2_2(mux_2528_nl, mux_2517_nl, fsm_output[8]);
  assign mux_2545_itm = MUX_s_1_2_2(mux_2544_nl, mux_2529_nl, fsm_output[9]);
  assign operator_64_false_slc_operator_64_false_acc_1_60_itm_mx0c1 = and_dcpl_261
      & and_dcpl_307;
  assign operator_64_false_slc_operator_64_false_acc_1_60_itm_mx0c2 = and_dcpl_239
      & and_dcpl_267;
  assign operator_64_false_slc_operator_64_false_acc_1_60_itm_mx0c3 = and_dcpl_257
      & and_dcpl_323;
  assign operator_64_false_slc_operator_64_false_acc_1_60_itm_mx0c4 = and_dcpl_244
      & and_dcpl_288;
  assign tmp_1_lpi_4_dfm_mx0c0 = and_dcpl_97 & and_dcpl_346;
  assign and_332_m1c = and_dcpl_244 & and_dcpl_106;
  assign and_334_m1c = and_dcpl_239 & and_dcpl_307;
  assign and_335_m1c = and_dcpl_253 & and_dcpl_256;
  assign and_338_m1c = and_dcpl_311 & and_dcpl_252;
  assign and_340_m1c = and_dcpl_261 & and_dcpl_313;
  assign and_342_m1c = and_dcpl_257 & and_dcpl_242 & and_dcpl_44;
  assign and_344_m1c = and_dcpl_268 & and_dcpl_317;
  assign and_346_m1c = and_dcpl_109 & and_dcpl_319;
  assign and_348_m1c = and_dcpl_239 & and_dcpl_321;
  assign and_350_m1c = and_dcpl_244 & and_dcpl_323;
  assign and_351_m1c = and_dcpl_248 & and_dcpl_279;
  assign and_352_m1c = and_dcpl_253 & and_dcpl_284;
  assign and_354_m1c = and_dcpl_257 & and_dcpl_255 & and_dcpl_70;
  assign and_356_m1c = and_dcpl_261 & and_dcpl_329;
  assign and_358_m1c = and_dcpl_264 & and_dcpl_331;
  assign or_508_nl = (~ (fsm_output[5])) | (fsm_output[1]);
  assign mux_1051_nl = MUX_s_1_2_2(or_508_nl, or_tmp_546, fsm_output[4]);
  assign and_125_nl = (~ mux_1051_nl) & and_dcpl_95 & (~ (fsm_output[2])) & (fsm_output[0])
      & (~ (fsm_output[7])) & and_dcpl;
  assign and_132_nl = and_dcpl_109 & and_dcpl_106;
  assign and_136_nl = and_dcpl_113 & and_dcpl_94 & (~ (fsm_output[7])) & and_dcpl;
  assign nor_811_nl = ~((fsm_output[1:0]!=2'b00) | (~ nor_tmp_1));
  assign nor_812_nl = ~((~ (fsm_output[0])) | (~ (fsm_output[1])) | (fsm_output[2])
      | (fsm_output[6]) | (fsm_output[3]));
  assign mux_1052_nl = MUX_s_1_2_2(nor_811_nl, nor_812_nl, fsm_output[7]);
  assign and_139_nl = mux_1052_nl & (fsm_output[5:4]==2'b00) & and_dcpl;
  assign and_144_nl = not_tmp_280 & (~ (fsm_output[3])) & (~ (fsm_output[6])) & (~
      (fsm_output[5])) & (fsm_output[7]) & and_dcpl;
  assign and_556_nl = (fsm_output[5:3]==3'b111);
  assign nor_808_nl = ~((fsm_output[5:3]!=3'b000));
  assign mux_1054_nl = MUX_s_1_2_2(and_556_nl, nor_808_nl, fsm_output[0]);
  assign and_149_nl = mux_1054_nl & (~ (fsm_output[6])) & and_dcpl_125;
  assign nor_806_nl = ~((fsm_output[6:4]!=3'b100));
  assign nor_807_nl = ~((fsm_output[6:4]!=3'b011));
  assign mux_1055_nl = MUX_s_1_2_2(nor_806_nl, nor_807_nl, fsm_output[0]);
  assign and_151_nl = mux_1055_nl & (fsm_output[3]) & and_dcpl_125;
  assign nor_804_nl = ~((~ (fsm_output[1])) | (fsm_output[6]) | (~ (fsm_output[3])));
  assign nor_805_nl = ~((fsm_output[1]) | (~ (fsm_output[6])) | (fsm_output[3]));
  assign mux_1056_nl = MUX_s_1_2_2(nor_804_nl, nor_805_nl, fsm_output[0]);
  assign and_156_nl = mux_1056_nl & (fsm_output[2]) & and_dcpl_131 & and_dcpl;
  assign nor_802_nl = ~((~ (fsm_output[7])) | (fsm_output[0]) | (~((fsm_output[4])
      & (fsm_output[5]) & (fsm_output[1]) & (fsm_output[6]))));
  assign nor_803_nl = ~((fsm_output[7]) | (~ (fsm_output[0])) | (fsm_output[4]) |
      (fsm_output[5]) | (fsm_output[1]) | (fsm_output[6]));
  assign mux_1057_nl = MUX_s_1_2_2(nor_802_nl, nor_803_nl, fsm_output[8]);
  assign and_159_nl = mux_1057_nl & and_dcpl_135 & (~ (fsm_output[9]));
  assign and_555_nl = (fsm_output[7]) & (fsm_output[0]) & (fsm_output[4]) & (fsm_output[6])
      & (~ (fsm_output[3]));
  assign nor_801_nl = ~((fsm_output[7]) | (fsm_output[0]) | (fsm_output[4]) | (fsm_output[6])
      | (~ (fsm_output[3])));
  assign mux_1058_nl = MUX_s_1_2_2(and_555_nl, nor_801_nl, fsm_output[8]);
  assign and_163_nl = mux_1058_nl & and_516_cse & (fsm_output[5]) & (~ (fsm_output[9]));
  assign and_171_nl = and_dcpl_147 & xor_dcpl & and_dcpl_143 & (~ (fsm_output[7]))
      & and_dcpl_44;
  assign nor_799_nl = ~((~ (fsm_output[4])) | (fsm_output[1]) | (fsm_output[2]) |
      (fsm_output[6]));
  assign nor_800_nl = ~((fsm_output[4]) | (~((fsm_output[1]) & (fsm_output[2]) &
      (fsm_output[6]))));
  assign mux_1059_nl = MUX_s_1_2_2(nor_799_nl, nor_800_nl, fsm_output[0]);
  assign and_175_nl = mux_1059_nl & (~ (fsm_output[3])) & (fsm_output[5]) & (~ (fsm_output[7]))
      & and_dcpl_44;
  assign nor_798_nl = ~((fsm_output[4:1]!=4'b0100));
  assign and_554_nl = (fsm_output[4:1]==4'b1011);
  assign mux_1060_nl = MUX_s_1_2_2(nor_798_nl, and_554_nl, fsm_output[0]);
  assign and_179_nl = mux_1060_nl & and_613_cse & (~ (fsm_output[7])) & and_dcpl_44;
  assign and_184_nl = not_tmp_292 & (~ (fsm_output[2])) & and_dcpl_159 & and_dcpl_44;
  assign and_188_nl = and_dcpl_96 & xor_dcpl & and_dcpl_158 & (fsm_output[7]) & and_dcpl_44;
  assign nor_795_nl = ~((fsm_output[4]) | (~ (fsm_output[5])) | (~ (fsm_output[1]))
      | (fsm_output[6]) | (fsm_output[3]));
  assign nor_796_nl = ~((~ (fsm_output[4])) | (fsm_output[5]) | (fsm_output[1]) |
      (~ and_711_cse));
  assign mux_1062_nl = MUX_s_1_2_2(nor_795_nl, nor_796_nl, fsm_output[0]);
  assign and_191_nl = mux_1062_nl & (~ (fsm_output[2])) & (fsm_output[7]) & and_dcpl_44;
  assign nor_793_nl = ~((~ (fsm_output[4])) | (fsm_output[5]) | (~ (fsm_output[1])));
  assign nor_794_nl = ~((fsm_output[4]) | (~ (fsm_output[5])) | (fsm_output[1]));
  assign mux_1063_nl = MUX_s_1_2_2(nor_793_nl, nor_794_nl, fsm_output[0]);
  assign and_196_nl = mux_1063_nl & (fsm_output[3]) & (fsm_output[6]) & (~ (fsm_output[2]))
      & (fsm_output[7]) & and_dcpl_44;
  assign and_552_nl = (fsm_output[8]) & (fsm_output[7]) & (fsm_output[0]) & (fsm_output[6])
      & (fsm_output[3]);
  assign nor_792_nl = ~((fsm_output[8]) | (fsm_output[7]) | (fsm_output[0]) | (fsm_output[6])
      | (fsm_output[3]));
  assign mux_1064_nl = MUX_s_1_2_2(and_552_nl, nor_792_nl, fsm_output[9]);
  assign and_200_nl = mux_1064_nl & and_dcpl_176 & (fsm_output[5:4]==2'b01);
  assign nor_790_nl = ~((fsm_output[5:4]!=2'b10));
  assign nor_791_nl = ~((fsm_output[5:4]!=2'b01));
  assign mux_1065_nl = MUX_s_1_2_2(nor_790_nl, nor_791_nl, fsm_output[0]);
  assign and_205_nl = mux_1065_nl & and_dcpl_95 & and_dcpl_176 & (~ (fsm_output[7]))
      & and_dcpl_70;
  assign nor_788_nl = ~((~ (fsm_output[4])) | (fsm_output[1]) | (~ (fsm_output[2]))
      | (fsm_output[6]) | (fsm_output[3]));
  assign nor_789_nl = ~((fsm_output[4]) | (~ (fsm_output[1])) | (fsm_output[2]) |
      (~ and_711_cse));
  assign mux_1066_nl = MUX_s_1_2_2(nor_788_nl, nor_789_nl, fsm_output[0]);
  assign and_208_nl = mux_1066_nl & (~ (fsm_output[5])) & (~ (fsm_output[7])) & and_dcpl_70;
  assign and_213_nl = not_tmp_280 & (fsm_output[3]) & (fsm_output[6]) & (~ (fsm_output[5]))
      & (~ (fsm_output[7])) & and_dcpl_70;
  assign and_218_nl = not_tmp_292 & (fsm_output[2]) & and_dcpl_192 & (~ (fsm_output[4]))
      & and_dcpl_70;
  assign and_223_nl = and_dcpl_199 & xor_dcpl & and_dcpl_192 & (fsm_output[7]) &
      and_dcpl_70;
  assign nor_786_nl = ~((fsm_output[4]) | (fsm_output[5]) | (~ (fsm_output[1])) |
      (fsm_output[3]));
  assign and_762_nl = (fsm_output[4]) & (fsm_output[5]) & (~ (fsm_output[1])) & (fsm_output[3]);
  assign mux_1067_nl = MUX_s_1_2_2(nor_786_nl, and_762_nl, fsm_output[0]);
  assign and_227_nl = mux_1067_nl & (~ (fsm_output[6])) & (fsm_output[2]) & (fsm_output[7])
      & and_dcpl_70;
  assign and_551_nl = (fsm_output[4]) & (fsm_output[5]) & (fsm_output[1]) & (~ (fsm_output[6]));
  assign nor_785_nl = ~((fsm_output[4]) | (fsm_output[5]) | (fsm_output[1]) | (~
      (fsm_output[6])));
  assign mux_1068_nl = MUX_s_1_2_2(and_551_nl, nor_785_nl, fsm_output[0]);
  assign and_231_nl = mux_1068_nl & (fsm_output[3]) & (fsm_output[2]) & (fsm_output[7])
      & and_dcpl_70;
  assign mux_1069_nl = MUX_s_1_2_2(or_tmp_33, or_tmp_591, fsm_output[0]);
  assign and_234_nl = (~ mux_1069_nl) & and_516_cse & and_dcpl_131 & and_dcpl_70;
  assign and_550_nl = (fsm_output[7]) & (fsm_output[0]) & (fsm_output[4]) & (fsm_output[5])
      & (fsm_output[6]);
  assign nor_784_nl = ~((fsm_output[7]) | (fsm_output[0]) | (fsm_output[4]) | (fsm_output[5])
      | (fsm_output[6]));
  assign mux_1070_nl = MUX_s_1_2_2(and_550_nl, nor_784_nl, fsm_output[8]);
  assign and_237_nl = mux_1070_nl & and_dcpl_135 & (fsm_output[1]) & (fsm_output[9]);
  assign nor_782_nl = ~((~ (fsm_output[7])) | (fsm_output[0]) | (~ (fsm_output[4]))
      | (fsm_output[1]) | (fsm_output[2]) | (~ (fsm_output[6])));
  assign nor_783_nl = ~((fsm_output[7]) | (~ (fsm_output[0])) | (fsm_output[4]) |
      (~ (fsm_output[1])) | (~ (fsm_output[2])) | (fsm_output[6]));
  assign mux_1071_nl = MUX_s_1_2_2(nor_782_nl, nor_783_nl, fsm_output[8]);
  assign and_240_nl = mux_1071_nl & (fsm_output[3]) & (fsm_output[5]) & (fsm_output[9]);
  assign nor_781_nl = ~((fsm_output[3:1]!=3'b000));
  assign and_549_nl = (fsm_output[3:1]==3'b111);
  assign mux_1072_nl = MUX_s_1_2_2(nor_781_nl, and_549_nl, fsm_output[0]);
  assign and_245_nl = mux_1072_nl & (~ (fsm_output[6])) & and_623_cse & (~ (fsm_output[7]))
      & nor_tmp_130;
  assign nor_779_nl = ~((fsm_output[4]) | (~ and_711_cse));
  assign nor_780_nl = ~((~ (fsm_output[4])) | (fsm_output[6]) | (fsm_output[3]));
  assign mux_1073_nl = MUX_s_1_2_2(nor_779_nl, nor_780_nl, fsm_output[0]);
  assign and_249_nl = mux_1073_nl & (~ (fsm_output[2])) & and_dcpl_225;
  assign and_250_nl = and_dcpl_113 & and_dcpl_225;
  assign nor_777_nl = ~((fsm_output[0]) | (~((fsm_output[1]) & (fsm_output[6]) &
      (fsm_output[3]))));
  assign nor_778_nl = ~((~ (fsm_output[0])) | (fsm_output[1]) | (fsm_output[6]) |
      (fsm_output[3]));
  assign mux_1074_nl = MUX_s_1_2_2(nor_777_nl, nor_778_nl, fsm_output[7]);
  assign and_254_nl = mux_1074_nl & (~ (fsm_output[2])) & (fsm_output[5]) & (~ (fsm_output[4]))
      & nor_tmp_130;
  assign vec_rsc_0_0_i_adra_d_pff = MUX1HOT_v_6_33_2((COMP_LOOP_1_operator_64_false_acc_tmp[9:4]),
      COMP_LOOP_acc_psp_sva, (operator_64_false_acc_cse_1_sva[9:4]), (COMP_LOOP_acc_cse_2_sva[9:4]),
      (operator_64_false_acc_cse_2_sva[9:4]), (COMP_LOOP_acc_7_psp_sva[8:3]), (operator_64_false_acc_cse_3_sva[9:4]),
      (COMP_LOOP_acc_cse_4_sva[9:4]), (operator_64_false_acc_cse_4_sva[9:4]), (COMP_LOOP_acc_8_psp_sva[7:2]),
      (operator_64_false_acc_cse_5_sva[9:4]), (COMP_LOOP_acc_cse_6_sva[9:4]), (operator_64_false_acc_cse_6_sva[9:4]),
      (COMP_LOOP_acc_9_psp_sva[8:3]), (operator_64_false_acc_cse_7_sva[9:4]), (COMP_LOOP_acc_cse_8_sva[9:4]),
      (operator_64_false_acc_cse_8_sva[9:4]), (COMP_LOOP_acc_10_psp_sva[6:1]), (operator_64_false_acc_cse_9_sva[9:4]),
      (COMP_LOOP_acc_cse_10_sva[9:4]), (operator_64_false_acc_cse_10_sva[9:4]), (COMP_LOOP_acc_11_psp_sva[8:3]),
      (operator_64_false_acc_cse_11_sva[9:4]), (COMP_LOOP_acc_cse_12_sva[9:4]), (operator_64_false_acc_cse_12_sva[9:4]),
      (COMP_LOOP_acc_12_psp_sva[7:2]), (operator_64_false_acc_cse_13_sva[9:4]), (COMP_LOOP_acc_cse_14_sva[9:4]),
      (operator_64_false_acc_cse_14_sva[9:4]), (COMP_LOOP_acc_13_psp_sva[8:3]), (operator_64_false_acc_cse_15_sva[9:4]),
      (COMP_LOOP_acc_cse_sva[9:4]), (operator_64_false_acc_cse_sva[9:4]), {and_dcpl_98
      , and_125_nl , and_132_nl , and_136_nl , and_139_nl , and_144_nl , and_149_nl
      , and_151_nl , and_156_nl , and_159_nl , and_163_nl , and_171_nl , and_175_nl
      , and_179_nl , and_184_nl , and_188_nl , and_191_nl , and_196_nl , and_200_nl
      , and_205_nl , and_208_nl , and_213_nl , and_218_nl , and_223_nl , and_227_nl
      , and_231_nl , and_234_nl , and_237_nl , and_240_nl , and_245_nl , and_249_nl
      , and_250_nl , and_254_nl});
  assign vec_rsc_0_0_i_da_d_pff = COMP_LOOP_1_modulo_dev_cmp_return_rsc_z;
  assign nor_765_nl = ~((operator_64_false_acc_cse_1_sva[3:0]!=4'b0000) | (fsm_output[2])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]));
  assign nor_766_nl = ~((COMP_LOOP_acc_cse_2_sva[3:0]!=4'b0000) | (fsm_output[2])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]));
  assign mux_1103_nl = MUX_s_1_2_2(nor_765_nl, nor_766_nl, fsm_output[4]);
  assign nor_767_nl = ~((operator_64_false_acc_cse_5_sva[3:0]!=4'b0000) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5])));
  assign nor_768_nl = ~((COMP_LOOP_acc_cse_6_sva[3:0]!=4'b0000) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5])));
  assign mux_1102_nl = MUX_s_1_2_2(nor_767_nl, nor_768_nl, fsm_output[4]);
  assign mux_1104_nl = MUX_s_1_2_2(mux_1103_nl, mux_1102_nl, fsm_output[8]);
  assign nand_18_nl = ~((fsm_output[1]) & mux_1104_nl);
  assign nor_769_nl = ~((operator_64_false_acc_cse_15_sva[3:0]!=4'b0000) | (fsm_output[2])
      | not_tmp_311);
  assign nor_770_nl = ~((COMP_LOOP_acc_cse_sva[3:0]!=4'b0000) | (fsm_output[2]) |
      not_tmp_311);
  assign mux_1100_nl = MUX_s_1_2_2(nor_769_nl, nor_770_nl, fsm_output[4]);
  assign nand_17_nl = ~((fsm_output[8]) & mux_1100_nl);
  assign or_711_nl = (COMP_LOOP_acc_cse_10_sva[3:0]!=4'b0000) | (fsm_output[2]) |
      (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign or_709_nl = (operator_64_false_acc_cse_9_sva[3:0]!=4'b0000) | (fsm_output[2])
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1098_nl = MUX_s_1_2_2(or_711_nl, or_709_nl, fsm_output[4]);
  assign or_708_nl = (fsm_output[4]) | (COMP_LOOP_acc_cse_14_sva[3:0]!=4'b0000) |
      (~ (fsm_output[2])) | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1099_nl = MUX_s_1_2_2(mux_1098_nl, or_708_nl, fsm_output[8]);
  assign mux_1101_nl = MUX_s_1_2_2(nand_17_nl, mux_1099_nl, fsm_output[1]);
  assign mux_1105_nl = MUX_s_1_2_2(nand_18_nl, mux_1101_nl, fsm_output[9]);
  assign or_706_nl = (COMP_LOOP_acc_cse_4_sva[3:0]!=4'b0000) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]);
  assign or_705_nl = (operator_64_false_acc_cse_3_sva[3:0]!=4'b0000) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign mux_1095_nl = MUX_s_1_2_2(or_706_nl, or_705_nl, fsm_output[4]);
  assign or_703_nl = (operator_64_false_acc_cse_7_sva[3:0]!=4'b0000) | (fsm_output[2])
      | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign or_701_nl = (COMP_LOOP_acc_cse_8_sva[3:0]!=4'b0000) | (fsm_output[2]) |
      (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign mux_1094_nl = MUX_s_1_2_2(or_703_nl, or_701_nl, fsm_output[4]);
  assign mux_1096_nl = MUX_s_1_2_2(mux_1095_nl, mux_1094_nl, fsm_output[8]);
  assign or_707_nl = (fsm_output[1]) | mux_1096_nl;
  assign or_698_nl = (operator_64_false_acc_cse_11_sva[3:0]!=4'b0000) | (~ (fsm_output[2]))
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign or_697_nl = (COMP_LOOP_acc_cse_12_sva[3:0]!=4'b0000) | (~ (fsm_output[2]))
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1092_nl = MUX_s_1_2_2(or_698_nl, or_697_nl, fsm_output[4]);
  assign or_699_nl = (fsm_output[8]) | mux_1092_nl;
  assign or_696_nl = (operator_64_false_acc_cse_13_sva[3:0]!=4'b0000) | (fsm_output[8])
      | (~ (fsm_output[4])) | (~ (fsm_output[2])) | (fsm_output[3]) | not_tmp_312;
  assign mux_1093_nl = MUX_s_1_2_2(or_699_nl, or_696_nl, fsm_output[1]);
  assign mux_1097_nl = MUX_s_1_2_2(or_707_nl, mux_1093_nl, fsm_output[9]);
  assign mux_1106_nl = MUX_s_1_2_2(mux_1105_nl, mux_1097_nl, fsm_output[7]);
  assign or_692_nl = (COMP_LOOP_acc_8_psp_sva[1:0]!=2'b00) | (fsm_output[4]) | (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b00)
      | (~ (fsm_output[2])) | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1087_nl = MUX_s_1_2_2(or_694_cse, or_692_nl, fsm_output[8]);
  assign mux_1088_nl = MUX_s_1_2_2(mux_1087_nl, nand_tmp_16, fsm_output[1]);
  assign or_691_nl = (~ (fsm_output[8])) | (COMP_LOOP_acc_8_psp_sva[1:0]!=2'b00)
      | (fsm_output[4]) | (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b00) | (~ (fsm_output[2]))
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1086_nl = MUX_s_1_2_2(or_691_nl, nand_tmp_16, fsm_output[1]);
  assign mux_1089_nl = MUX_s_1_2_2(mux_1088_nl, mux_1086_nl, STAGE_VEC_LOOP_j_sva_9_0[3]);
  assign nor_771_nl = ~((operator_64_false_acc_cse_10_sva[3:0]!=4'b0000) | (fsm_output[2])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]));
  assign nor_772_nl = ~((COMP_LOOP_acc_11_psp_sva[2:0]!=3'b000) | (STAGE_VEC_LOOP_j_sva_9_0[0])
      | (fsm_output[2]) | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]));
  assign mux_1083_nl = MUX_s_1_2_2(nor_771_nl, nor_772_nl, fsm_output[4]);
  assign nor_773_nl = ~((operator_64_false_acc_cse_14_sva[3:0]!=4'b0000) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5])));
  assign nor_774_nl = ~((COMP_LOOP_acc_13_psp_sva[2:0]!=3'b000) | (STAGE_VEC_LOOP_j_sva_9_0[0])
      | (~ (fsm_output[2])) | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5])));
  assign mux_1082_nl = MUX_s_1_2_2(nor_773_nl, nor_774_nl, fsm_output[4]);
  assign mux_1084_nl = MUX_s_1_2_2(mux_1083_nl, mux_1082_nl, fsm_output[8]);
  assign nand_15_nl = ~((fsm_output[1]) & mux_1084_nl);
  assign mux_1090_nl = MUX_s_1_2_2(mux_1089_nl, nand_15_nl, fsm_output[9]);
  assign or_680_nl = (operator_64_false_acc_cse_4_sva[3:0]!=4'b0000) | (fsm_output[4:2]!=3'b101)
      | not_tmp_312;
  assign or_678_nl = (STAGE_VEC_LOOP_j_sva_9_0[2:0]!=3'b000) | (COMP_LOOP_acc_10_psp_sva[0])
      | (fsm_output[2]) | not_tmp_311;
  assign or_676_nl = (operator_64_false_acc_cse_8_sva[3:0]!=4'b0000) | (fsm_output[2])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]);
  assign mux_1078_nl = MUX_s_1_2_2(or_678_nl, or_676_nl, fsm_output[4]);
  assign mux_1079_nl = MUX_s_1_2_2(or_680_nl, mux_1078_nl, fsm_output[8]);
  assign or_674_nl = (operator_64_false_acc_cse_2_sva[3:0]!=4'b0000) | (fsm_output[2])
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign or_673_nl = (COMP_LOOP_acc_7_psp_sva[2:0]!=3'b000) | (STAGE_VEC_LOOP_j_sva_9_0[0])
      | (fsm_output[2]) | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1077_nl = MUX_s_1_2_2(or_674_nl, or_673_nl, fsm_output[4]);
  assign or_675_nl = (fsm_output[8]) | mux_1077_nl;
  assign mux_1080_nl = MUX_s_1_2_2(mux_1079_nl, or_675_nl, fsm_output[1]);
  assign or_671_nl = (COMP_LOOP_acc_12_psp_sva[1:0]!=2'b00) | (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b00)
      | (~ (fsm_output[2])) | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]);
  assign or_670_nl = (operator_64_false_acc_cse_12_sva[3:0]!=4'b0000) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign mux_1075_nl = MUX_s_1_2_2(or_671_nl, or_670_nl, fsm_output[4]);
  assign or_668_nl = (fsm_output[4]) | (operator_64_false_acc_cse_sva[3:0]!=4'b0000)
      | (fsm_output[2]) | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign mux_1076_nl = MUX_s_1_2_2(mux_1075_nl, or_668_nl, fsm_output[8]);
  assign or_672_nl = (fsm_output[1]) | mux_1076_nl;
  assign mux_1081_nl = MUX_s_1_2_2(mux_1080_nl, or_672_nl, fsm_output[9]);
  assign mux_1091_nl = MUX_s_1_2_2(mux_1090_nl, mux_1081_nl, fsm_output[7]);
  assign mux_1107_nl = MUX_s_1_2_2(mux_1106_nl, mux_1091_nl, fsm_output[0]);
  assign vec_rsc_0_0_i_wea_d_pff = ~ mux_1107_nl;
  assign or_775_nl = (operator_64_false_acc_cse_2_sva[3:0]!=4'b0000) | (fsm_output[4])
      | (fsm_output[0]) | (fsm_output[5]) | not_tmp_322;
  assign or_773_nl = (COMP_LOOP_acc_cse_2_sva[3:0]!=4'b0000) | (~ (fsm_output[0]))
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[5])
      | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign or_772_nl = (COMP_LOOP_1_operator_64_false_acc_tmp[3:0]!=4'b0000) | (fsm_output[5])
      | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign or_771_nl = (STAGE_VEC_LOOP_j_sva_9_0[3:0]!=4'b0000) | (fsm_output[5]) |
      (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign mux_1137_nl = MUX_s_1_2_2(or_772_nl, or_771_nl, fsm_output[0]);
  assign mux_1138_nl = MUX_s_1_2_2(or_773_nl, mux_1137_nl, fsm_output[4]);
  assign mux_1139_nl = MUX_s_1_2_2(or_775_nl, mux_1138_nl, fsm_output[1]);
  assign or_770_nl = (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b000) | (STAGE_VEC_LOOP_j_sva_9_0[0])
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[5])
      | not_tmp_322;
  assign or_768_nl = (operator_64_false_acc_cse_11_sva[3:0]!=4'b0000) | (fsm_output[5])
      | not_tmp_322;
  assign mux_1134_nl = MUX_s_1_2_2(or_770_nl, or_768_nl, fsm_output[0]);
  assign or_766_nl = (fsm_output[0]) | (operator_64_false_acc_cse_10_sva[3:0]!=4'b0000)
      | (fsm_output[5]) | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign mux_1135_nl = MUX_s_1_2_2(mux_1134_nl, or_766_nl, fsm_output[4]);
  assign or_764_nl = (~ (fsm_output[4])) | (~ (fsm_output[0])) | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      | (COMP_LOOP_acc_cse_10_sva[3:0]!=4'b0000) | (fsm_output[5]) | (fsm_output[6])
      | (fsm_output[3]) | (fsm_output[2]);
  assign mux_1136_nl = MUX_s_1_2_2(mux_1135_nl, or_764_nl, fsm_output[1]);
  assign mux_1140_nl = MUX_s_1_2_2(mux_1139_nl, mux_1136_nl, fsm_output[9]);
  assign or_763_nl = (COMP_LOOP_acc_9_psp_sva[2:0]!=3'b000) | (STAGE_VEC_LOOP_j_sva_9_0[0])
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (~
      (fsm_output[5])) | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign or_762_nl = (operator_64_false_acc_cse_7_sva[3:0]!=4'b0000) | (~ (fsm_output[5]))
      | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign mux_1130_nl = MUX_s_1_2_2(or_763_nl, or_762_nl, fsm_output[0]);
  assign or_761_nl = (operator_64_false_acc_cse_6_sva[3:0]!=4'b0000) | (fsm_output[0])
      | (~ (fsm_output[5])) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign mux_1131_nl = MUX_s_1_2_2(mux_1130_nl, or_761_nl, fsm_output[4]);
  assign or_760_nl = (COMP_LOOP_acc_cse_6_sva[3:0]!=4'b0000) | (fsm_output[4]) |
      (~ (fsm_output[0])) | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      | (fsm_output[6:5]!=2'b01) | nand_442_cse;
  assign mux_1132_nl = MUX_s_1_2_2(mux_1131_nl, or_760_nl, fsm_output[1]);
  assign or_758_nl = (COMP_LOOP_acc_cse_sva[3:0]!=4'b0000) | (~ operator_64_false_slc_operator_64_false_acc_1_60_itm)
      | (~ (fsm_output[0])) | (~ (fsm_output[5])) | (~ (fsm_output[6])) | (~ (fsm_output[3]))
      | (fsm_output[2]);
  assign or_757_nl = (COMP_LOOP_acc_13_psp_sva[2:0]!=3'b000) | (STAGE_VEC_LOOP_j_sva_9_0[0])
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (~
      (fsm_output[5])) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign or_756_nl = (operator_64_false_acc_cse_15_sva[3:0]!=4'b0000) | (~ (fsm_output[5]))
      | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign mux_1127_nl = MUX_s_1_2_2(or_757_nl, or_756_nl, fsm_output[0]);
  assign mux_1128_nl = MUX_s_1_2_2(or_758_nl, mux_1127_nl, fsm_output[4]);
  assign or_755_nl = (operator_64_false_acc_cse_sva[3:0]!=4'b0000) | (fsm_output[4])
      | (fsm_output[0]) | (~ (fsm_output[5])) | (~ (fsm_output[6])) | (~ (fsm_output[3]))
      | (fsm_output[2]);
  assign mux_1129_nl = MUX_s_1_2_2(mux_1128_nl, or_755_nl, fsm_output[1]);
  assign mux_1133_nl = MUX_s_1_2_2(mux_1132_nl, mux_1129_nl, fsm_output[9]);
  assign mux_1141_nl = MUX_s_1_2_2(mux_1140_nl, mux_1133_nl, fsm_output[8]);
  assign or_754_nl = (COMP_LOOP_acc_7_psp_sva[2:0]!=3'b000) | (STAGE_VEC_LOOP_j_sva_9_0[0])
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[5])
      | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign or_752_nl = (operator_64_false_acc_cse_3_sva[3:0]!=4'b0000) | (fsm_output[5])
      | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign mux_1122_nl = MUX_s_1_2_2(or_754_nl, or_752_nl, fsm_output[0]);
  assign or_750_nl = (~ operator_64_false_slc_operator_64_false_acc_1_60_itm) | (COMP_LOOP_acc_cse_4_sva[3:0]!=4'b0000)
      | (~ (fsm_output[0])) | (~ (fsm_output[5])) | (fsm_output[6]) | nand_442_cse;
  assign mux_1123_nl = MUX_s_1_2_2(mux_1122_nl, or_750_nl, fsm_output[4]);
  assign or_748_nl = (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b00) | (COMP_LOOP_acc_8_psp_sva[1:0]!=2'b00)
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm);
  assign mux_1119_nl = MUX_s_1_2_2(nand_tmp_19, or_tmp_669, or_748_nl);
  assign or_747_nl = (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b00) | (COMP_LOOP_acc_8_psp_sva[1:0]!=2'b00)
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (~
      (fsm_output[5])) | (~ (fsm_output[6])) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign or_745_nl = (operator_64_false_acc_cse_4_sva[3:0]!=4'b0000);
  assign mux_1120_nl = MUX_s_1_2_2(mux_1119_nl, or_747_nl, or_745_nl);
  assign or_744_nl = (operator_64_false_acc_cse_5_sva[3:0]!=4'b0000) | (~ (fsm_output[5]))
      | (~ (fsm_output[6])) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign mux_1121_nl = MUX_s_1_2_2(mux_1120_nl, or_744_nl, fsm_output[0]);
  assign nand_20_nl = ~((fsm_output[4]) & (~ mux_1121_nl));
  assign mux_1124_nl = MUX_s_1_2_2(mux_1123_nl, nand_20_nl, fsm_output[1]);
  assign or_742_nl = (COMP_LOOP_acc_cse_12_sva[3:0]!=4'b0000) | (~ operator_64_false_slc_operator_64_false_acc_1_60_itm)
      | (~ (fsm_output[0])) | (fsm_output[5]) | (fsm_output[6]) | (fsm_output[3])
      | (~ (fsm_output[2]));
  assign or_740_nl = (operator_64_false_acc_cse_14_sva[3:0]!=4'b0000) | (fsm_output[0])
      | (~ (fsm_output[5])) | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign mux_1117_nl = MUX_s_1_2_2(or_742_nl, or_740_nl, fsm_output[4]);
  assign or_739_nl = (operator_64_false_acc_cse_12_sva[3:0]!=4'b0000) | (fsm_output[0])
      | (fsm_output[5]) | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign or_737_nl = (COMP_LOOP_acc_12_psp_sva[1:0]!=2'b00) | (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b00)
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[6:5]!=2'b01)
      | nand_442_cse;
  assign or_730_nl = (operator_64_false_acc_cse_13_sva[3:0]!=4'b0000);
  assign mux_1113_nl = MUX_s_1_2_2(mux_1112_cse, nand_437_cse, or_730_nl);
  assign or_729_nl = (operator_64_false_acc_cse_13_sva[3:0]!=4'b0000) | (fsm_output[6:5]!=2'b01)
      | nand_442_cse;
  assign or_727_nl = (COMP_LOOP_acc_cse_14_sva[3:0]!=4'b0000);
  assign mux_1114_nl = MUX_s_1_2_2(mux_1113_nl, or_729_nl, or_727_nl);
  assign mux_1115_nl = MUX_s_1_2_2(or_737_nl, mux_1114_nl, fsm_output[0]);
  assign mux_1116_nl = MUX_s_1_2_2(or_739_nl, mux_1115_nl, fsm_output[4]);
  assign mux_1118_nl = MUX_s_1_2_2(mux_1117_nl, mux_1116_nl, fsm_output[1]);
  assign mux_1125_nl = MUX_s_1_2_2(mux_1124_nl, mux_1118_nl, fsm_output[9]);
  assign or_725_nl = (COMP_LOOP_acc_cse_8_sva[3:0]!=4'b0000) | (fsm_output[4]) |
      (~ operator_64_false_slc_operator_64_false_acc_1_60_itm) | (~ (fsm_output[0]))
      | (~ (fsm_output[5])) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign or_724_nl = (operator_64_false_acc_cse_8_sva[3:0]!=4'b0000) | (fsm_output[0])
      | (~ (fsm_output[5])) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign or_723_nl = (STAGE_VEC_LOOP_j_sva_9_0[2:0]!=3'b000) | (COMP_LOOP_acc_10_psp_sva[0])
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[5])
      | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign or_722_nl = (operator_64_false_acc_cse_9_sva[3:0]!=4'b0000) | (fsm_output[5])
      | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign mux_1108_nl = MUX_s_1_2_2(or_723_nl, or_722_nl, fsm_output[0]);
  assign mux_1109_nl = MUX_s_1_2_2(or_724_nl, mux_1108_nl, fsm_output[4]);
  assign mux_1110_nl = MUX_s_1_2_2(or_725_nl, mux_1109_nl, fsm_output[1]);
  assign or_726_nl = (fsm_output[9]) | mux_1110_nl;
  assign mux_1126_nl = MUX_s_1_2_2(mux_1125_nl, or_726_nl, fsm_output[8]);
  assign mux_1142_nl = MUX_s_1_2_2(mux_1141_nl, mux_1126_nl, fsm_output[7]);
  assign vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d = ~ mux_1142_nl;
  assign nor_753_nl = ~((operator_64_false_acc_cse_1_sva[3:0]!=4'b0001) | (fsm_output[2])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]));
  assign nor_754_nl = ~((COMP_LOOP_acc_cse_2_sva[3:0]!=4'b0001) | (fsm_output[2])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]));
  assign mux_1171_nl = MUX_s_1_2_2(nor_753_nl, nor_754_nl, fsm_output[4]);
  assign nor_755_nl = ~((operator_64_false_acc_cse_5_sva[3:0]!=4'b0001) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5])));
  assign nor_756_nl = ~((COMP_LOOP_acc_cse_6_sva[3:0]!=4'b0001) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5])));
  assign mux_1170_nl = MUX_s_1_2_2(nor_755_nl, nor_756_nl, fsm_output[4]);
  assign mux_1172_nl = MUX_s_1_2_2(mux_1171_nl, mux_1170_nl, fsm_output[8]);
  assign nand_24_nl = ~((fsm_output[1]) & mux_1172_nl);
  assign nor_757_nl = ~((operator_64_false_acc_cse_15_sva[3:0]!=4'b0001) | (fsm_output[2])
      | not_tmp_311);
  assign nor_758_nl = ~((COMP_LOOP_acc_cse_sva[3:0]!=4'b0001) | (fsm_output[2]) |
      not_tmp_311);
  assign mux_1168_nl = MUX_s_1_2_2(nor_757_nl, nor_758_nl, fsm_output[4]);
  assign nand_23_nl = ~((fsm_output[8]) & mux_1168_nl);
  assign or_820_nl = (COMP_LOOP_acc_cse_10_sva[3:0]!=4'b0001) | (fsm_output[2]) |
      (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign or_818_nl = (operator_64_false_acc_cse_9_sva[3:0]!=4'b0001) | (fsm_output[2])
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1166_nl = MUX_s_1_2_2(or_820_nl, or_818_nl, fsm_output[4]);
  assign or_817_nl = (fsm_output[4]) | (COMP_LOOP_acc_cse_14_sva[3:0]!=4'b0001) |
      (~ (fsm_output[2])) | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1167_nl = MUX_s_1_2_2(mux_1166_nl, or_817_nl, fsm_output[8]);
  assign mux_1169_nl = MUX_s_1_2_2(nand_23_nl, mux_1167_nl, fsm_output[1]);
  assign mux_1173_nl = MUX_s_1_2_2(nand_24_nl, mux_1169_nl, fsm_output[9]);
  assign or_815_nl = (COMP_LOOP_acc_cse_4_sva[3:0]!=4'b0001) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]);
  assign or_814_nl = (operator_64_false_acc_cse_3_sva[3:0]!=4'b0001) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign mux_1163_nl = MUX_s_1_2_2(or_815_nl, or_814_nl, fsm_output[4]);
  assign or_812_nl = (operator_64_false_acc_cse_7_sva[3:0]!=4'b0001) | (fsm_output[2])
      | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign or_810_nl = (COMP_LOOP_acc_cse_8_sva[3:0]!=4'b0001) | (fsm_output[2]) |
      (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign mux_1162_nl = MUX_s_1_2_2(or_812_nl, or_810_nl, fsm_output[4]);
  assign mux_1164_nl = MUX_s_1_2_2(mux_1163_nl, mux_1162_nl, fsm_output[8]);
  assign or_816_nl = (fsm_output[1]) | mux_1164_nl;
  assign or_807_nl = (operator_64_false_acc_cse_11_sva[3:0]!=4'b0001) | (~ (fsm_output[2]))
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign or_806_nl = (COMP_LOOP_acc_cse_12_sva[3:0]!=4'b0001) | (~ (fsm_output[2]))
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1160_nl = MUX_s_1_2_2(or_807_nl, or_806_nl, fsm_output[4]);
  assign or_808_nl = (fsm_output[8]) | mux_1160_nl;
  assign or_805_nl = (operator_64_false_acc_cse_13_sva[3:0]!=4'b0001) | (fsm_output[8])
      | (~ (fsm_output[4])) | (~ (fsm_output[2])) | (fsm_output[3]) | not_tmp_312;
  assign mux_1161_nl = MUX_s_1_2_2(or_808_nl, or_805_nl, fsm_output[1]);
  assign mux_1165_nl = MUX_s_1_2_2(or_816_nl, mux_1161_nl, fsm_output[9]);
  assign mux_1174_nl = MUX_s_1_2_2(mux_1173_nl, mux_1165_nl, fsm_output[7]);
  assign or_801_nl = (COMP_LOOP_acc_8_psp_sva[1:0]!=2'b00) | (fsm_output[4]) | (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b01)
      | (~ (fsm_output[2])) | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1155_nl = MUX_s_1_2_2(or_803_cse, or_801_nl, fsm_output[8]);
  assign mux_1156_nl = MUX_s_1_2_2(mux_1155_nl, nand_tmp_22, fsm_output[1]);
  assign or_800_nl = (~ (fsm_output[8])) | (COMP_LOOP_acc_8_psp_sva[1:0]!=2'b00)
      | (fsm_output[4]) | (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b01) | (~ (fsm_output[2]))
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1154_nl = MUX_s_1_2_2(or_800_nl, nand_tmp_22, fsm_output[1]);
  assign mux_1157_nl = MUX_s_1_2_2(mux_1156_nl, mux_1154_nl, STAGE_VEC_LOOP_j_sva_9_0[3]);
  assign nor_759_nl = ~((operator_64_false_acc_cse_10_sva[3:0]!=4'b0001) | (fsm_output[2])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]));
  assign nor_760_nl = ~((COMP_LOOP_acc_11_psp_sva[2:0]!=3'b000) | (~ (STAGE_VEC_LOOP_j_sva_9_0[0]))
      | (fsm_output[2]) | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]));
  assign mux_1151_nl = MUX_s_1_2_2(nor_759_nl, nor_760_nl, fsm_output[4]);
  assign nor_761_nl = ~((operator_64_false_acc_cse_14_sva[3:0]!=4'b0001) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5])));
  assign nor_762_nl = ~((COMP_LOOP_acc_13_psp_sva[2:0]!=3'b000) | (~ (STAGE_VEC_LOOP_j_sva_9_0[0]))
      | (~ (fsm_output[2])) | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5])));
  assign mux_1150_nl = MUX_s_1_2_2(nor_761_nl, nor_762_nl, fsm_output[4]);
  assign mux_1152_nl = MUX_s_1_2_2(mux_1151_nl, mux_1150_nl, fsm_output[8]);
  assign nand_21_nl = ~((fsm_output[1]) & mux_1152_nl);
  assign mux_1158_nl = MUX_s_1_2_2(mux_1157_nl, nand_21_nl, fsm_output[9]);
  assign or_789_nl = (operator_64_false_acc_cse_4_sva[3:0]!=4'b0001) | (fsm_output[4:2]!=3'b101)
      | not_tmp_312;
  assign or_787_nl = (STAGE_VEC_LOOP_j_sva_9_0[2:0]!=3'b001) | (COMP_LOOP_acc_10_psp_sva[0])
      | (fsm_output[2]) | not_tmp_311;
  assign or_785_nl = (operator_64_false_acc_cse_8_sva[3:0]!=4'b0001) | (fsm_output[2])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]);
  assign mux_1146_nl = MUX_s_1_2_2(or_787_nl, or_785_nl, fsm_output[4]);
  assign mux_1147_nl = MUX_s_1_2_2(or_789_nl, mux_1146_nl, fsm_output[8]);
  assign or_783_nl = (operator_64_false_acc_cse_2_sva[3:0]!=4'b0001) | (fsm_output[2])
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign or_782_nl = (COMP_LOOP_acc_7_psp_sva[2:0]!=3'b000) | (~ (STAGE_VEC_LOOP_j_sva_9_0[0]))
      | (fsm_output[2]) | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1145_nl = MUX_s_1_2_2(or_783_nl, or_782_nl, fsm_output[4]);
  assign or_784_nl = (fsm_output[8]) | mux_1145_nl;
  assign mux_1148_nl = MUX_s_1_2_2(mux_1147_nl, or_784_nl, fsm_output[1]);
  assign or_780_nl = (COMP_LOOP_acc_12_psp_sva[1:0]!=2'b00) | (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b01)
      | (~ (fsm_output[2])) | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]);
  assign or_779_nl = (operator_64_false_acc_cse_12_sva[3:0]!=4'b0001) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign mux_1143_nl = MUX_s_1_2_2(or_780_nl, or_779_nl, fsm_output[4]);
  assign or_777_nl = (fsm_output[4]) | (operator_64_false_acc_cse_sva[3:0]!=4'b0001)
      | (fsm_output[2]) | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign mux_1144_nl = MUX_s_1_2_2(mux_1143_nl, or_777_nl, fsm_output[8]);
  assign or_781_nl = (fsm_output[1]) | mux_1144_nl;
  assign mux_1149_nl = MUX_s_1_2_2(mux_1148_nl, or_781_nl, fsm_output[9]);
  assign mux_1159_nl = MUX_s_1_2_2(mux_1158_nl, mux_1149_nl, fsm_output[7]);
  assign mux_1175_nl = MUX_s_1_2_2(mux_1174_nl, mux_1159_nl, fsm_output[0]);
  assign vec_rsc_0_1_i_wea_d_pff = ~ mux_1175_nl;
  assign or_881_nl = (operator_64_false_acc_cse_2_sva[3:0]!=4'b0001) | (fsm_output[4])
      | (fsm_output[0]) | (fsm_output[5]) | not_tmp_322;
  assign or_879_nl = (COMP_LOOP_acc_cse_2_sva[3:0]!=4'b0001) | (~ (fsm_output[0]))
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[5])
      | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign or_878_nl = (COMP_LOOP_1_operator_64_false_acc_tmp[3:0]!=4'b0001) | (fsm_output[5])
      | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign or_877_nl = (STAGE_VEC_LOOP_j_sva_9_0[3:0]!=4'b0001) | (fsm_output[5]) |
      (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign mux_1205_nl = MUX_s_1_2_2(or_878_nl, or_877_nl, fsm_output[0]);
  assign mux_1206_nl = MUX_s_1_2_2(or_879_nl, mux_1205_nl, fsm_output[4]);
  assign mux_1207_nl = MUX_s_1_2_2(or_881_nl, mux_1206_nl, fsm_output[1]);
  assign or_876_nl = (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b000) | (~ (STAGE_VEC_LOOP_j_sva_9_0[0]))
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[5])
      | not_tmp_322;
  assign or_874_nl = (operator_64_false_acc_cse_11_sva[3:0]!=4'b0001) | (fsm_output[5])
      | not_tmp_322;
  assign mux_1202_nl = MUX_s_1_2_2(or_876_nl, or_874_nl, fsm_output[0]);
  assign or_872_nl = (fsm_output[0]) | (operator_64_false_acc_cse_10_sva[3:0]!=4'b0001)
      | (fsm_output[5]) | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign mux_1203_nl = MUX_s_1_2_2(mux_1202_nl, or_872_nl, fsm_output[4]);
  assign or_870_nl = (COMP_LOOP_acc_cse_10_sva[3:0]!=4'b0001) | (~ (fsm_output[4]))
      | (~ (fsm_output[0])) | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      | (fsm_output[5]) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign mux_1204_nl = MUX_s_1_2_2(mux_1203_nl, or_870_nl, fsm_output[1]);
  assign mux_1208_nl = MUX_s_1_2_2(mux_1207_nl, mux_1204_nl, fsm_output[9]);
  assign or_869_nl = (COMP_LOOP_acc_9_psp_sva[2:0]!=3'b000) | (~ (STAGE_VEC_LOOP_j_sva_9_0[0]))
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (~
      (fsm_output[5])) | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign or_868_nl = (operator_64_false_acc_cse_7_sva[3:0]!=4'b0001) | (~ (fsm_output[5]))
      | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign mux_1198_nl = MUX_s_1_2_2(or_869_nl, or_868_nl, fsm_output[0]);
  assign or_867_nl = (operator_64_false_acc_cse_6_sva[3:0]!=4'b0001) | (fsm_output[0])
      | (~ (fsm_output[5])) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign mux_1199_nl = MUX_s_1_2_2(mux_1198_nl, or_867_nl, fsm_output[4]);
  assign or_866_nl = (COMP_LOOP_acc_cse_6_sva[3:0]!=4'b0001) | (fsm_output[4]) |
      (~ (fsm_output[0])) | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      | (fsm_output[6:5]!=2'b01) | nand_442_cse;
  assign mux_1200_nl = MUX_s_1_2_2(mux_1199_nl, or_866_nl, fsm_output[1]);
  assign or_864_nl = (COMP_LOOP_acc_cse_sva[3:0]!=4'b0001) | (~ operator_64_false_slc_operator_64_false_acc_1_60_itm)
      | (~ (fsm_output[0])) | (~ (fsm_output[5])) | (~ (fsm_output[6])) | (~ (fsm_output[3]))
      | (fsm_output[2]);
  assign or_863_nl = (COMP_LOOP_acc_13_psp_sva[2:0]!=3'b000) | (~ (STAGE_VEC_LOOP_j_sva_9_0[0]))
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (~
      (fsm_output[5])) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign or_862_nl = (operator_64_false_acc_cse_15_sva[3:0]!=4'b0001) | (~ (fsm_output[5]))
      | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign mux_1195_nl = MUX_s_1_2_2(or_863_nl, or_862_nl, fsm_output[0]);
  assign mux_1196_nl = MUX_s_1_2_2(or_864_nl, mux_1195_nl, fsm_output[4]);
  assign or_861_nl = (operator_64_false_acc_cse_sva[3:0]!=4'b0001) | (fsm_output[4])
      | (fsm_output[0]) | (~ (fsm_output[5])) | (~ (fsm_output[6])) | (~ (fsm_output[3]))
      | (fsm_output[2]);
  assign mux_1197_nl = MUX_s_1_2_2(mux_1196_nl, or_861_nl, fsm_output[1]);
  assign mux_1201_nl = MUX_s_1_2_2(mux_1200_nl, mux_1197_nl, fsm_output[9]);
  assign mux_1209_nl = MUX_s_1_2_2(mux_1208_nl, mux_1201_nl, fsm_output[8]);
  assign or_860_nl = (COMP_LOOP_acc_7_psp_sva[2:0]!=3'b000) | (~ (STAGE_VEC_LOOP_j_sva_9_0[0]))
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[5])
      | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign or_858_nl = (operator_64_false_acc_cse_3_sva[3:0]!=4'b0001) | (fsm_output[5])
      | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign mux_1190_nl = MUX_s_1_2_2(or_860_nl, or_858_nl, fsm_output[0]);
  assign or_856_nl = (~ operator_64_false_slc_operator_64_false_acc_1_60_itm) | (COMP_LOOP_acc_cse_4_sva[3:0]!=4'b0001)
      | (~ (fsm_output[0])) | (~ (fsm_output[5])) | (fsm_output[6]) | nand_442_cse;
  assign mux_1191_nl = MUX_s_1_2_2(mux_1190_nl, or_856_nl, fsm_output[4]);
  assign or_854_nl = (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b01) | (COMP_LOOP_acc_8_psp_sva[1:0]!=2'b00)
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (~
      (fsm_output[5])) | (~ (fsm_output[6])) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign or_852_nl = (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b01) | (COMP_LOOP_acc_8_psp_sva[1:0]!=2'b00)
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm);
  assign mux_1187_nl = MUX_s_1_2_2(nand_tmp_19, or_tmp_669, or_852_nl);
  assign nor_277_nl = ~((operator_64_false_acc_cse_4_sva[3:0]!=4'b0001));
  assign mux_1188_nl = MUX_s_1_2_2(or_854_nl, mux_1187_nl, nor_277_nl);
  assign or_851_nl = (operator_64_false_acc_cse_5_sva[3:0]!=4'b0001) | (~ (fsm_output[5]))
      | (~ (fsm_output[6])) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign mux_1189_nl = MUX_s_1_2_2(mux_1188_nl, or_851_nl, fsm_output[0]);
  assign nand_26_nl = ~((fsm_output[4]) & (~ mux_1189_nl));
  assign mux_1192_nl = MUX_s_1_2_2(mux_1191_nl, nand_26_nl, fsm_output[1]);
  assign or_849_nl = (COMP_LOOP_acc_cse_12_sva[3:0]!=4'b0001) | (~ operator_64_false_slc_operator_64_false_acc_1_60_itm)
      | (~ (fsm_output[0])) | (fsm_output[5]) | (fsm_output[6]) | (fsm_output[3])
      | (~ (fsm_output[2]));
  assign or_847_nl = (operator_64_false_acc_cse_14_sva[3:0]!=4'b0001) | (fsm_output[0])
      | (~ (fsm_output[5])) | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign mux_1185_nl = MUX_s_1_2_2(or_849_nl, or_847_nl, fsm_output[4]);
  assign or_846_nl = (operator_64_false_acc_cse_12_sva[3:0]!=4'b0001) | (fsm_output[0])
      | (fsm_output[5]) | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign or_844_nl = (COMP_LOOP_acc_12_psp_sva[1:0]!=2'b00) | (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b01)
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[6:5]!=2'b01)
      | nand_442_cse;
  assign or_842_nl = (operator_64_false_acc_cse_13_sva[3:0]!=4'b0001) | (fsm_output[6:5]!=2'b01)
      | nand_442_cse;
  assign nor_275_nl = ~((operator_64_false_acc_cse_13_sva[3:0]!=4'b0001));
  assign mux_1181_nl = MUX_s_1_2_2(nand_437_cse, mux_1112_cse, nor_275_nl);
  assign nor_274_nl = ~((COMP_LOOP_acc_cse_14_sva[3:0]!=4'b0001));
  assign mux_1182_nl = MUX_s_1_2_2(or_842_nl, mux_1181_nl, nor_274_nl);
  assign mux_1183_nl = MUX_s_1_2_2(or_844_nl, mux_1182_nl, fsm_output[0]);
  assign mux_1184_nl = MUX_s_1_2_2(or_846_nl, mux_1183_nl, fsm_output[4]);
  assign mux_1186_nl = MUX_s_1_2_2(mux_1185_nl, mux_1184_nl, fsm_output[1]);
  assign mux_1193_nl = MUX_s_1_2_2(mux_1192_nl, mux_1186_nl, fsm_output[9]);
  assign or_834_nl = (COMP_LOOP_acc_cse_8_sva[3:0]!=4'b0001) | (fsm_output[4]) |
      (~ operator_64_false_slc_operator_64_false_acc_1_60_itm) | (~ (fsm_output[0]))
      | (~ (fsm_output[5])) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign or_833_nl = (operator_64_false_acc_cse_8_sva[3:0]!=4'b0001) | (fsm_output[0])
      | (~ (fsm_output[5])) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign or_832_nl = (STAGE_VEC_LOOP_j_sva_9_0[2:0]!=3'b001) | (COMP_LOOP_acc_10_psp_sva[0])
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[5])
      | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign or_831_nl = (operator_64_false_acc_cse_9_sva[3:0]!=4'b0001) | (fsm_output[5])
      | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign mux_1176_nl = MUX_s_1_2_2(or_832_nl, or_831_nl, fsm_output[0]);
  assign mux_1177_nl = MUX_s_1_2_2(or_833_nl, mux_1176_nl, fsm_output[4]);
  assign mux_1178_nl = MUX_s_1_2_2(or_834_nl, mux_1177_nl, fsm_output[1]);
  assign or_835_nl = (fsm_output[9]) | mux_1178_nl;
  assign mux_1194_nl = MUX_s_1_2_2(mux_1193_nl, or_835_nl, fsm_output[8]);
  assign mux_1210_nl = MUX_s_1_2_2(mux_1209_nl, mux_1194_nl, fsm_output[7]);
  assign vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d = ~ mux_1210_nl;
  assign nor_741_nl = ~((operator_64_false_acc_cse_1_sva[3:0]!=4'b0010) | (fsm_output[2])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]));
  assign nor_742_nl = ~((COMP_LOOP_acc_cse_2_sva[3:0]!=4'b0010) | (fsm_output[2])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]));
  assign mux_1239_nl = MUX_s_1_2_2(nor_741_nl, nor_742_nl, fsm_output[4]);
  assign nor_743_nl = ~((operator_64_false_acc_cse_5_sva[3:0]!=4'b0010) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5])));
  assign nor_744_nl = ~((COMP_LOOP_acc_cse_6_sva[3:0]!=4'b0010) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5])));
  assign mux_1238_nl = MUX_s_1_2_2(nor_743_nl, nor_744_nl, fsm_output[4]);
  assign mux_1240_nl = MUX_s_1_2_2(mux_1239_nl, mux_1238_nl, fsm_output[8]);
  assign nand_30_nl = ~((fsm_output[1]) & mux_1240_nl);
  assign nor_745_nl = ~((operator_64_false_acc_cse_15_sva[3:0]!=4'b0010) | (fsm_output[2])
      | not_tmp_311);
  assign nor_746_nl = ~((COMP_LOOP_acc_cse_sva[3:0]!=4'b0010) | (fsm_output[2]) |
      not_tmp_311);
  assign mux_1236_nl = MUX_s_1_2_2(nor_745_nl, nor_746_nl, fsm_output[4]);
  assign nand_29_nl = ~((fsm_output[8]) & mux_1236_nl);
  assign or_926_nl = (COMP_LOOP_acc_cse_10_sva[3:0]!=4'b0010) | (fsm_output[2]) |
      (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign or_924_nl = (operator_64_false_acc_cse_9_sva[3:0]!=4'b0010) | (fsm_output[2])
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1234_nl = MUX_s_1_2_2(or_926_nl, or_924_nl, fsm_output[4]);
  assign or_923_nl = (fsm_output[4]) | (COMP_LOOP_acc_cse_14_sva[3:0]!=4'b0010) |
      (~ (fsm_output[2])) | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1235_nl = MUX_s_1_2_2(mux_1234_nl, or_923_nl, fsm_output[8]);
  assign mux_1237_nl = MUX_s_1_2_2(nand_29_nl, mux_1235_nl, fsm_output[1]);
  assign mux_1241_nl = MUX_s_1_2_2(nand_30_nl, mux_1237_nl, fsm_output[9]);
  assign or_921_nl = (COMP_LOOP_acc_cse_4_sva[3:0]!=4'b0010) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]);
  assign or_920_nl = (operator_64_false_acc_cse_3_sva[3:0]!=4'b0010) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign mux_1231_nl = MUX_s_1_2_2(or_921_nl, or_920_nl, fsm_output[4]);
  assign or_918_nl = (operator_64_false_acc_cse_7_sva[3:0]!=4'b0010) | (fsm_output[2])
      | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign or_916_nl = (COMP_LOOP_acc_cse_8_sva[3:0]!=4'b0010) | (fsm_output[2]) |
      (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign mux_1230_nl = MUX_s_1_2_2(or_918_nl, or_916_nl, fsm_output[4]);
  assign mux_1232_nl = MUX_s_1_2_2(mux_1231_nl, mux_1230_nl, fsm_output[8]);
  assign or_922_nl = (fsm_output[1]) | mux_1232_nl;
  assign or_913_nl = (operator_64_false_acc_cse_11_sva[3:0]!=4'b0010) | (~ (fsm_output[2]))
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign or_912_nl = (COMP_LOOP_acc_cse_12_sva[3:0]!=4'b0010) | (~ (fsm_output[2]))
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1228_nl = MUX_s_1_2_2(or_913_nl, or_912_nl, fsm_output[4]);
  assign or_914_nl = (fsm_output[8]) | mux_1228_nl;
  assign or_911_nl = (operator_64_false_acc_cse_13_sva[3:0]!=4'b0010) | (fsm_output[8])
      | (~ (fsm_output[4])) | (~ (fsm_output[2])) | (fsm_output[3]) | not_tmp_312;
  assign mux_1229_nl = MUX_s_1_2_2(or_914_nl, or_911_nl, fsm_output[1]);
  assign mux_1233_nl = MUX_s_1_2_2(or_922_nl, mux_1229_nl, fsm_output[9]);
  assign mux_1242_nl = MUX_s_1_2_2(mux_1241_nl, mux_1233_nl, fsm_output[7]);
  assign or_907_nl = (COMP_LOOP_acc_8_psp_sva[1:0]!=2'b00) | (fsm_output[4]) | (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b10)
      | (~ (fsm_output[2])) | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1223_nl = MUX_s_1_2_2(or_909_cse, or_907_nl, fsm_output[8]);
  assign mux_1224_nl = MUX_s_1_2_2(mux_1223_nl, nand_tmp_28, fsm_output[1]);
  assign or_906_nl = (~ (fsm_output[8])) | (COMP_LOOP_acc_8_psp_sva[1:0]!=2'b00)
      | (fsm_output[4]) | (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b10) | (~ (fsm_output[2]))
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1222_nl = MUX_s_1_2_2(or_906_nl, nand_tmp_28, fsm_output[1]);
  assign mux_1225_nl = MUX_s_1_2_2(mux_1224_nl, mux_1222_nl, STAGE_VEC_LOOP_j_sva_9_0[3]);
  assign nor_747_nl = ~((operator_64_false_acc_cse_10_sva[3:0]!=4'b0010) | (fsm_output[2])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]));
  assign nor_748_nl = ~((COMP_LOOP_acc_11_psp_sva[2:0]!=3'b001) | (STAGE_VEC_LOOP_j_sva_9_0[0])
      | (fsm_output[2]) | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]));
  assign mux_1219_nl = MUX_s_1_2_2(nor_747_nl, nor_748_nl, fsm_output[4]);
  assign nor_749_nl = ~((operator_64_false_acc_cse_14_sva[3:0]!=4'b0010) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5])));
  assign nor_750_nl = ~((COMP_LOOP_acc_13_psp_sva[2:0]!=3'b001) | (STAGE_VEC_LOOP_j_sva_9_0[0])
      | (~ (fsm_output[2])) | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5])));
  assign mux_1218_nl = MUX_s_1_2_2(nor_749_nl, nor_750_nl, fsm_output[4]);
  assign mux_1220_nl = MUX_s_1_2_2(mux_1219_nl, mux_1218_nl, fsm_output[8]);
  assign nand_27_nl = ~((fsm_output[1]) & mux_1220_nl);
  assign mux_1226_nl = MUX_s_1_2_2(mux_1225_nl, nand_27_nl, fsm_output[9]);
  assign or_895_nl = (operator_64_false_acc_cse_4_sva[3:0]!=4'b0010) | (fsm_output[4:2]!=3'b101)
      | not_tmp_312;
  assign or_893_nl = (STAGE_VEC_LOOP_j_sva_9_0[2:0]!=3'b010) | (COMP_LOOP_acc_10_psp_sva[0])
      | (fsm_output[2]) | not_tmp_311;
  assign or_891_nl = (operator_64_false_acc_cse_8_sva[3:0]!=4'b0010) | (fsm_output[2])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]);
  assign mux_1214_nl = MUX_s_1_2_2(or_893_nl, or_891_nl, fsm_output[4]);
  assign mux_1215_nl = MUX_s_1_2_2(or_895_nl, mux_1214_nl, fsm_output[8]);
  assign or_889_nl = (operator_64_false_acc_cse_2_sva[3:0]!=4'b0010) | (fsm_output[2])
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign or_888_nl = (COMP_LOOP_acc_7_psp_sva[2:0]!=3'b001) | (STAGE_VEC_LOOP_j_sva_9_0[0])
      | (fsm_output[2]) | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1213_nl = MUX_s_1_2_2(or_889_nl, or_888_nl, fsm_output[4]);
  assign or_890_nl = (fsm_output[8]) | mux_1213_nl;
  assign mux_1216_nl = MUX_s_1_2_2(mux_1215_nl, or_890_nl, fsm_output[1]);
  assign or_886_nl = (COMP_LOOP_acc_12_psp_sva[1:0]!=2'b00) | (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b10)
      | (~ (fsm_output[2])) | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]);
  assign or_885_nl = (operator_64_false_acc_cse_12_sva[3:0]!=4'b0010) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign mux_1211_nl = MUX_s_1_2_2(or_886_nl, or_885_nl, fsm_output[4]);
  assign or_883_nl = (fsm_output[4]) | (operator_64_false_acc_cse_sva[3:0]!=4'b0010)
      | (fsm_output[2]) | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign mux_1212_nl = MUX_s_1_2_2(mux_1211_nl, or_883_nl, fsm_output[8]);
  assign or_887_nl = (fsm_output[1]) | mux_1212_nl;
  assign mux_1217_nl = MUX_s_1_2_2(mux_1216_nl, or_887_nl, fsm_output[9]);
  assign mux_1227_nl = MUX_s_1_2_2(mux_1226_nl, mux_1217_nl, fsm_output[7]);
  assign mux_1243_nl = MUX_s_1_2_2(mux_1242_nl, mux_1227_nl, fsm_output[0]);
  assign vec_rsc_0_2_i_wea_d_pff = ~ mux_1243_nl;
  assign or_990_nl = (operator_64_false_acc_cse_2_sva[3:0]!=4'b0010) | (fsm_output[4])
      | (fsm_output[0]) | (fsm_output[5]) | not_tmp_322;
  assign or_988_nl = (COMP_LOOP_acc_cse_2_sva[3:0]!=4'b0010) | (~ (fsm_output[0]))
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[5])
      | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign or_987_nl = (COMP_LOOP_1_operator_64_false_acc_tmp[3:0]!=4'b0010) | (fsm_output[5])
      | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign or_986_nl = (STAGE_VEC_LOOP_j_sva_9_0[3:0]!=4'b0010) | (fsm_output[5]) |
      (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign mux_1273_nl = MUX_s_1_2_2(or_987_nl, or_986_nl, fsm_output[0]);
  assign mux_1274_nl = MUX_s_1_2_2(or_988_nl, mux_1273_nl, fsm_output[4]);
  assign mux_1275_nl = MUX_s_1_2_2(or_990_nl, mux_1274_nl, fsm_output[1]);
  assign or_985_nl = (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b001) | (STAGE_VEC_LOOP_j_sva_9_0[0])
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[5])
      | not_tmp_322;
  assign or_983_nl = (operator_64_false_acc_cse_11_sva[3:0]!=4'b0010) | (fsm_output[5])
      | not_tmp_322;
  assign mux_1270_nl = MUX_s_1_2_2(or_985_nl, or_983_nl, fsm_output[0]);
  assign or_981_nl = (fsm_output[0]) | (operator_64_false_acc_cse_10_sva[3:0]!=4'b0010)
      | (fsm_output[5]) | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign mux_1271_nl = MUX_s_1_2_2(mux_1270_nl, or_981_nl, fsm_output[4]);
  assign or_979_nl = (~ (fsm_output[4])) | (~ (fsm_output[0])) | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      | (COMP_LOOP_acc_cse_10_sva[3:0]!=4'b0010) | (fsm_output[5]) | (fsm_output[6])
      | (fsm_output[3]) | (fsm_output[2]);
  assign mux_1272_nl = MUX_s_1_2_2(mux_1271_nl, or_979_nl, fsm_output[1]);
  assign mux_1276_nl = MUX_s_1_2_2(mux_1275_nl, mux_1272_nl, fsm_output[9]);
  assign or_978_nl = (COMP_LOOP_acc_9_psp_sva[2:0]!=3'b001) | (STAGE_VEC_LOOP_j_sva_9_0[0])
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (~
      (fsm_output[5])) | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign or_977_nl = (operator_64_false_acc_cse_7_sva[3:0]!=4'b0010) | (~ (fsm_output[5]))
      | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign mux_1266_nl = MUX_s_1_2_2(or_978_nl, or_977_nl, fsm_output[0]);
  assign or_976_nl = (operator_64_false_acc_cse_6_sva[3:0]!=4'b0010) | (fsm_output[0])
      | (~ (fsm_output[5])) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign mux_1267_nl = MUX_s_1_2_2(mux_1266_nl, or_976_nl, fsm_output[4]);
  assign or_975_nl = (COMP_LOOP_acc_cse_6_sva[3:0]!=4'b0010) | (fsm_output[4]) |
      (~ (fsm_output[0])) | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      | (fsm_output[6:5]!=2'b01) | nand_442_cse;
  assign mux_1268_nl = MUX_s_1_2_2(mux_1267_nl, or_975_nl, fsm_output[1]);
  assign or_973_nl = (~ operator_64_false_slc_operator_64_false_acc_1_60_itm) | (~
      (fsm_output[0])) | (COMP_LOOP_acc_cse_sva[3:0]!=4'b0010) | (~ (fsm_output[5]))
      | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign or_972_nl = (COMP_LOOP_acc_13_psp_sva[2:0]!=3'b001) | (STAGE_VEC_LOOP_j_sva_9_0[0])
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (~
      (fsm_output[5])) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign or_971_nl = (operator_64_false_acc_cse_15_sva[3:0]!=4'b0010) | (~ (fsm_output[5]))
      | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign mux_1263_nl = MUX_s_1_2_2(or_972_nl, or_971_nl, fsm_output[0]);
  assign mux_1264_nl = MUX_s_1_2_2(or_973_nl, mux_1263_nl, fsm_output[4]);
  assign or_970_nl = (operator_64_false_acc_cse_sva[3:0]!=4'b0010) | (fsm_output[4])
      | (fsm_output[0]) | (~ (fsm_output[5])) | (~ (fsm_output[6])) | (~ (fsm_output[3]))
      | (fsm_output[2]);
  assign mux_1265_nl = MUX_s_1_2_2(mux_1264_nl, or_970_nl, fsm_output[1]);
  assign mux_1269_nl = MUX_s_1_2_2(mux_1268_nl, mux_1265_nl, fsm_output[9]);
  assign mux_1277_nl = MUX_s_1_2_2(mux_1276_nl, mux_1269_nl, fsm_output[8]);
  assign or_969_nl = (COMP_LOOP_acc_7_psp_sva[2:0]!=3'b001) | (STAGE_VEC_LOOP_j_sva_9_0[0])
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[5])
      | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign or_967_nl = (operator_64_false_acc_cse_3_sva[3:0]!=4'b0010) | (fsm_output[5])
      | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign mux_1258_nl = MUX_s_1_2_2(or_969_nl, or_967_nl, fsm_output[0]);
  assign or_965_nl = (~ operator_64_false_slc_operator_64_false_acc_1_60_itm) | (COMP_LOOP_acc_cse_4_sva[3:0]!=4'b0010)
      | (~ (fsm_output[0])) | (~ (fsm_output[5])) | (fsm_output[6]) | nand_442_cse;
  assign mux_1259_nl = MUX_s_1_2_2(mux_1258_nl, or_965_nl, fsm_output[4]);
  assign or_963_nl = (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b10) | (COMP_LOOP_acc_8_psp_sva[1:0]!=2'b00)
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm);
  assign mux_1255_nl = MUX_s_1_2_2(nand_tmp_19, or_tmp_669, or_963_nl);
  assign or_962_nl = (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b10) | (COMP_LOOP_acc_8_psp_sva[1:0]!=2'b00)
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (~
      (fsm_output[5])) | (~ (fsm_output[6])) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign or_960_nl = (operator_64_false_acc_cse_4_sva[3:0]!=4'b0010);
  assign mux_1256_nl = MUX_s_1_2_2(mux_1255_nl, or_962_nl, or_960_nl);
  assign or_959_nl = (operator_64_false_acc_cse_5_sva[3:0]!=4'b0010) | (~ (fsm_output[5]))
      | (~ (fsm_output[6])) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign mux_1257_nl = MUX_s_1_2_2(mux_1256_nl, or_959_nl, fsm_output[0]);
  assign nand_32_nl = ~((fsm_output[4]) & (~ mux_1257_nl));
  assign mux_1260_nl = MUX_s_1_2_2(mux_1259_nl, nand_32_nl, fsm_output[1]);
  assign or_957_nl = (~ operator_64_false_slc_operator_64_false_acc_1_60_itm) | (~
      (fsm_output[0])) | (COMP_LOOP_acc_cse_12_sva[3:0]!=4'b0010) | (fsm_output[5])
      | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign or_955_nl = (operator_64_false_acc_cse_14_sva[3:0]!=4'b0010) | (fsm_output[0])
      | (~ (fsm_output[5])) | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign mux_1253_nl = MUX_s_1_2_2(or_957_nl, or_955_nl, fsm_output[4]);
  assign or_954_nl = (operator_64_false_acc_cse_12_sva[3:0]!=4'b0010) | (fsm_output[0])
      | (fsm_output[5]) | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign or_952_nl = (COMP_LOOP_acc_12_psp_sva[1:0]!=2'b00) | (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b10)
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[6:5]!=2'b01)
      | nand_442_cse;
  assign or_945_nl = (operator_64_false_acc_cse_13_sva[3:0]!=4'b0010);
  assign mux_1249_nl = MUX_s_1_2_2(mux_1112_cse, nand_437_cse, or_945_nl);
  assign or_944_nl = (operator_64_false_acc_cse_13_sva[3:0]!=4'b0010) | (fsm_output[6:5]!=2'b01)
      | nand_442_cse;
  assign or_942_nl = (COMP_LOOP_acc_cse_14_sva[3:0]!=4'b0010);
  assign mux_1250_nl = MUX_s_1_2_2(mux_1249_nl, or_944_nl, or_942_nl);
  assign mux_1251_nl = MUX_s_1_2_2(or_952_nl, mux_1250_nl, fsm_output[0]);
  assign mux_1252_nl = MUX_s_1_2_2(or_954_nl, mux_1251_nl, fsm_output[4]);
  assign mux_1254_nl = MUX_s_1_2_2(mux_1253_nl, mux_1252_nl, fsm_output[1]);
  assign mux_1261_nl = MUX_s_1_2_2(mux_1260_nl, mux_1254_nl, fsm_output[9]);
  assign or_940_nl = (COMP_LOOP_acc_cse_8_sva[3:0]!=4'b0010) | (fsm_output[4]) |
      (~ operator_64_false_slc_operator_64_false_acc_1_60_itm) | (~ (fsm_output[0]))
      | (~ (fsm_output[5])) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign or_939_nl = (operator_64_false_acc_cse_8_sva[3:0]!=4'b0010) | (fsm_output[0])
      | (~ (fsm_output[5])) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign or_938_nl = (STAGE_VEC_LOOP_j_sva_9_0[2:0]!=3'b010) | (COMP_LOOP_acc_10_psp_sva[0])
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[5])
      | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign or_937_nl = (operator_64_false_acc_cse_9_sva[3:0]!=4'b0010) | (fsm_output[5])
      | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign mux_1244_nl = MUX_s_1_2_2(or_938_nl, or_937_nl, fsm_output[0]);
  assign mux_1245_nl = MUX_s_1_2_2(or_939_nl, mux_1244_nl, fsm_output[4]);
  assign mux_1246_nl = MUX_s_1_2_2(or_940_nl, mux_1245_nl, fsm_output[1]);
  assign or_941_nl = (fsm_output[9]) | mux_1246_nl;
  assign mux_1262_nl = MUX_s_1_2_2(mux_1261_nl, or_941_nl, fsm_output[8]);
  assign mux_1278_nl = MUX_s_1_2_2(mux_1277_nl, mux_1262_nl, fsm_output[7]);
  assign vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d = ~ mux_1278_nl;
  assign nor_729_nl = ~((operator_64_false_acc_cse_1_sva[3:0]!=4'b0011) | (fsm_output[2])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]));
  assign nor_730_nl = ~((COMP_LOOP_acc_cse_2_sva[3:0]!=4'b0011) | (fsm_output[2])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]));
  assign mux_1307_nl = MUX_s_1_2_2(nor_729_nl, nor_730_nl, fsm_output[4]);
  assign nor_731_nl = ~((operator_64_false_acc_cse_5_sva[3:0]!=4'b0011) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5])));
  assign nor_732_nl = ~((COMP_LOOP_acc_cse_6_sva[3:0]!=4'b0011) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5])));
  assign mux_1306_nl = MUX_s_1_2_2(nor_731_nl, nor_732_nl, fsm_output[4]);
  assign mux_1308_nl = MUX_s_1_2_2(mux_1307_nl, mux_1306_nl, fsm_output[8]);
  assign nand_36_nl = ~((fsm_output[1]) & mux_1308_nl);
  assign nor_733_nl = ~((operator_64_false_acc_cse_15_sva[3:0]!=4'b0011) | (fsm_output[2])
      | not_tmp_311);
  assign nor_734_nl = ~((COMP_LOOP_acc_cse_sva[3:0]!=4'b0011) | (fsm_output[2]) |
      not_tmp_311);
  assign mux_1304_nl = MUX_s_1_2_2(nor_733_nl, nor_734_nl, fsm_output[4]);
  assign nand_35_nl = ~((fsm_output[8]) & mux_1304_nl);
  assign or_1035_nl = (COMP_LOOP_acc_cse_10_sva[3:0]!=4'b0011) | (fsm_output[2])
      | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign or_1033_nl = (operator_64_false_acc_cse_9_sva[3:0]!=4'b0011) | (fsm_output[2])
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1302_nl = MUX_s_1_2_2(or_1035_nl, or_1033_nl, fsm_output[4]);
  assign or_1032_nl = (fsm_output[4]) | (COMP_LOOP_acc_cse_14_sva[3:0]!=4'b0011)
      | (~ (fsm_output[2])) | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1303_nl = MUX_s_1_2_2(mux_1302_nl, or_1032_nl, fsm_output[8]);
  assign mux_1305_nl = MUX_s_1_2_2(nand_35_nl, mux_1303_nl, fsm_output[1]);
  assign mux_1309_nl = MUX_s_1_2_2(nand_36_nl, mux_1305_nl, fsm_output[9]);
  assign or_1030_nl = (COMP_LOOP_acc_cse_4_sva[3:0]!=4'b0011) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]);
  assign or_1029_nl = (operator_64_false_acc_cse_3_sva[3:0]!=4'b0011) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign mux_1299_nl = MUX_s_1_2_2(or_1030_nl, or_1029_nl, fsm_output[4]);
  assign or_1027_nl = (operator_64_false_acc_cse_7_sva[3:0]!=4'b0011) | (fsm_output[2])
      | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign or_1025_nl = (COMP_LOOP_acc_cse_8_sva[3:0]!=4'b0011) | (fsm_output[2]) |
      (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign mux_1298_nl = MUX_s_1_2_2(or_1027_nl, or_1025_nl, fsm_output[4]);
  assign mux_1300_nl = MUX_s_1_2_2(mux_1299_nl, mux_1298_nl, fsm_output[8]);
  assign or_1031_nl = (fsm_output[1]) | mux_1300_nl;
  assign or_1022_nl = (operator_64_false_acc_cse_11_sva[3:0]!=4'b0011) | (~ (fsm_output[2]))
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign or_1021_nl = (COMP_LOOP_acc_cse_12_sva[3:0]!=4'b0011) | (~ (fsm_output[2]))
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1296_nl = MUX_s_1_2_2(or_1022_nl, or_1021_nl, fsm_output[4]);
  assign or_1023_nl = (fsm_output[8]) | mux_1296_nl;
  assign or_1020_nl = (operator_64_false_acc_cse_13_sva[3:0]!=4'b0011) | (fsm_output[8])
      | (~ (fsm_output[4])) | (~ (fsm_output[2])) | (fsm_output[3]) | not_tmp_312;
  assign mux_1297_nl = MUX_s_1_2_2(or_1023_nl, or_1020_nl, fsm_output[1]);
  assign mux_1301_nl = MUX_s_1_2_2(or_1031_nl, mux_1297_nl, fsm_output[9]);
  assign mux_1310_nl = MUX_s_1_2_2(mux_1309_nl, mux_1301_nl, fsm_output[7]);
  assign or_1016_nl = (COMP_LOOP_acc_8_psp_sva[1:0]!=2'b00) | (fsm_output[4]) | (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b11)
      | (~ (fsm_output[2])) | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1291_nl = MUX_s_1_2_2(or_1018_cse, or_1016_nl, fsm_output[8]);
  assign mux_1292_nl = MUX_s_1_2_2(mux_1291_nl, nand_tmp_34, fsm_output[1]);
  assign or_1015_nl = (~ (fsm_output[8])) | (COMP_LOOP_acc_8_psp_sva[1:0]!=2'b00)
      | (fsm_output[4]) | (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b11) | (~ (fsm_output[2]))
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1290_nl = MUX_s_1_2_2(or_1015_nl, nand_tmp_34, fsm_output[1]);
  assign mux_1293_nl = MUX_s_1_2_2(mux_1292_nl, mux_1290_nl, STAGE_VEC_LOOP_j_sva_9_0[3]);
  assign nor_735_nl = ~((operator_64_false_acc_cse_10_sva[3:0]!=4'b0011) | (fsm_output[2])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]));
  assign nor_736_nl = ~((COMP_LOOP_acc_11_psp_sva[2:0]!=3'b001) | (~ (STAGE_VEC_LOOP_j_sva_9_0[0]))
      | (fsm_output[2]) | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]));
  assign mux_1287_nl = MUX_s_1_2_2(nor_735_nl, nor_736_nl, fsm_output[4]);
  assign nor_737_nl = ~((operator_64_false_acc_cse_14_sva[3:0]!=4'b0011) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5])));
  assign nor_738_nl = ~((COMP_LOOP_acc_13_psp_sva[2:0]!=3'b001) | (~ (STAGE_VEC_LOOP_j_sva_9_0[0]))
      | (~ (fsm_output[2])) | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5])));
  assign mux_1286_nl = MUX_s_1_2_2(nor_737_nl, nor_738_nl, fsm_output[4]);
  assign mux_1288_nl = MUX_s_1_2_2(mux_1287_nl, mux_1286_nl, fsm_output[8]);
  assign nand_33_nl = ~((fsm_output[1]) & mux_1288_nl);
  assign mux_1294_nl = MUX_s_1_2_2(mux_1293_nl, nand_33_nl, fsm_output[9]);
  assign or_1004_nl = (operator_64_false_acc_cse_4_sva[3:0]!=4'b0011) | (fsm_output[4:2]!=3'b101)
      | not_tmp_312;
  assign or_1002_nl = (STAGE_VEC_LOOP_j_sva_9_0[2:0]!=3'b011) | (COMP_LOOP_acc_10_psp_sva[0])
      | (fsm_output[2]) | not_tmp_311;
  assign or_1000_nl = (operator_64_false_acc_cse_8_sva[3:0]!=4'b0011) | (fsm_output[2])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]);
  assign mux_1282_nl = MUX_s_1_2_2(or_1002_nl, or_1000_nl, fsm_output[4]);
  assign mux_1283_nl = MUX_s_1_2_2(or_1004_nl, mux_1282_nl, fsm_output[8]);
  assign or_998_nl = (operator_64_false_acc_cse_2_sva[3:0]!=4'b0011) | (fsm_output[2])
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign or_997_nl = (COMP_LOOP_acc_7_psp_sva[2:0]!=3'b001) | (~ (STAGE_VEC_LOOP_j_sva_9_0[0]))
      | (fsm_output[2]) | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1281_nl = MUX_s_1_2_2(or_998_nl, or_997_nl, fsm_output[4]);
  assign or_999_nl = (fsm_output[8]) | mux_1281_nl;
  assign mux_1284_nl = MUX_s_1_2_2(mux_1283_nl, or_999_nl, fsm_output[1]);
  assign or_995_nl = (COMP_LOOP_acc_12_psp_sva[1:0]!=2'b00) | (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b11)
      | (~ (fsm_output[2])) | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]);
  assign or_994_nl = (operator_64_false_acc_cse_12_sva[3:0]!=4'b0011) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign mux_1279_nl = MUX_s_1_2_2(or_995_nl, or_994_nl, fsm_output[4]);
  assign or_992_nl = (fsm_output[4]) | (operator_64_false_acc_cse_sva[3:0]!=4'b0011)
      | (fsm_output[2]) | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign mux_1280_nl = MUX_s_1_2_2(mux_1279_nl, or_992_nl, fsm_output[8]);
  assign or_996_nl = (fsm_output[1]) | mux_1280_nl;
  assign mux_1285_nl = MUX_s_1_2_2(mux_1284_nl, or_996_nl, fsm_output[9]);
  assign mux_1295_nl = MUX_s_1_2_2(mux_1294_nl, mux_1285_nl, fsm_output[7]);
  assign mux_1311_nl = MUX_s_1_2_2(mux_1310_nl, mux_1295_nl, fsm_output[0]);
  assign vec_rsc_0_3_i_wea_d_pff = ~ mux_1311_nl;
  assign or_1096_nl = (operator_64_false_acc_cse_2_sva[3:0]!=4'b0011) | (fsm_output[4])
      | (fsm_output[0]) | (fsm_output[5]) | not_tmp_322;
  assign or_1094_nl = (COMP_LOOP_acc_cse_2_sva[3:0]!=4'b0011) | (~ (fsm_output[0]))
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[5])
      | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign or_1093_nl = (COMP_LOOP_1_operator_64_false_acc_tmp[3:0]!=4'b0011) | (fsm_output[5])
      | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign or_1092_nl = (STAGE_VEC_LOOP_j_sva_9_0[3:0]!=4'b0011) | (fsm_output[5])
      | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign mux_1341_nl = MUX_s_1_2_2(or_1093_nl, or_1092_nl, fsm_output[0]);
  assign mux_1342_nl = MUX_s_1_2_2(or_1094_nl, mux_1341_nl, fsm_output[4]);
  assign mux_1343_nl = MUX_s_1_2_2(or_1096_nl, mux_1342_nl, fsm_output[1]);
  assign or_1091_nl = (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b001) | (~ (STAGE_VEC_LOOP_j_sva_9_0[0]))
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[5])
      | not_tmp_322;
  assign or_1089_nl = (operator_64_false_acc_cse_11_sva[3:0]!=4'b0011) | (fsm_output[5])
      | not_tmp_322;
  assign mux_1338_nl = MUX_s_1_2_2(or_1091_nl, or_1089_nl, fsm_output[0]);
  assign or_1087_nl = (fsm_output[0]) | (operator_64_false_acc_cse_10_sva[3:0]!=4'b0011)
      | (fsm_output[5]) | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign mux_1339_nl = MUX_s_1_2_2(mux_1338_nl, or_1087_nl, fsm_output[4]);
  assign or_1085_nl = (COMP_LOOP_acc_cse_10_sva[3:0]!=4'b0011) | (~ (fsm_output[4]))
      | (~ (fsm_output[0])) | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      | (fsm_output[5]) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign mux_1340_nl = MUX_s_1_2_2(mux_1339_nl, or_1085_nl, fsm_output[1]);
  assign mux_1344_nl = MUX_s_1_2_2(mux_1343_nl, mux_1340_nl, fsm_output[9]);
  assign or_1084_nl = (COMP_LOOP_acc_9_psp_sva[2:0]!=3'b001) | (~ (STAGE_VEC_LOOP_j_sva_9_0[0]))
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (~
      (fsm_output[5])) | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign or_1083_nl = (operator_64_false_acc_cse_7_sva[3:0]!=4'b0011) | (~ (fsm_output[5]))
      | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign mux_1334_nl = MUX_s_1_2_2(or_1084_nl, or_1083_nl, fsm_output[0]);
  assign or_1082_nl = (operator_64_false_acc_cse_6_sva[3:0]!=4'b0011) | (fsm_output[0])
      | (~ (fsm_output[5])) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign mux_1335_nl = MUX_s_1_2_2(mux_1334_nl, or_1082_nl, fsm_output[4]);
  assign or_1081_nl = (COMP_LOOP_acc_cse_6_sva[3:0]!=4'b0011) | (fsm_output[4]) |
      (~ (fsm_output[0])) | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      | (fsm_output[6:5]!=2'b01) | nand_442_cse;
  assign mux_1336_nl = MUX_s_1_2_2(mux_1335_nl, or_1081_nl, fsm_output[1]);
  assign nand_357_nl = ~(operator_64_false_slc_operator_64_false_acc_1_60_itm & (fsm_output[0])
      & (COMP_LOOP_acc_cse_sva[3:0]==4'b0011) & (fsm_output[5]) & (fsm_output[6])
      & (fsm_output[3]) & (~ (fsm_output[2])));
  assign or_1078_nl = (COMP_LOOP_acc_13_psp_sva[2:0]!=3'b001) | (~ (STAGE_VEC_LOOP_j_sva_9_0[0]))
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (~
      (fsm_output[5])) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign or_1077_nl = (operator_64_false_acc_cse_15_sva[3:0]!=4'b0011) | (~ (fsm_output[5]))
      | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign mux_1331_nl = MUX_s_1_2_2(or_1078_nl, or_1077_nl, fsm_output[0]);
  assign mux_1332_nl = MUX_s_1_2_2(nand_357_nl, mux_1331_nl, fsm_output[4]);
  assign or_1076_nl = (operator_64_false_acc_cse_sva[3:0]!=4'b0011) | (fsm_output[4])
      | (fsm_output[0]) | (~ (fsm_output[5])) | (~ (fsm_output[6])) | (~ (fsm_output[3]))
      | (fsm_output[2]);
  assign mux_1333_nl = MUX_s_1_2_2(mux_1332_nl, or_1076_nl, fsm_output[1]);
  assign mux_1337_nl = MUX_s_1_2_2(mux_1336_nl, mux_1333_nl, fsm_output[9]);
  assign mux_1345_nl = MUX_s_1_2_2(mux_1344_nl, mux_1337_nl, fsm_output[8]);
  assign or_1075_nl = (COMP_LOOP_acc_7_psp_sva[2:0]!=3'b001) | (~ (STAGE_VEC_LOOP_j_sva_9_0[0]))
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[5])
      | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign or_1073_nl = (operator_64_false_acc_cse_3_sva[3:0]!=4'b0011) | (fsm_output[5])
      | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign mux_1326_nl = MUX_s_1_2_2(or_1075_nl, or_1073_nl, fsm_output[0]);
  assign or_1071_nl = (~ operator_64_false_slc_operator_64_false_acc_1_60_itm) |
      (COMP_LOOP_acc_cse_4_sva[3:0]!=4'b0011) | (~ (fsm_output[0])) | (~ (fsm_output[5]))
      | (fsm_output[6]) | nand_442_cse;
  assign mux_1327_nl = MUX_s_1_2_2(mux_1326_nl, or_1071_nl, fsm_output[4]);
  assign or_1069_nl = (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b11) | (COMP_LOOP_acc_8_psp_sva[1:0]!=2'b00)
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (~
      (fsm_output[5])) | (~ (fsm_output[6])) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign or_1067_nl = (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b11) | (COMP_LOOP_acc_8_psp_sva[1:0]!=2'b00)
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm);
  assign mux_1323_nl = MUX_s_1_2_2(nand_tmp_19, or_tmp_669, or_1067_nl);
  assign nor_288_nl = ~((operator_64_false_acc_cse_4_sva[3:0]!=4'b0011));
  assign mux_1324_nl = MUX_s_1_2_2(or_1069_nl, mux_1323_nl, nor_288_nl);
  assign or_1066_nl = (operator_64_false_acc_cse_5_sva[3:0]!=4'b0011) | (~ (fsm_output[5]))
      | (~ (fsm_output[6])) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign mux_1325_nl = MUX_s_1_2_2(mux_1324_nl, or_1066_nl, fsm_output[0]);
  assign nand_38_nl = ~((fsm_output[4]) & (~ mux_1325_nl));
  assign mux_1328_nl = MUX_s_1_2_2(mux_1327_nl, nand_38_nl, fsm_output[1]);
  assign or_1064_nl = (~ operator_64_false_slc_operator_64_false_acc_1_60_itm) |
      (~ (fsm_output[0])) | (COMP_LOOP_acc_cse_12_sva[3:0]!=4'b0011) | (fsm_output[5])
      | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign or_1062_nl = (operator_64_false_acc_cse_14_sva[3:0]!=4'b0011) | (fsm_output[0])
      | (~ (fsm_output[5])) | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign mux_1321_nl = MUX_s_1_2_2(or_1064_nl, or_1062_nl, fsm_output[4]);
  assign or_1061_nl = (operator_64_false_acc_cse_12_sva[3:0]!=4'b0011) | (fsm_output[0])
      | (fsm_output[5]) | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign or_1059_nl = (COMP_LOOP_acc_12_psp_sva[1:0]!=2'b00) | (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b11)
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[6:5]!=2'b01)
      | nand_442_cse;
  assign or_1057_nl = (operator_64_false_acc_cse_13_sva[3:0]!=4'b0011) | (fsm_output[6:5]!=2'b01)
      | nand_442_cse;
  assign nor_286_nl = ~((operator_64_false_acc_cse_13_sva[3:0]!=4'b0011));
  assign mux_1317_nl = MUX_s_1_2_2(nand_437_cse, mux_1112_cse, nor_286_nl);
  assign nor_285_nl = ~((COMP_LOOP_acc_cse_14_sva[3:0]!=4'b0011));
  assign mux_1318_nl = MUX_s_1_2_2(or_1057_nl, mux_1317_nl, nor_285_nl);
  assign mux_1319_nl = MUX_s_1_2_2(or_1059_nl, mux_1318_nl, fsm_output[0]);
  assign mux_1320_nl = MUX_s_1_2_2(or_1061_nl, mux_1319_nl, fsm_output[4]);
  assign mux_1322_nl = MUX_s_1_2_2(mux_1321_nl, mux_1320_nl, fsm_output[1]);
  assign mux_1329_nl = MUX_s_1_2_2(mux_1328_nl, mux_1322_nl, fsm_output[9]);
  assign or_1049_nl = (COMP_LOOP_acc_cse_8_sva[3:0]!=4'b0011) | (fsm_output[4]) |
      (~ operator_64_false_slc_operator_64_false_acc_1_60_itm) | (~ (fsm_output[0]))
      | (~ (fsm_output[5])) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign or_1048_nl = (operator_64_false_acc_cse_8_sva[3:0]!=4'b0011) | (fsm_output[0])
      | (~ (fsm_output[5])) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign or_1047_nl = (STAGE_VEC_LOOP_j_sva_9_0[2:0]!=3'b011) | (COMP_LOOP_acc_10_psp_sva[0])
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[5])
      | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign or_1046_nl = (operator_64_false_acc_cse_9_sva[3:0]!=4'b0011) | (fsm_output[5])
      | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign mux_1312_nl = MUX_s_1_2_2(or_1047_nl, or_1046_nl, fsm_output[0]);
  assign mux_1313_nl = MUX_s_1_2_2(or_1048_nl, mux_1312_nl, fsm_output[4]);
  assign mux_1314_nl = MUX_s_1_2_2(or_1049_nl, mux_1313_nl, fsm_output[1]);
  assign or_1050_nl = (fsm_output[9]) | mux_1314_nl;
  assign mux_1330_nl = MUX_s_1_2_2(mux_1329_nl, or_1050_nl, fsm_output[8]);
  assign mux_1346_nl = MUX_s_1_2_2(mux_1345_nl, mux_1330_nl, fsm_output[7]);
  assign vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d = ~ mux_1346_nl;
  assign nor_717_nl = ~((operator_64_false_acc_cse_1_sva[3:0]!=4'b0100) | (fsm_output[2])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]));
  assign nor_718_nl = ~((COMP_LOOP_acc_cse_2_sva[3:0]!=4'b0100) | (fsm_output[2])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]));
  assign mux_1375_nl = MUX_s_1_2_2(nor_717_nl, nor_718_nl, fsm_output[4]);
  assign nor_719_nl = ~((operator_64_false_acc_cse_5_sva[3:0]!=4'b0100) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5])));
  assign nor_720_nl = ~((COMP_LOOP_acc_cse_6_sva[3:0]!=4'b0100) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5])));
  assign mux_1374_nl = MUX_s_1_2_2(nor_719_nl, nor_720_nl, fsm_output[4]);
  assign mux_1376_nl = MUX_s_1_2_2(mux_1375_nl, mux_1374_nl, fsm_output[8]);
  assign nand_42_nl = ~((fsm_output[1]) & mux_1376_nl);
  assign nor_721_nl = ~((operator_64_false_acc_cse_15_sva[3:0]!=4'b0100) | (fsm_output[2])
      | not_tmp_311);
  assign nor_722_nl = ~((COMP_LOOP_acc_cse_sva[3:0]!=4'b0100) | (fsm_output[2]) |
      not_tmp_311);
  assign mux_1372_nl = MUX_s_1_2_2(nor_721_nl, nor_722_nl, fsm_output[4]);
  assign nand_41_nl = ~((fsm_output[8]) & mux_1372_nl);
  assign or_1141_nl = (COMP_LOOP_acc_cse_10_sva[3:0]!=4'b0100) | (fsm_output[2])
      | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign or_1139_nl = (operator_64_false_acc_cse_9_sva[3:0]!=4'b0100) | (fsm_output[2])
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1370_nl = MUX_s_1_2_2(or_1141_nl, or_1139_nl, fsm_output[4]);
  assign or_1138_nl = (fsm_output[4]) | (COMP_LOOP_acc_cse_14_sva[3:0]!=4'b0100)
      | (~ (fsm_output[2])) | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1371_nl = MUX_s_1_2_2(mux_1370_nl, or_1138_nl, fsm_output[8]);
  assign mux_1373_nl = MUX_s_1_2_2(nand_41_nl, mux_1371_nl, fsm_output[1]);
  assign mux_1377_nl = MUX_s_1_2_2(nand_42_nl, mux_1373_nl, fsm_output[9]);
  assign or_1136_nl = (COMP_LOOP_acc_cse_4_sva[3:0]!=4'b0100) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]);
  assign or_1135_nl = (operator_64_false_acc_cse_3_sva[3:0]!=4'b0100) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign mux_1367_nl = MUX_s_1_2_2(or_1136_nl, or_1135_nl, fsm_output[4]);
  assign or_1133_nl = (operator_64_false_acc_cse_7_sva[3:0]!=4'b0100) | (fsm_output[2])
      | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign or_1131_nl = (COMP_LOOP_acc_cse_8_sva[3:0]!=4'b0100) | (fsm_output[2]) |
      (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign mux_1366_nl = MUX_s_1_2_2(or_1133_nl, or_1131_nl, fsm_output[4]);
  assign mux_1368_nl = MUX_s_1_2_2(mux_1367_nl, mux_1366_nl, fsm_output[8]);
  assign or_1137_nl = (fsm_output[1]) | mux_1368_nl;
  assign or_1128_nl = (operator_64_false_acc_cse_11_sva[3:0]!=4'b0100) | (~ (fsm_output[2]))
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign or_1127_nl = (COMP_LOOP_acc_cse_12_sva[3:0]!=4'b0100) | (~ (fsm_output[2]))
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1364_nl = MUX_s_1_2_2(or_1128_nl, or_1127_nl, fsm_output[4]);
  assign or_1129_nl = (fsm_output[8]) | mux_1364_nl;
  assign or_1126_nl = (operator_64_false_acc_cse_13_sva[3:0]!=4'b0100) | (fsm_output[8])
      | (~ (fsm_output[4])) | (~ (fsm_output[2])) | (fsm_output[3]) | not_tmp_312;
  assign mux_1365_nl = MUX_s_1_2_2(or_1129_nl, or_1126_nl, fsm_output[1]);
  assign mux_1369_nl = MUX_s_1_2_2(or_1137_nl, mux_1365_nl, fsm_output[9]);
  assign mux_1378_nl = MUX_s_1_2_2(mux_1377_nl, mux_1369_nl, fsm_output[7]);
  assign or_1122_nl = (COMP_LOOP_acc_8_psp_sva[1:0]!=2'b01) | (fsm_output[4]) | (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b00)
      | (~ (fsm_output[2])) | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1359_nl = MUX_s_1_2_2(or_1124_cse, or_1122_nl, fsm_output[8]);
  assign mux_1360_nl = MUX_s_1_2_2(mux_1359_nl, nand_tmp_40, fsm_output[1]);
  assign or_1121_nl = (~ (fsm_output[8])) | (COMP_LOOP_acc_8_psp_sva[1:0]!=2'b01)
      | (fsm_output[4]) | (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b00) | (~ (fsm_output[2]))
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1358_nl = MUX_s_1_2_2(or_1121_nl, nand_tmp_40, fsm_output[1]);
  assign mux_1361_nl = MUX_s_1_2_2(mux_1360_nl, mux_1358_nl, STAGE_VEC_LOOP_j_sva_9_0[3]);
  assign nor_723_nl = ~((operator_64_false_acc_cse_10_sva[3:0]!=4'b0100) | (fsm_output[2])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]));
  assign nor_724_nl = ~((COMP_LOOP_acc_11_psp_sva[2:0]!=3'b010) | (STAGE_VEC_LOOP_j_sva_9_0[0])
      | (fsm_output[2]) | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]));
  assign mux_1355_nl = MUX_s_1_2_2(nor_723_nl, nor_724_nl, fsm_output[4]);
  assign nor_725_nl = ~((operator_64_false_acc_cse_14_sva[3:0]!=4'b0100) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5])));
  assign nor_726_nl = ~((COMP_LOOP_acc_13_psp_sva[2:0]!=3'b010) | (STAGE_VEC_LOOP_j_sva_9_0[0])
      | (~ (fsm_output[2])) | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5])));
  assign mux_1354_nl = MUX_s_1_2_2(nor_725_nl, nor_726_nl, fsm_output[4]);
  assign mux_1356_nl = MUX_s_1_2_2(mux_1355_nl, mux_1354_nl, fsm_output[8]);
  assign nand_39_nl = ~((fsm_output[1]) & mux_1356_nl);
  assign mux_1362_nl = MUX_s_1_2_2(mux_1361_nl, nand_39_nl, fsm_output[9]);
  assign or_1110_nl = (operator_64_false_acc_cse_4_sva[3:0]!=4'b0100) | (fsm_output[4:2]!=3'b101)
      | not_tmp_312;
  assign or_1108_nl = (STAGE_VEC_LOOP_j_sva_9_0[2:0]!=3'b100) | (COMP_LOOP_acc_10_psp_sva[0])
      | (fsm_output[2]) | not_tmp_311;
  assign or_1106_nl = (operator_64_false_acc_cse_8_sva[3:0]!=4'b0100) | (fsm_output[2])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]);
  assign mux_1350_nl = MUX_s_1_2_2(or_1108_nl, or_1106_nl, fsm_output[4]);
  assign mux_1351_nl = MUX_s_1_2_2(or_1110_nl, mux_1350_nl, fsm_output[8]);
  assign or_1104_nl = (operator_64_false_acc_cse_2_sva[3:0]!=4'b0100) | (fsm_output[2])
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign or_1103_nl = (COMP_LOOP_acc_7_psp_sva[2:0]!=3'b010) | (STAGE_VEC_LOOP_j_sva_9_0[0])
      | (fsm_output[2]) | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1349_nl = MUX_s_1_2_2(or_1104_nl, or_1103_nl, fsm_output[4]);
  assign or_1105_nl = (fsm_output[8]) | mux_1349_nl;
  assign mux_1352_nl = MUX_s_1_2_2(mux_1351_nl, or_1105_nl, fsm_output[1]);
  assign or_1101_nl = (COMP_LOOP_acc_12_psp_sva[1:0]!=2'b01) | (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b00)
      | (~ (fsm_output[2])) | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]);
  assign or_1100_nl = (operator_64_false_acc_cse_12_sva[3:0]!=4'b0100) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign mux_1347_nl = MUX_s_1_2_2(or_1101_nl, or_1100_nl, fsm_output[4]);
  assign or_1098_nl = (fsm_output[4]) | (operator_64_false_acc_cse_sva[3:0]!=4'b0100)
      | (fsm_output[2]) | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign mux_1348_nl = MUX_s_1_2_2(mux_1347_nl, or_1098_nl, fsm_output[8]);
  assign or_1102_nl = (fsm_output[1]) | mux_1348_nl;
  assign mux_1353_nl = MUX_s_1_2_2(mux_1352_nl, or_1102_nl, fsm_output[9]);
  assign mux_1363_nl = MUX_s_1_2_2(mux_1362_nl, mux_1353_nl, fsm_output[7]);
  assign mux_1379_nl = MUX_s_1_2_2(mux_1378_nl, mux_1363_nl, fsm_output[0]);
  assign vec_rsc_0_4_i_wea_d_pff = ~ mux_1379_nl;
  assign or_1205_nl = (operator_64_false_acc_cse_2_sva[3:0]!=4'b0100) | (fsm_output[4])
      | (fsm_output[0]) | (fsm_output[5]) | not_tmp_322;
  assign or_1203_nl = (COMP_LOOP_acc_cse_2_sva[3:0]!=4'b0100) | (~ (fsm_output[0]))
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[5])
      | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign or_1202_nl = (COMP_LOOP_1_operator_64_false_acc_tmp[3:0]!=4'b0100) | (fsm_output[5])
      | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign or_1201_nl = (STAGE_VEC_LOOP_j_sva_9_0[3:0]!=4'b0100) | (fsm_output[5])
      | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign mux_1409_nl = MUX_s_1_2_2(or_1202_nl, or_1201_nl, fsm_output[0]);
  assign mux_1410_nl = MUX_s_1_2_2(or_1203_nl, mux_1409_nl, fsm_output[4]);
  assign mux_1411_nl = MUX_s_1_2_2(or_1205_nl, mux_1410_nl, fsm_output[1]);
  assign or_1200_nl = (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b010) | (STAGE_VEC_LOOP_j_sva_9_0[0])
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[5])
      | not_tmp_322;
  assign or_1198_nl = (operator_64_false_acc_cse_11_sva[3:0]!=4'b0100) | (fsm_output[5])
      | not_tmp_322;
  assign mux_1406_nl = MUX_s_1_2_2(or_1200_nl, or_1198_nl, fsm_output[0]);
  assign or_1196_nl = (fsm_output[0]) | (operator_64_false_acc_cse_10_sva[3:0]!=4'b0100)
      | (fsm_output[5]) | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign mux_1407_nl = MUX_s_1_2_2(mux_1406_nl, or_1196_nl, fsm_output[4]);
  assign or_1194_nl = (~ (fsm_output[4])) | (~ (fsm_output[0])) | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      | (COMP_LOOP_acc_cse_10_sva[3:0]!=4'b0100) | (fsm_output[5]) | (fsm_output[6])
      | (fsm_output[3]) | (fsm_output[2]);
  assign mux_1408_nl = MUX_s_1_2_2(mux_1407_nl, or_1194_nl, fsm_output[1]);
  assign mux_1412_nl = MUX_s_1_2_2(mux_1411_nl, mux_1408_nl, fsm_output[9]);
  assign or_1193_nl = (COMP_LOOP_acc_9_psp_sva[2:0]!=3'b010) | (STAGE_VEC_LOOP_j_sva_9_0[0])
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (~
      (fsm_output[5])) | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign or_1192_nl = (operator_64_false_acc_cse_7_sva[3:0]!=4'b0100) | (~ (fsm_output[5]))
      | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign mux_1402_nl = MUX_s_1_2_2(or_1193_nl, or_1192_nl, fsm_output[0]);
  assign or_1191_nl = (operator_64_false_acc_cse_6_sva[3:0]!=4'b0100) | (fsm_output[0])
      | (~ (fsm_output[5])) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign mux_1403_nl = MUX_s_1_2_2(mux_1402_nl, or_1191_nl, fsm_output[4]);
  assign or_1190_nl = (COMP_LOOP_acc_cse_6_sva[3:0]!=4'b0100) | (fsm_output[4]) |
      (~ (fsm_output[0])) | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      | (fsm_output[6:5]!=2'b01) | nand_442_cse;
  assign mux_1404_nl = MUX_s_1_2_2(mux_1403_nl, or_1190_nl, fsm_output[1]);
  assign or_1188_nl = (COMP_LOOP_acc_cse_sva[3:0]!=4'b0100) | (~ operator_64_false_slc_operator_64_false_acc_1_60_itm)
      | (~ (fsm_output[0])) | (~ (fsm_output[5])) | (~ (fsm_output[6])) | (~ (fsm_output[3]))
      | (fsm_output[2]);
  assign or_1187_nl = (COMP_LOOP_acc_13_psp_sva[2:0]!=3'b010) | (STAGE_VEC_LOOP_j_sva_9_0[0])
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (~
      (fsm_output[5])) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign or_1186_nl = (operator_64_false_acc_cse_15_sva[3:0]!=4'b0100) | (~ (fsm_output[5]))
      | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign mux_1399_nl = MUX_s_1_2_2(or_1187_nl, or_1186_nl, fsm_output[0]);
  assign mux_1400_nl = MUX_s_1_2_2(or_1188_nl, mux_1399_nl, fsm_output[4]);
  assign or_1185_nl = (operator_64_false_acc_cse_sva[3:0]!=4'b0100) | (fsm_output[4])
      | (fsm_output[0]) | (~ (fsm_output[5])) | (~ (fsm_output[6])) | (~ (fsm_output[3]))
      | (fsm_output[2]);
  assign mux_1401_nl = MUX_s_1_2_2(mux_1400_nl, or_1185_nl, fsm_output[1]);
  assign mux_1405_nl = MUX_s_1_2_2(mux_1404_nl, mux_1401_nl, fsm_output[9]);
  assign mux_1413_nl = MUX_s_1_2_2(mux_1412_nl, mux_1405_nl, fsm_output[8]);
  assign or_1184_nl = (COMP_LOOP_acc_7_psp_sva[2:0]!=3'b010) | (STAGE_VEC_LOOP_j_sva_9_0[0])
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[5])
      | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign or_1182_nl = (operator_64_false_acc_cse_3_sva[3:0]!=4'b0100) | (fsm_output[5])
      | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign mux_1394_nl = MUX_s_1_2_2(or_1184_nl, or_1182_nl, fsm_output[0]);
  assign or_1180_nl = (~ operator_64_false_slc_operator_64_false_acc_1_60_itm) |
      (COMP_LOOP_acc_cse_4_sva[3:0]!=4'b0100) | (~ (fsm_output[0])) | (~ (fsm_output[5]))
      | (fsm_output[6]) | nand_442_cse;
  assign mux_1395_nl = MUX_s_1_2_2(mux_1394_nl, or_1180_nl, fsm_output[4]);
  assign or_1178_nl = (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b00) | (COMP_LOOP_acc_8_psp_sva[1:0]!=2'b01)
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm);
  assign mux_1391_nl = MUX_s_1_2_2(nand_tmp_19, or_tmp_669, or_1178_nl);
  assign or_1177_nl = (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b00) | (COMP_LOOP_acc_8_psp_sva[1:0]!=2'b01)
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (~
      (fsm_output[5])) | (~ (fsm_output[6])) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign or_1175_nl = (operator_64_false_acc_cse_4_sva[3:0]!=4'b0100);
  assign mux_1392_nl = MUX_s_1_2_2(mux_1391_nl, or_1177_nl, or_1175_nl);
  assign or_1174_nl = (operator_64_false_acc_cse_5_sva[3:0]!=4'b0100) | (~ (fsm_output[5]))
      | (~ (fsm_output[6])) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign mux_1393_nl = MUX_s_1_2_2(mux_1392_nl, or_1174_nl, fsm_output[0]);
  assign nand_44_nl = ~((fsm_output[4]) & (~ mux_1393_nl));
  assign mux_1396_nl = MUX_s_1_2_2(mux_1395_nl, nand_44_nl, fsm_output[1]);
  assign or_1172_nl = (COMP_LOOP_acc_cse_12_sva[3:0]!=4'b0100) | (~ operator_64_false_slc_operator_64_false_acc_1_60_itm)
      | (~ (fsm_output[0])) | (fsm_output[5]) | (fsm_output[6]) | (fsm_output[3])
      | (~ (fsm_output[2]));
  assign or_1170_nl = (operator_64_false_acc_cse_14_sva[3:0]!=4'b0100) | (fsm_output[0])
      | (~ (fsm_output[5])) | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign mux_1389_nl = MUX_s_1_2_2(or_1172_nl, or_1170_nl, fsm_output[4]);
  assign or_1169_nl = (operator_64_false_acc_cse_12_sva[3:0]!=4'b0100) | (fsm_output[0])
      | (fsm_output[5]) | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign or_1167_nl = (COMP_LOOP_acc_12_psp_sva[1:0]!=2'b01) | (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b00)
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[6:5]!=2'b01)
      | nand_442_cse;
  assign or_1160_nl = (operator_64_false_acc_cse_13_sva[3:0]!=4'b0100);
  assign mux_1385_nl = MUX_s_1_2_2(mux_1112_cse, nand_437_cse, or_1160_nl);
  assign or_1159_nl = (operator_64_false_acc_cse_13_sva[3:0]!=4'b0100) | (fsm_output[6:5]!=2'b01)
      | nand_442_cse;
  assign or_1157_nl = (COMP_LOOP_acc_cse_14_sva[3:0]!=4'b0100);
  assign mux_1386_nl = MUX_s_1_2_2(mux_1385_nl, or_1159_nl, or_1157_nl);
  assign mux_1387_nl = MUX_s_1_2_2(or_1167_nl, mux_1386_nl, fsm_output[0]);
  assign mux_1388_nl = MUX_s_1_2_2(or_1169_nl, mux_1387_nl, fsm_output[4]);
  assign mux_1390_nl = MUX_s_1_2_2(mux_1389_nl, mux_1388_nl, fsm_output[1]);
  assign mux_1397_nl = MUX_s_1_2_2(mux_1396_nl, mux_1390_nl, fsm_output[9]);
  assign or_1155_nl = (COMP_LOOP_acc_cse_8_sva[3:0]!=4'b0100) | (fsm_output[4]) |
      (~ operator_64_false_slc_operator_64_false_acc_1_60_itm) | (~ (fsm_output[0]))
      | (~ (fsm_output[5])) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign or_1154_nl = (operator_64_false_acc_cse_8_sva[3:0]!=4'b0100) | (fsm_output[0])
      | (~ (fsm_output[5])) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign or_1153_nl = (STAGE_VEC_LOOP_j_sva_9_0[2:0]!=3'b100) | (COMP_LOOP_acc_10_psp_sva[0])
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[5])
      | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign or_1152_nl = (operator_64_false_acc_cse_9_sva[3:0]!=4'b0100) | (fsm_output[5])
      | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign mux_1380_nl = MUX_s_1_2_2(or_1153_nl, or_1152_nl, fsm_output[0]);
  assign mux_1381_nl = MUX_s_1_2_2(or_1154_nl, mux_1380_nl, fsm_output[4]);
  assign mux_1382_nl = MUX_s_1_2_2(or_1155_nl, mux_1381_nl, fsm_output[1]);
  assign or_1156_nl = (fsm_output[9]) | mux_1382_nl;
  assign mux_1398_nl = MUX_s_1_2_2(mux_1397_nl, or_1156_nl, fsm_output[8]);
  assign mux_1414_nl = MUX_s_1_2_2(mux_1413_nl, mux_1398_nl, fsm_output[7]);
  assign vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d = ~ mux_1414_nl;
  assign nor_705_nl = ~((operator_64_false_acc_cse_1_sva[3:0]!=4'b0101) | (fsm_output[2])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]));
  assign nor_706_nl = ~((COMP_LOOP_acc_cse_2_sva[3:0]!=4'b0101) | (fsm_output[2])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]));
  assign mux_1443_nl = MUX_s_1_2_2(nor_705_nl, nor_706_nl, fsm_output[4]);
  assign nor_707_nl = ~((operator_64_false_acc_cse_5_sva[3:0]!=4'b0101) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5])));
  assign nor_708_nl = ~((COMP_LOOP_acc_cse_6_sva[3:0]!=4'b0101) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5])));
  assign mux_1442_nl = MUX_s_1_2_2(nor_707_nl, nor_708_nl, fsm_output[4]);
  assign mux_1444_nl = MUX_s_1_2_2(mux_1443_nl, mux_1442_nl, fsm_output[8]);
  assign nand_48_nl = ~((fsm_output[1]) & mux_1444_nl);
  assign nor_709_nl = ~((operator_64_false_acc_cse_15_sva[3:0]!=4'b0101) | (fsm_output[2])
      | not_tmp_311);
  assign nor_710_nl = ~((COMP_LOOP_acc_cse_sva[3:0]!=4'b0101) | (fsm_output[2]) |
      not_tmp_311);
  assign mux_1440_nl = MUX_s_1_2_2(nor_709_nl, nor_710_nl, fsm_output[4]);
  assign nand_47_nl = ~((fsm_output[8]) & mux_1440_nl);
  assign or_1250_nl = (COMP_LOOP_acc_cse_10_sva[3:0]!=4'b0101) | (fsm_output[2])
      | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign or_1248_nl = (operator_64_false_acc_cse_9_sva[3:0]!=4'b0101) | (fsm_output[2])
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1438_nl = MUX_s_1_2_2(or_1250_nl, or_1248_nl, fsm_output[4]);
  assign or_1247_nl = (fsm_output[4]) | (COMP_LOOP_acc_cse_14_sva[3:0]!=4'b0101)
      | (~ (fsm_output[2])) | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1439_nl = MUX_s_1_2_2(mux_1438_nl, or_1247_nl, fsm_output[8]);
  assign mux_1441_nl = MUX_s_1_2_2(nand_47_nl, mux_1439_nl, fsm_output[1]);
  assign mux_1445_nl = MUX_s_1_2_2(nand_48_nl, mux_1441_nl, fsm_output[9]);
  assign or_1245_nl = (COMP_LOOP_acc_cse_4_sva[3:0]!=4'b0101) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]);
  assign or_1244_nl = (operator_64_false_acc_cse_3_sva[3:0]!=4'b0101) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign mux_1435_nl = MUX_s_1_2_2(or_1245_nl, or_1244_nl, fsm_output[4]);
  assign or_1242_nl = (operator_64_false_acc_cse_7_sva[3:0]!=4'b0101) | (fsm_output[2])
      | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign or_1240_nl = (COMP_LOOP_acc_cse_8_sva[3:0]!=4'b0101) | (fsm_output[2]) |
      (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign mux_1434_nl = MUX_s_1_2_2(or_1242_nl, or_1240_nl, fsm_output[4]);
  assign mux_1436_nl = MUX_s_1_2_2(mux_1435_nl, mux_1434_nl, fsm_output[8]);
  assign or_1246_nl = (fsm_output[1]) | mux_1436_nl;
  assign or_1237_nl = (operator_64_false_acc_cse_11_sva[3:0]!=4'b0101) | (~ (fsm_output[2]))
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign or_1236_nl = (COMP_LOOP_acc_cse_12_sva[3:0]!=4'b0101) | (~ (fsm_output[2]))
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1432_nl = MUX_s_1_2_2(or_1237_nl, or_1236_nl, fsm_output[4]);
  assign or_1238_nl = (fsm_output[8]) | mux_1432_nl;
  assign or_1235_nl = (operator_64_false_acc_cse_13_sva[3:0]!=4'b0101) | (fsm_output[8])
      | (~ (fsm_output[4])) | (~ (fsm_output[2])) | (fsm_output[3]) | not_tmp_312;
  assign mux_1433_nl = MUX_s_1_2_2(or_1238_nl, or_1235_nl, fsm_output[1]);
  assign mux_1437_nl = MUX_s_1_2_2(or_1246_nl, mux_1433_nl, fsm_output[9]);
  assign mux_1446_nl = MUX_s_1_2_2(mux_1445_nl, mux_1437_nl, fsm_output[7]);
  assign or_1231_nl = (COMP_LOOP_acc_8_psp_sva[1:0]!=2'b01) | (fsm_output[4]) | (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b01)
      | (~ (fsm_output[2])) | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1427_nl = MUX_s_1_2_2(or_1233_cse, or_1231_nl, fsm_output[8]);
  assign mux_1428_nl = MUX_s_1_2_2(mux_1427_nl, nand_tmp_46, fsm_output[1]);
  assign or_1230_nl = (~ (fsm_output[8])) | (COMP_LOOP_acc_8_psp_sva[1:0]!=2'b01)
      | (fsm_output[4]) | (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b01) | (~ (fsm_output[2]))
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1426_nl = MUX_s_1_2_2(or_1230_nl, nand_tmp_46, fsm_output[1]);
  assign mux_1429_nl = MUX_s_1_2_2(mux_1428_nl, mux_1426_nl, STAGE_VEC_LOOP_j_sva_9_0[3]);
  assign nor_711_nl = ~((operator_64_false_acc_cse_10_sva[3:0]!=4'b0101) | (fsm_output[2])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]));
  assign nor_712_nl = ~((COMP_LOOP_acc_11_psp_sva[2:0]!=3'b010) | (~ (STAGE_VEC_LOOP_j_sva_9_0[0]))
      | (fsm_output[2]) | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]));
  assign mux_1423_nl = MUX_s_1_2_2(nor_711_nl, nor_712_nl, fsm_output[4]);
  assign nor_713_nl = ~((operator_64_false_acc_cse_14_sva[3:0]!=4'b0101) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5])));
  assign nor_714_nl = ~((COMP_LOOP_acc_13_psp_sva[2:0]!=3'b010) | (~ (STAGE_VEC_LOOP_j_sva_9_0[0]))
      | (~ (fsm_output[2])) | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5])));
  assign mux_1422_nl = MUX_s_1_2_2(nor_713_nl, nor_714_nl, fsm_output[4]);
  assign mux_1424_nl = MUX_s_1_2_2(mux_1423_nl, mux_1422_nl, fsm_output[8]);
  assign nand_45_nl = ~((fsm_output[1]) & mux_1424_nl);
  assign mux_1430_nl = MUX_s_1_2_2(mux_1429_nl, nand_45_nl, fsm_output[9]);
  assign or_1219_nl = (operator_64_false_acc_cse_4_sva[3:0]!=4'b0101) | (fsm_output[4:2]!=3'b101)
      | not_tmp_312;
  assign or_1217_nl = (STAGE_VEC_LOOP_j_sva_9_0[2:0]!=3'b101) | (COMP_LOOP_acc_10_psp_sva[0])
      | (fsm_output[2]) | not_tmp_311;
  assign or_1215_nl = (operator_64_false_acc_cse_8_sva[3:0]!=4'b0101) | (fsm_output[2])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]);
  assign mux_1418_nl = MUX_s_1_2_2(or_1217_nl, or_1215_nl, fsm_output[4]);
  assign mux_1419_nl = MUX_s_1_2_2(or_1219_nl, mux_1418_nl, fsm_output[8]);
  assign or_1213_nl = (operator_64_false_acc_cse_2_sva[3:0]!=4'b0101) | (fsm_output[2])
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign or_1212_nl = (COMP_LOOP_acc_7_psp_sva[2:0]!=3'b010) | (~ (STAGE_VEC_LOOP_j_sva_9_0[0]))
      | (fsm_output[2]) | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1417_nl = MUX_s_1_2_2(or_1213_nl, or_1212_nl, fsm_output[4]);
  assign or_1214_nl = (fsm_output[8]) | mux_1417_nl;
  assign mux_1420_nl = MUX_s_1_2_2(mux_1419_nl, or_1214_nl, fsm_output[1]);
  assign or_1210_nl = (COMP_LOOP_acc_12_psp_sva[1:0]!=2'b01) | (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b01)
      | (~ (fsm_output[2])) | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]);
  assign or_1209_nl = (operator_64_false_acc_cse_12_sva[3:0]!=4'b0101) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign mux_1415_nl = MUX_s_1_2_2(or_1210_nl, or_1209_nl, fsm_output[4]);
  assign or_1207_nl = (fsm_output[4]) | (operator_64_false_acc_cse_sva[3:0]!=4'b0101)
      | (fsm_output[2]) | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign mux_1416_nl = MUX_s_1_2_2(mux_1415_nl, or_1207_nl, fsm_output[8]);
  assign or_1211_nl = (fsm_output[1]) | mux_1416_nl;
  assign mux_1421_nl = MUX_s_1_2_2(mux_1420_nl, or_1211_nl, fsm_output[9]);
  assign mux_1431_nl = MUX_s_1_2_2(mux_1430_nl, mux_1421_nl, fsm_output[7]);
  assign mux_1447_nl = MUX_s_1_2_2(mux_1446_nl, mux_1431_nl, fsm_output[0]);
  assign vec_rsc_0_5_i_wea_d_pff = ~ mux_1447_nl;
  assign or_1311_nl = (operator_64_false_acc_cse_2_sva[3:0]!=4'b0101) | (fsm_output[4])
      | (fsm_output[0]) | (fsm_output[5]) | not_tmp_322;
  assign or_1309_nl = (COMP_LOOP_acc_cse_2_sva[3:0]!=4'b0101) | (~ (fsm_output[0]))
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[5])
      | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign or_1308_nl = (COMP_LOOP_1_operator_64_false_acc_tmp[3:0]!=4'b0101) | (fsm_output[5])
      | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign or_1307_nl = (STAGE_VEC_LOOP_j_sva_9_0[3:0]!=4'b0101) | (fsm_output[5])
      | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign mux_1477_nl = MUX_s_1_2_2(or_1308_nl, or_1307_nl, fsm_output[0]);
  assign mux_1478_nl = MUX_s_1_2_2(or_1309_nl, mux_1477_nl, fsm_output[4]);
  assign mux_1479_nl = MUX_s_1_2_2(or_1311_nl, mux_1478_nl, fsm_output[1]);
  assign or_1306_nl = (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b010) | (~ (STAGE_VEC_LOOP_j_sva_9_0[0]))
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[5])
      | not_tmp_322;
  assign or_1304_nl = (operator_64_false_acc_cse_11_sva[3:0]!=4'b0101) | (fsm_output[5])
      | not_tmp_322;
  assign mux_1474_nl = MUX_s_1_2_2(or_1306_nl, or_1304_nl, fsm_output[0]);
  assign or_1302_nl = (fsm_output[0]) | (operator_64_false_acc_cse_10_sva[3:0]!=4'b0101)
      | (fsm_output[5]) | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign mux_1475_nl = MUX_s_1_2_2(mux_1474_nl, or_1302_nl, fsm_output[4]);
  assign or_1300_nl = (COMP_LOOP_acc_cse_10_sva[3:0]!=4'b0101) | (~ (fsm_output[4]))
      | (~ (fsm_output[0])) | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      | (fsm_output[5]) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign mux_1476_nl = MUX_s_1_2_2(mux_1475_nl, or_1300_nl, fsm_output[1]);
  assign mux_1480_nl = MUX_s_1_2_2(mux_1479_nl, mux_1476_nl, fsm_output[9]);
  assign or_1299_nl = (COMP_LOOP_acc_9_psp_sva[2:0]!=3'b010) | (~ (STAGE_VEC_LOOP_j_sva_9_0[0]))
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (~
      (fsm_output[5])) | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign or_1298_nl = (operator_64_false_acc_cse_7_sva[3:0]!=4'b0101) | (~ (fsm_output[5]))
      | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign mux_1470_nl = MUX_s_1_2_2(or_1299_nl, or_1298_nl, fsm_output[0]);
  assign or_1297_nl = (operator_64_false_acc_cse_6_sva[3:0]!=4'b0101) | (fsm_output[0])
      | (~ (fsm_output[5])) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign mux_1471_nl = MUX_s_1_2_2(mux_1470_nl, or_1297_nl, fsm_output[4]);
  assign or_1296_nl = (COMP_LOOP_acc_cse_6_sva[3:0]!=4'b0101) | (fsm_output[4]) |
      (~ (fsm_output[0])) | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      | (fsm_output[6:5]!=2'b01) | nand_442_cse;
  assign mux_1472_nl = MUX_s_1_2_2(mux_1471_nl, or_1296_nl, fsm_output[1]);
  assign nand_346_nl = ~((COMP_LOOP_acc_cse_sva[3:0]==4'b0101) & operator_64_false_slc_operator_64_false_acc_1_60_itm
      & (fsm_output[0]) & (fsm_output[5]) & (fsm_output[6]) & (fsm_output[3]) & (~
      (fsm_output[2])));
  assign or_1293_nl = (COMP_LOOP_acc_13_psp_sva[2:0]!=3'b010) | (~ (STAGE_VEC_LOOP_j_sva_9_0[0]))
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (~
      (fsm_output[5])) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign or_1292_nl = (operator_64_false_acc_cse_15_sva[3:0]!=4'b0101) | (~ (fsm_output[5]))
      | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign mux_1467_nl = MUX_s_1_2_2(or_1293_nl, or_1292_nl, fsm_output[0]);
  assign mux_1468_nl = MUX_s_1_2_2(nand_346_nl, mux_1467_nl, fsm_output[4]);
  assign or_1291_nl = (operator_64_false_acc_cse_sva[3:0]!=4'b0101) | (fsm_output[4])
      | (fsm_output[0]) | (~ (fsm_output[5])) | (~ (fsm_output[6])) | (~ (fsm_output[3]))
      | (fsm_output[2]);
  assign mux_1469_nl = MUX_s_1_2_2(mux_1468_nl, or_1291_nl, fsm_output[1]);
  assign mux_1473_nl = MUX_s_1_2_2(mux_1472_nl, mux_1469_nl, fsm_output[9]);
  assign mux_1481_nl = MUX_s_1_2_2(mux_1480_nl, mux_1473_nl, fsm_output[8]);
  assign or_1290_nl = (COMP_LOOP_acc_7_psp_sva[2:0]!=3'b010) | (~ (STAGE_VEC_LOOP_j_sva_9_0[0]))
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[5])
      | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign or_1288_nl = (operator_64_false_acc_cse_3_sva[3:0]!=4'b0101) | (fsm_output[5])
      | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign mux_1462_nl = MUX_s_1_2_2(or_1290_nl, or_1288_nl, fsm_output[0]);
  assign or_1286_nl = (~ operator_64_false_slc_operator_64_false_acc_1_60_itm) |
      (COMP_LOOP_acc_cse_4_sva[3:0]!=4'b0101) | (~ (fsm_output[0])) | (~ (fsm_output[5]))
      | (fsm_output[6]) | nand_442_cse;
  assign mux_1463_nl = MUX_s_1_2_2(mux_1462_nl, or_1286_nl, fsm_output[4]);
  assign or_1284_nl = (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b01) | (COMP_LOOP_acc_8_psp_sva[1:0]!=2'b01)
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (~
      (fsm_output[5])) | (~ (fsm_output[6])) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign or_1282_nl = (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b01) | (COMP_LOOP_acc_8_psp_sva[1:0]!=2'b01)
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm);
  assign mux_1459_nl = MUX_s_1_2_2(nand_tmp_19, or_tmp_669, or_1282_nl);
  assign nor_299_nl = ~((operator_64_false_acc_cse_4_sva[3:0]!=4'b0101));
  assign mux_1460_nl = MUX_s_1_2_2(or_1284_nl, mux_1459_nl, nor_299_nl);
  assign or_1281_nl = (operator_64_false_acc_cse_5_sva[3:0]!=4'b0101) | (~ (fsm_output[5]))
      | (~ (fsm_output[6])) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign mux_1461_nl = MUX_s_1_2_2(mux_1460_nl, or_1281_nl, fsm_output[0]);
  assign nand_50_nl = ~((fsm_output[4]) & (~ mux_1461_nl));
  assign mux_1464_nl = MUX_s_1_2_2(mux_1463_nl, nand_50_nl, fsm_output[1]);
  assign or_1279_nl = (COMP_LOOP_acc_cse_12_sva[3:0]!=4'b0101) | (~ operator_64_false_slc_operator_64_false_acc_1_60_itm)
      | (~ (fsm_output[0])) | (fsm_output[5]) | (fsm_output[6]) | (fsm_output[3])
      | (~ (fsm_output[2]));
  assign or_1277_nl = (operator_64_false_acc_cse_14_sva[3:0]!=4'b0101) | (fsm_output[0])
      | (~ (fsm_output[5])) | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign mux_1457_nl = MUX_s_1_2_2(or_1279_nl, or_1277_nl, fsm_output[4]);
  assign or_1276_nl = (operator_64_false_acc_cse_12_sva[3:0]!=4'b0101) | (fsm_output[0])
      | (fsm_output[5]) | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign or_1274_nl = (COMP_LOOP_acc_12_psp_sva[1:0]!=2'b01) | (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b01)
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[6:5]!=2'b01)
      | nand_442_cse;
  assign or_1272_nl = (operator_64_false_acc_cse_13_sva[3:0]!=4'b0101) | (fsm_output[6:5]!=2'b01)
      | nand_442_cse;
  assign nor_297_nl = ~((operator_64_false_acc_cse_13_sva[3:0]!=4'b0101));
  assign mux_1453_nl = MUX_s_1_2_2(nand_437_cse, mux_1112_cse, nor_297_nl);
  assign nor_296_nl = ~((COMP_LOOP_acc_cse_14_sva[3:0]!=4'b0101));
  assign mux_1454_nl = MUX_s_1_2_2(or_1272_nl, mux_1453_nl, nor_296_nl);
  assign mux_1455_nl = MUX_s_1_2_2(or_1274_nl, mux_1454_nl, fsm_output[0]);
  assign mux_1456_nl = MUX_s_1_2_2(or_1276_nl, mux_1455_nl, fsm_output[4]);
  assign mux_1458_nl = MUX_s_1_2_2(mux_1457_nl, mux_1456_nl, fsm_output[1]);
  assign mux_1465_nl = MUX_s_1_2_2(mux_1464_nl, mux_1458_nl, fsm_output[9]);
  assign or_1264_nl = (COMP_LOOP_acc_cse_8_sva[3:0]!=4'b0101) | (fsm_output[4]) |
      (~ operator_64_false_slc_operator_64_false_acc_1_60_itm) | (~ (fsm_output[0]))
      | (~ (fsm_output[5])) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign or_1263_nl = (operator_64_false_acc_cse_8_sva[3:0]!=4'b0101) | (fsm_output[0])
      | (~ (fsm_output[5])) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign or_1262_nl = (STAGE_VEC_LOOP_j_sva_9_0[2:0]!=3'b101) | (COMP_LOOP_acc_10_psp_sva[0])
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[5])
      | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign or_1261_nl = (operator_64_false_acc_cse_9_sva[3:0]!=4'b0101) | (fsm_output[5])
      | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign mux_1448_nl = MUX_s_1_2_2(or_1262_nl, or_1261_nl, fsm_output[0]);
  assign mux_1449_nl = MUX_s_1_2_2(or_1263_nl, mux_1448_nl, fsm_output[4]);
  assign mux_1450_nl = MUX_s_1_2_2(or_1264_nl, mux_1449_nl, fsm_output[1]);
  assign or_1265_nl = (fsm_output[9]) | mux_1450_nl;
  assign mux_1466_nl = MUX_s_1_2_2(mux_1465_nl, or_1265_nl, fsm_output[8]);
  assign mux_1482_nl = MUX_s_1_2_2(mux_1481_nl, mux_1466_nl, fsm_output[7]);
  assign vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d = ~ mux_1482_nl;
  assign nor_693_nl = ~((operator_64_false_acc_cse_1_sva[3:0]!=4'b0110) | (fsm_output[2])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]));
  assign nor_694_nl = ~((COMP_LOOP_acc_cse_2_sva[3:0]!=4'b0110) | (fsm_output[2])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]));
  assign mux_1511_nl = MUX_s_1_2_2(nor_693_nl, nor_694_nl, fsm_output[4]);
  assign nor_695_nl = ~((operator_64_false_acc_cse_5_sva[3:0]!=4'b0110) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5])));
  assign nor_696_nl = ~((COMP_LOOP_acc_cse_6_sva[3:0]!=4'b0110) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5])));
  assign mux_1510_nl = MUX_s_1_2_2(nor_695_nl, nor_696_nl, fsm_output[4]);
  assign mux_1512_nl = MUX_s_1_2_2(mux_1511_nl, mux_1510_nl, fsm_output[8]);
  assign nand_54_nl = ~((fsm_output[1]) & mux_1512_nl);
  assign nor_697_nl = ~((operator_64_false_acc_cse_15_sva[3:0]!=4'b0110) | (fsm_output[2])
      | not_tmp_311);
  assign nor_698_nl = ~((COMP_LOOP_acc_cse_sva[3:0]!=4'b0110) | (fsm_output[2]) |
      not_tmp_311);
  assign mux_1508_nl = MUX_s_1_2_2(nor_697_nl, nor_698_nl, fsm_output[4]);
  assign nand_53_nl = ~((fsm_output[8]) & mux_1508_nl);
  assign or_1356_nl = (COMP_LOOP_acc_cse_10_sva[3:0]!=4'b0110) | (fsm_output[2])
      | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign or_1354_nl = (operator_64_false_acc_cse_9_sva[3:0]!=4'b0110) | (fsm_output[2])
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1506_nl = MUX_s_1_2_2(or_1356_nl, or_1354_nl, fsm_output[4]);
  assign or_1353_nl = (fsm_output[4]) | (COMP_LOOP_acc_cse_14_sva[3:0]!=4'b0110)
      | (~ (fsm_output[2])) | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1507_nl = MUX_s_1_2_2(mux_1506_nl, or_1353_nl, fsm_output[8]);
  assign mux_1509_nl = MUX_s_1_2_2(nand_53_nl, mux_1507_nl, fsm_output[1]);
  assign mux_1513_nl = MUX_s_1_2_2(nand_54_nl, mux_1509_nl, fsm_output[9]);
  assign or_1351_nl = (COMP_LOOP_acc_cse_4_sva[3:0]!=4'b0110) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]);
  assign or_1350_nl = (operator_64_false_acc_cse_3_sva[3:0]!=4'b0110) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign mux_1503_nl = MUX_s_1_2_2(or_1351_nl, or_1350_nl, fsm_output[4]);
  assign or_1348_nl = (operator_64_false_acc_cse_7_sva[3:0]!=4'b0110) | (fsm_output[2])
      | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign or_1346_nl = (COMP_LOOP_acc_cse_8_sva[3:0]!=4'b0110) | (fsm_output[2]) |
      (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign mux_1502_nl = MUX_s_1_2_2(or_1348_nl, or_1346_nl, fsm_output[4]);
  assign mux_1504_nl = MUX_s_1_2_2(mux_1503_nl, mux_1502_nl, fsm_output[8]);
  assign or_1352_nl = (fsm_output[1]) | mux_1504_nl;
  assign or_1343_nl = (operator_64_false_acc_cse_11_sva[3:0]!=4'b0110) | (~ (fsm_output[2]))
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign or_1342_nl = (COMP_LOOP_acc_cse_12_sva[3:0]!=4'b0110) | (~ (fsm_output[2]))
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1500_nl = MUX_s_1_2_2(or_1343_nl, or_1342_nl, fsm_output[4]);
  assign or_1344_nl = (fsm_output[8]) | mux_1500_nl;
  assign or_1341_nl = (operator_64_false_acc_cse_13_sva[3:0]!=4'b0110) | (fsm_output[8])
      | (~ (fsm_output[4])) | (~ (fsm_output[2])) | (fsm_output[3]) | not_tmp_312;
  assign mux_1501_nl = MUX_s_1_2_2(or_1344_nl, or_1341_nl, fsm_output[1]);
  assign mux_1505_nl = MUX_s_1_2_2(or_1352_nl, mux_1501_nl, fsm_output[9]);
  assign mux_1514_nl = MUX_s_1_2_2(mux_1513_nl, mux_1505_nl, fsm_output[7]);
  assign or_1337_nl = (COMP_LOOP_acc_8_psp_sva[1:0]!=2'b01) | (fsm_output[4]) | (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b10)
      | (~ (fsm_output[2])) | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1495_nl = MUX_s_1_2_2(or_1339_cse, or_1337_nl, fsm_output[8]);
  assign mux_1496_nl = MUX_s_1_2_2(mux_1495_nl, nand_tmp_52, fsm_output[1]);
  assign or_1336_nl = (~ (fsm_output[8])) | (COMP_LOOP_acc_8_psp_sva[1:0]!=2'b01)
      | (fsm_output[4]) | (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b10) | (~ (fsm_output[2]))
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1494_nl = MUX_s_1_2_2(or_1336_nl, nand_tmp_52, fsm_output[1]);
  assign mux_1497_nl = MUX_s_1_2_2(mux_1496_nl, mux_1494_nl, STAGE_VEC_LOOP_j_sva_9_0[3]);
  assign nor_699_nl = ~((operator_64_false_acc_cse_10_sva[3:0]!=4'b0110) | (fsm_output[2])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]));
  assign nor_700_nl = ~((COMP_LOOP_acc_11_psp_sva[2:0]!=3'b011) | (STAGE_VEC_LOOP_j_sva_9_0[0])
      | (fsm_output[2]) | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]));
  assign mux_1491_nl = MUX_s_1_2_2(nor_699_nl, nor_700_nl, fsm_output[4]);
  assign nor_701_nl = ~((operator_64_false_acc_cse_14_sva[3:0]!=4'b0110) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5])));
  assign nor_702_nl = ~((COMP_LOOP_acc_13_psp_sva[2:0]!=3'b011) | (STAGE_VEC_LOOP_j_sva_9_0[0])
      | (~ (fsm_output[2])) | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5])));
  assign mux_1490_nl = MUX_s_1_2_2(nor_701_nl, nor_702_nl, fsm_output[4]);
  assign mux_1492_nl = MUX_s_1_2_2(mux_1491_nl, mux_1490_nl, fsm_output[8]);
  assign nand_51_nl = ~((fsm_output[1]) & mux_1492_nl);
  assign mux_1498_nl = MUX_s_1_2_2(mux_1497_nl, nand_51_nl, fsm_output[9]);
  assign or_1325_nl = (operator_64_false_acc_cse_4_sva[3:0]!=4'b0110) | (fsm_output[4:2]!=3'b101)
      | not_tmp_312;
  assign or_1323_nl = (STAGE_VEC_LOOP_j_sva_9_0[2:0]!=3'b110) | (COMP_LOOP_acc_10_psp_sva[0])
      | (fsm_output[2]) | not_tmp_311;
  assign or_1321_nl = (operator_64_false_acc_cse_8_sva[3:0]!=4'b0110) | (fsm_output[2])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]);
  assign mux_1486_nl = MUX_s_1_2_2(or_1323_nl, or_1321_nl, fsm_output[4]);
  assign mux_1487_nl = MUX_s_1_2_2(or_1325_nl, mux_1486_nl, fsm_output[8]);
  assign or_1319_nl = (operator_64_false_acc_cse_2_sva[3:0]!=4'b0110) | (fsm_output[2])
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign or_1318_nl = (COMP_LOOP_acc_7_psp_sva[2:0]!=3'b011) | (STAGE_VEC_LOOP_j_sva_9_0[0])
      | (fsm_output[2]) | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1485_nl = MUX_s_1_2_2(or_1319_nl, or_1318_nl, fsm_output[4]);
  assign or_1320_nl = (fsm_output[8]) | mux_1485_nl;
  assign mux_1488_nl = MUX_s_1_2_2(mux_1487_nl, or_1320_nl, fsm_output[1]);
  assign or_1316_nl = (COMP_LOOP_acc_12_psp_sva[1:0]!=2'b01) | (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b10)
      | (~ (fsm_output[2])) | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]);
  assign or_1315_nl = (operator_64_false_acc_cse_12_sva[3:0]!=4'b0110) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign mux_1483_nl = MUX_s_1_2_2(or_1316_nl, or_1315_nl, fsm_output[4]);
  assign or_1313_nl = (fsm_output[4]) | (operator_64_false_acc_cse_sva[3:0]!=4'b0110)
      | (fsm_output[2]) | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign mux_1484_nl = MUX_s_1_2_2(mux_1483_nl, or_1313_nl, fsm_output[8]);
  assign or_1317_nl = (fsm_output[1]) | mux_1484_nl;
  assign mux_1489_nl = MUX_s_1_2_2(mux_1488_nl, or_1317_nl, fsm_output[9]);
  assign mux_1499_nl = MUX_s_1_2_2(mux_1498_nl, mux_1489_nl, fsm_output[7]);
  assign mux_1515_nl = MUX_s_1_2_2(mux_1514_nl, mux_1499_nl, fsm_output[0]);
  assign vec_rsc_0_6_i_wea_d_pff = ~ mux_1515_nl;
  assign or_1420_nl = (operator_64_false_acc_cse_2_sva[3:0]!=4'b0110) | (fsm_output[4])
      | (fsm_output[0]) | (fsm_output[5]) | not_tmp_322;
  assign or_1418_nl = (COMP_LOOP_acc_cse_2_sva[3:0]!=4'b0110) | (~ (fsm_output[0]))
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[5])
      | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign or_1417_nl = (COMP_LOOP_1_operator_64_false_acc_tmp[3:0]!=4'b0110) | (fsm_output[5])
      | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign or_1416_nl = (STAGE_VEC_LOOP_j_sva_9_0[3:0]!=4'b0110) | (fsm_output[5])
      | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign mux_1545_nl = MUX_s_1_2_2(or_1417_nl, or_1416_nl, fsm_output[0]);
  assign mux_1546_nl = MUX_s_1_2_2(or_1418_nl, mux_1545_nl, fsm_output[4]);
  assign mux_1547_nl = MUX_s_1_2_2(or_1420_nl, mux_1546_nl, fsm_output[1]);
  assign or_1415_nl = (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b011) | (STAGE_VEC_LOOP_j_sva_9_0[0])
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[5])
      | not_tmp_322;
  assign or_1413_nl = (operator_64_false_acc_cse_11_sva[3:0]!=4'b0110) | (fsm_output[5])
      | not_tmp_322;
  assign mux_1542_nl = MUX_s_1_2_2(or_1415_nl, or_1413_nl, fsm_output[0]);
  assign or_1411_nl = (fsm_output[0]) | (operator_64_false_acc_cse_10_sva[3:0]!=4'b0110)
      | (fsm_output[5]) | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign mux_1543_nl = MUX_s_1_2_2(mux_1542_nl, or_1411_nl, fsm_output[4]);
  assign or_1409_nl = (~ (fsm_output[4])) | (~ (fsm_output[0])) | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      | (COMP_LOOP_acc_cse_10_sva[3:0]!=4'b0110) | (fsm_output[5]) | (fsm_output[6])
      | (fsm_output[3]) | (fsm_output[2]);
  assign mux_1544_nl = MUX_s_1_2_2(mux_1543_nl, or_1409_nl, fsm_output[1]);
  assign mux_1548_nl = MUX_s_1_2_2(mux_1547_nl, mux_1544_nl, fsm_output[9]);
  assign or_1408_nl = (COMP_LOOP_acc_9_psp_sva[2:0]!=3'b011) | (STAGE_VEC_LOOP_j_sva_9_0[0])
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (~
      (fsm_output[5])) | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign or_1407_nl = (operator_64_false_acc_cse_7_sva[3:0]!=4'b0110) | (~ (fsm_output[5]))
      | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign mux_1538_nl = MUX_s_1_2_2(or_1408_nl, or_1407_nl, fsm_output[0]);
  assign or_1406_nl = (operator_64_false_acc_cse_6_sva[3:0]!=4'b0110) | (fsm_output[0])
      | (~ (fsm_output[5])) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign mux_1539_nl = MUX_s_1_2_2(mux_1538_nl, or_1406_nl, fsm_output[4]);
  assign or_1405_nl = (COMP_LOOP_acc_cse_6_sva[3:0]!=4'b0110) | (fsm_output[4]) |
      (~ (fsm_output[0])) | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      | (fsm_output[6:5]!=2'b01) | nand_442_cse;
  assign mux_1540_nl = MUX_s_1_2_2(mux_1539_nl, or_1405_nl, fsm_output[1]);
  assign nand_340_nl = ~(operator_64_false_slc_operator_64_false_acc_1_60_itm & (fsm_output[0])
      & (COMP_LOOP_acc_cse_sva[3:0]==4'b0110) & (fsm_output[5]) & (fsm_output[6])
      & (fsm_output[3]) & (~ (fsm_output[2])));
  assign or_1402_nl = (COMP_LOOP_acc_13_psp_sva[2:0]!=3'b011) | (STAGE_VEC_LOOP_j_sva_9_0[0])
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (~
      (fsm_output[5])) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign or_1401_nl = (operator_64_false_acc_cse_15_sva[3:0]!=4'b0110) | (~ (fsm_output[5]))
      | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign mux_1535_nl = MUX_s_1_2_2(or_1402_nl, or_1401_nl, fsm_output[0]);
  assign mux_1536_nl = MUX_s_1_2_2(nand_340_nl, mux_1535_nl, fsm_output[4]);
  assign or_1400_nl = (operator_64_false_acc_cse_sva[3:0]!=4'b0110) | (fsm_output[4])
      | (fsm_output[0]) | (~ (fsm_output[5])) | (~ (fsm_output[6])) | (~ (fsm_output[3]))
      | (fsm_output[2]);
  assign mux_1537_nl = MUX_s_1_2_2(mux_1536_nl, or_1400_nl, fsm_output[1]);
  assign mux_1541_nl = MUX_s_1_2_2(mux_1540_nl, mux_1537_nl, fsm_output[9]);
  assign mux_1549_nl = MUX_s_1_2_2(mux_1548_nl, mux_1541_nl, fsm_output[8]);
  assign or_1399_nl = (COMP_LOOP_acc_7_psp_sva[2:0]!=3'b011) | (STAGE_VEC_LOOP_j_sva_9_0[0])
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[5])
      | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign or_1397_nl = (operator_64_false_acc_cse_3_sva[3:0]!=4'b0110) | (fsm_output[5])
      | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign mux_1530_nl = MUX_s_1_2_2(or_1399_nl, or_1397_nl, fsm_output[0]);
  assign or_1395_nl = (~ operator_64_false_slc_operator_64_false_acc_1_60_itm) |
      (COMP_LOOP_acc_cse_4_sva[3:0]!=4'b0110) | (~ (fsm_output[0])) | (~ (fsm_output[5]))
      | (fsm_output[6]) | nand_442_cse;
  assign mux_1531_nl = MUX_s_1_2_2(mux_1530_nl, or_1395_nl, fsm_output[4]);
  assign or_1393_nl = (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b10) | (COMP_LOOP_acc_8_psp_sva[1:0]!=2'b01)
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm);
  assign mux_1527_nl = MUX_s_1_2_2(nand_tmp_19, or_tmp_669, or_1393_nl);
  assign or_1392_nl = (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b10) | (COMP_LOOP_acc_8_psp_sva[1:0]!=2'b01)
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (~
      (fsm_output[5])) | (~ (fsm_output[6])) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign or_1390_nl = (operator_64_false_acc_cse_4_sva[3:0]!=4'b0110);
  assign mux_1528_nl = MUX_s_1_2_2(mux_1527_nl, or_1392_nl, or_1390_nl);
  assign or_1389_nl = (operator_64_false_acc_cse_5_sva[3:0]!=4'b0110) | (~ (fsm_output[5]))
      | (~ (fsm_output[6])) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign mux_1529_nl = MUX_s_1_2_2(mux_1528_nl, or_1389_nl, fsm_output[0]);
  assign nand_56_nl = ~((fsm_output[4]) & (~ mux_1529_nl));
  assign mux_1532_nl = MUX_s_1_2_2(mux_1531_nl, nand_56_nl, fsm_output[1]);
  assign or_1387_nl = (~ operator_64_false_slc_operator_64_false_acc_1_60_itm) |
      (~ (fsm_output[0])) | (COMP_LOOP_acc_cse_12_sva[3:0]!=4'b0110) | (fsm_output[5])
      | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign or_1385_nl = (operator_64_false_acc_cse_14_sva[3:0]!=4'b0110) | (fsm_output[0])
      | (~ (fsm_output[5])) | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign mux_1525_nl = MUX_s_1_2_2(or_1387_nl, or_1385_nl, fsm_output[4]);
  assign or_1384_nl = (operator_64_false_acc_cse_12_sva[3:0]!=4'b0110) | (fsm_output[0])
      | (fsm_output[5]) | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign or_1382_nl = (COMP_LOOP_acc_12_psp_sva[1:0]!=2'b01) | (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b10)
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[6:5]!=2'b01)
      | nand_442_cse;
  assign or_1375_nl = (operator_64_false_acc_cse_13_sva[3:0]!=4'b0110);
  assign mux_1521_nl = MUX_s_1_2_2(mux_1112_cse, nand_437_cse, or_1375_nl);
  assign or_1374_nl = (operator_64_false_acc_cse_13_sva[3:0]!=4'b0110) | (fsm_output[6:5]!=2'b01)
      | nand_442_cse;
  assign or_1372_nl = (COMP_LOOP_acc_cse_14_sva[3:0]!=4'b0110);
  assign mux_1522_nl = MUX_s_1_2_2(mux_1521_nl, or_1374_nl, or_1372_nl);
  assign mux_1523_nl = MUX_s_1_2_2(or_1382_nl, mux_1522_nl, fsm_output[0]);
  assign mux_1524_nl = MUX_s_1_2_2(or_1384_nl, mux_1523_nl, fsm_output[4]);
  assign mux_1526_nl = MUX_s_1_2_2(mux_1525_nl, mux_1524_nl, fsm_output[1]);
  assign mux_1533_nl = MUX_s_1_2_2(mux_1532_nl, mux_1526_nl, fsm_output[9]);
  assign or_1370_nl = (COMP_LOOP_acc_cse_8_sva[3:0]!=4'b0110) | (fsm_output[4]) |
      (~ operator_64_false_slc_operator_64_false_acc_1_60_itm) | (~ (fsm_output[0]))
      | (~ (fsm_output[5])) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign or_1369_nl = (operator_64_false_acc_cse_8_sva[3:0]!=4'b0110) | (fsm_output[0])
      | (~ (fsm_output[5])) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign or_1368_nl = (STAGE_VEC_LOOP_j_sva_9_0[2:0]!=3'b110) | (COMP_LOOP_acc_10_psp_sva[0])
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[5])
      | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign or_1367_nl = (operator_64_false_acc_cse_9_sva[3:0]!=4'b0110) | (fsm_output[5])
      | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign mux_1516_nl = MUX_s_1_2_2(or_1368_nl, or_1367_nl, fsm_output[0]);
  assign mux_1517_nl = MUX_s_1_2_2(or_1369_nl, mux_1516_nl, fsm_output[4]);
  assign mux_1518_nl = MUX_s_1_2_2(or_1370_nl, mux_1517_nl, fsm_output[1]);
  assign or_1371_nl = (fsm_output[9]) | mux_1518_nl;
  assign mux_1534_nl = MUX_s_1_2_2(mux_1533_nl, or_1371_nl, fsm_output[8]);
  assign mux_1550_nl = MUX_s_1_2_2(mux_1549_nl, mux_1534_nl, fsm_output[7]);
  assign vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d = ~ mux_1550_nl;
  assign nor_681_nl = ~((operator_64_false_acc_cse_1_sva[3:0]!=4'b0111) | (fsm_output[2])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]));
  assign nor_682_nl = ~((COMP_LOOP_acc_cse_2_sva[3:0]!=4'b0111) | (fsm_output[2])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]));
  assign mux_1579_nl = MUX_s_1_2_2(nor_681_nl, nor_682_nl, fsm_output[4]);
  assign and_773_nl = (operator_64_false_acc_cse_5_sva[3:0]==4'b0111) & (fsm_output[2])
      & (fsm_output[3]) & (~ (fsm_output[6])) & (fsm_output[5]);
  assign and_779_nl = (COMP_LOOP_acc_cse_6_sva[3:0]==4'b0111) & (fsm_output[2]) &
      (fsm_output[3]) & (~ (fsm_output[6])) & (fsm_output[5]);
  assign mux_1578_nl = MUX_s_1_2_2(and_773_nl, and_779_nl, fsm_output[4]);
  assign mux_1580_nl = MUX_s_1_2_2(mux_1579_nl, mux_1578_nl, fsm_output[8]);
  assign nand_60_nl = ~((fsm_output[1]) & mux_1580_nl);
  assign nor_685_nl = ~((operator_64_false_acc_cse_15_sva[3:0]!=4'b0111) | (fsm_output[2])
      | not_tmp_311);
  assign nor_686_nl = ~((COMP_LOOP_acc_cse_sva[3:0]!=4'b0111) | (fsm_output[2]) |
      not_tmp_311);
  assign mux_1576_nl = MUX_s_1_2_2(nor_685_nl, nor_686_nl, fsm_output[4]);
  assign nand_59_nl = ~((fsm_output[8]) & mux_1576_nl);
  assign or_1465_nl = (COMP_LOOP_acc_cse_10_sva[3:0]!=4'b0111) | (fsm_output[2])
      | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign or_1463_nl = (operator_64_false_acc_cse_9_sva[3:0]!=4'b0111) | (fsm_output[2])
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1574_nl = MUX_s_1_2_2(or_1465_nl, or_1463_nl, fsm_output[4]);
  assign or_1462_nl = (fsm_output[4]) | (COMP_LOOP_acc_cse_14_sva[3:0]!=4'b0111)
      | (~ (fsm_output[2])) | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1575_nl = MUX_s_1_2_2(mux_1574_nl, or_1462_nl, fsm_output[8]);
  assign mux_1577_nl = MUX_s_1_2_2(nand_59_nl, mux_1575_nl, fsm_output[1]);
  assign mux_1581_nl = MUX_s_1_2_2(nand_60_nl, mux_1577_nl, fsm_output[9]);
  assign nand_331_nl = ~((COMP_LOOP_acc_cse_4_sva[3:0]==4'b0111) & (fsm_output[2])
      & (fsm_output[3]) & (fsm_output[6]) & (~ (fsm_output[5])));
  assign nand_472_nl = ~((operator_64_false_acc_cse_3_sva[3:0]==4'b0111) & (fsm_output[2])
      & (fsm_output[3]) & (~ (fsm_output[6])) & (fsm_output[5]));
  assign mux_1571_nl = MUX_s_1_2_2(nand_331_nl, nand_472_nl, fsm_output[4]);
  assign or_1457_nl = (operator_64_false_acc_cse_7_sva[3:0]!=4'b0111) | (fsm_output[2])
      | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign or_1455_nl = (COMP_LOOP_acc_cse_8_sva[3:0]!=4'b0111) | (fsm_output[2]) |
      (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign mux_1570_nl = MUX_s_1_2_2(or_1457_nl, or_1455_nl, fsm_output[4]);
  assign mux_1572_nl = MUX_s_1_2_2(mux_1571_nl, mux_1570_nl, fsm_output[8]);
  assign or_1461_nl = (fsm_output[1]) | mux_1572_nl;
  assign or_1452_nl = (operator_64_false_acc_cse_11_sva[3:0]!=4'b0111) | (~ (fsm_output[2]))
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign or_1451_nl = (COMP_LOOP_acc_cse_12_sva[3:0]!=4'b0111) | (~ (fsm_output[2]))
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1568_nl = MUX_s_1_2_2(or_1452_nl, or_1451_nl, fsm_output[4]);
  assign or_1453_nl = (fsm_output[8]) | mux_1568_nl;
  assign or_1450_nl = (operator_64_false_acc_cse_13_sva[3:0]!=4'b0111) | (fsm_output[8])
      | (~ (fsm_output[4])) | (~ (fsm_output[2])) | (fsm_output[3]) | not_tmp_312;
  assign mux_1569_nl = MUX_s_1_2_2(or_1453_nl, or_1450_nl, fsm_output[1]);
  assign mux_1573_nl = MUX_s_1_2_2(or_1461_nl, mux_1569_nl, fsm_output[9]);
  assign mux_1582_nl = MUX_s_1_2_2(mux_1581_nl, mux_1573_nl, fsm_output[7]);
  assign or_1446_nl = (COMP_LOOP_acc_8_psp_sva[1:0]!=2'b01) | (fsm_output[4]) | (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b11)
      | (~ (fsm_output[2])) | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1563_nl = MUX_s_1_2_2(or_1448_cse, or_1446_nl, fsm_output[8]);
  assign mux_1564_nl = MUX_s_1_2_2(mux_1563_nl, nand_tmp_58, fsm_output[1]);
  assign or_1445_nl = (~ (fsm_output[8])) | (COMP_LOOP_acc_8_psp_sva[1:0]!=2'b01)
      | (fsm_output[4]) | (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b11) | (~ (fsm_output[2]))
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1562_nl = MUX_s_1_2_2(or_1445_nl, nand_tmp_58, fsm_output[1]);
  assign mux_1565_nl = MUX_s_1_2_2(mux_1564_nl, mux_1562_nl, STAGE_VEC_LOOP_j_sva_9_0[3]);
  assign nor_687_nl = ~((operator_64_false_acc_cse_10_sva[3:0]!=4'b0111) | (fsm_output[2])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]));
  assign nor_688_nl = ~((COMP_LOOP_acc_11_psp_sva[2:0]!=3'b011) | (~ (STAGE_VEC_LOOP_j_sva_9_0[0]))
      | (fsm_output[2]) | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]));
  assign mux_1559_nl = MUX_s_1_2_2(nor_687_nl, nor_688_nl, fsm_output[4]);
  assign and_789_nl = (operator_64_false_acc_cse_14_sva[3:0]==4'b0111) & (fsm_output[2])
      & (fsm_output[3]) & (~ (fsm_output[6])) & (fsm_output[5]);
  assign and_790_nl = (COMP_LOOP_acc_13_psp_sva[2:0]==3'b011) & (STAGE_VEC_LOOP_j_sva_9_0[0])
      & (fsm_output[2]) & (fsm_output[3]) & (~ (fsm_output[6])) & (fsm_output[5]);
  assign mux_1558_nl = MUX_s_1_2_2(and_789_nl, and_790_nl, fsm_output[4]);
  assign mux_1560_nl = MUX_s_1_2_2(mux_1559_nl, mux_1558_nl, fsm_output[8]);
  assign nand_57_nl = ~((fsm_output[1]) & mux_1560_nl);
  assign mux_1566_nl = MUX_s_1_2_2(mux_1565_nl, nand_57_nl, fsm_output[9]);
  assign or_1434_nl = (~((operator_64_false_acc_cse_4_sva[3:0]==4'b0111) & (fsm_output[4:2]==3'b101)))
      | not_tmp_312;
  assign or_1432_nl = (STAGE_VEC_LOOP_j_sva_9_0[2:0]!=3'b111) | (COMP_LOOP_acc_10_psp_sva[0])
      | (fsm_output[2]) | not_tmp_311;
  assign or_1430_nl = (operator_64_false_acc_cse_8_sva[3:0]!=4'b0111) | (fsm_output[2])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]);
  assign mux_1554_nl = MUX_s_1_2_2(or_1432_nl, or_1430_nl, fsm_output[4]);
  assign mux_1555_nl = MUX_s_1_2_2(or_1434_nl, mux_1554_nl, fsm_output[8]);
  assign or_1428_nl = (operator_64_false_acc_cse_2_sva[3:0]!=4'b0111) | (fsm_output[2])
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign or_1427_nl = (COMP_LOOP_acc_7_psp_sva[2:0]!=3'b011) | (~ (STAGE_VEC_LOOP_j_sva_9_0[0]))
      | (fsm_output[2]) | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1553_nl = MUX_s_1_2_2(or_1428_nl, or_1427_nl, fsm_output[4]);
  assign or_1429_nl = (fsm_output[8]) | mux_1553_nl;
  assign mux_1556_nl = MUX_s_1_2_2(mux_1555_nl, or_1429_nl, fsm_output[1]);
  assign nand_336_nl = ~((COMP_LOOP_acc_12_psp_sva[1:0]==2'b01) & (STAGE_VEC_LOOP_j_sva_9_0[1:0]==2'b11)
      & (fsm_output[2]) & (fsm_output[3]) & (fsm_output[6]) & (~ (fsm_output[5])));
  assign nand_453_nl = ~((operator_64_false_acc_cse_12_sva[3:0]==4'b0111) & (fsm_output[2])
      & (fsm_output[3]) & (~ (fsm_output[6])) & (fsm_output[5]));
  assign mux_1551_nl = MUX_s_1_2_2(nand_336_nl, nand_453_nl, fsm_output[4]);
  assign or_1422_nl = (fsm_output[4]) | (operator_64_false_acc_cse_sva[3:0]!=4'b0111)
      | (fsm_output[2]) | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign mux_1552_nl = MUX_s_1_2_2(mux_1551_nl, or_1422_nl, fsm_output[8]);
  assign or_1426_nl = (fsm_output[1]) | mux_1552_nl;
  assign mux_1557_nl = MUX_s_1_2_2(mux_1556_nl, or_1426_nl, fsm_output[9]);
  assign mux_1567_nl = MUX_s_1_2_2(mux_1566_nl, mux_1557_nl, fsm_output[7]);
  assign mux_1583_nl = MUX_s_1_2_2(mux_1582_nl, mux_1567_nl, fsm_output[0]);
  assign vec_rsc_0_7_i_wea_d_pff = ~ mux_1583_nl;
  assign or_1526_nl = (operator_64_false_acc_cse_2_sva[3:0]!=4'b0111) | (fsm_output[4])
      | (fsm_output[0]) | (fsm_output[5]) | not_tmp_322;
  assign nand_317_nl = ~((COMP_LOOP_acc_cse_2_sva[3:0]==4'b0111) & (fsm_output[0])
      & COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm & (~ (fsm_output[5]))
      & (fsm_output[6]) & (fsm_output[3]) & (~ (fsm_output[2])));
  assign or_1523_nl = (COMP_LOOP_1_operator_64_false_acc_tmp[3:0]!=4'b0111) | (fsm_output[5])
      | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign or_1522_nl = (STAGE_VEC_LOOP_j_sva_9_0[3:0]!=4'b0111) | (fsm_output[5])
      | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign mux_1613_nl = MUX_s_1_2_2(or_1523_nl, or_1522_nl, fsm_output[0]);
  assign mux_1614_nl = MUX_s_1_2_2(nand_317_nl, mux_1613_nl, fsm_output[4]);
  assign mux_1615_nl = MUX_s_1_2_2(or_1526_nl, mux_1614_nl, fsm_output[1]);
  assign or_1521_nl = (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b011) | (~ (STAGE_VEC_LOOP_j_sva_9_0[0]))
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[5])
      | not_tmp_322;
  assign or_1519_nl = (operator_64_false_acc_cse_11_sva[3:0]!=4'b0111) | (fsm_output[5])
      | not_tmp_322;
  assign mux_1610_nl = MUX_s_1_2_2(or_1521_nl, or_1519_nl, fsm_output[0]);
  assign or_1517_nl = (fsm_output[0]) | (operator_64_false_acc_cse_10_sva[3:0]!=4'b0111)
      | (fsm_output[5]) | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign mux_1611_nl = MUX_s_1_2_2(mux_1610_nl, or_1517_nl, fsm_output[4]);
  assign or_1515_nl = (COMP_LOOP_acc_cse_10_sva[3:0]!=4'b0111) | (~ (fsm_output[4]))
      | (~ (fsm_output[0])) | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      | (fsm_output[5]) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign mux_1612_nl = MUX_s_1_2_2(mux_1611_nl, or_1515_nl, fsm_output[1]);
  assign mux_1616_nl = MUX_s_1_2_2(mux_1615_nl, mux_1612_nl, fsm_output[9]);
  assign nand_318_nl = ~((COMP_LOOP_acc_9_psp_sva[2:0]==3'b011) & (STAGE_VEC_LOOP_j_sva_9_0[0])
      & COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm & (fsm_output[5])
      & (fsm_output[6]) & (fsm_output[3]) & (~ (fsm_output[2])));
  assign nand_319_nl = ~((operator_64_false_acc_cse_7_sva[3:0]==4'b0111) & (fsm_output[5])
      & (fsm_output[6]) & (fsm_output[3]) & (~ (fsm_output[2])));
  assign mux_1606_nl = MUX_s_1_2_2(nand_318_nl, nand_319_nl, fsm_output[0]);
  assign or_1512_nl = (operator_64_false_acc_cse_6_sva[3:0]!=4'b0111) | (fsm_output[0])
      | (~ (fsm_output[5])) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign mux_1607_nl = MUX_s_1_2_2(mux_1606_nl, or_1512_nl, fsm_output[4]);
  assign or_1511_nl = (COMP_LOOP_acc_cse_6_sva[3:0]!=4'b0111) | (fsm_output[4]) |
      (~ (fsm_output[0])) | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      | (fsm_output[6:5]!=2'b01) | nand_442_cse;
  assign mux_1608_nl = MUX_s_1_2_2(mux_1607_nl, or_1511_nl, fsm_output[1]);
  assign nand_320_nl = ~(operator_64_false_slc_operator_64_false_acc_1_60_itm & (fsm_output[0])
      & (COMP_LOOP_acc_cse_sva[3:0]==4'b0111) & (fsm_output[5]) & (fsm_output[6])
      & (fsm_output[3]) & (~ (fsm_output[2])));
  assign or_1508_nl = (COMP_LOOP_acc_13_psp_sva[2:0]!=3'b011) | (~ (STAGE_VEC_LOOP_j_sva_9_0[0]))
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (~
      (fsm_output[5])) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign or_1507_nl = (operator_64_false_acc_cse_15_sva[3:0]!=4'b0111) | (~ (fsm_output[5]))
      | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign mux_1603_nl = MUX_s_1_2_2(or_1508_nl, or_1507_nl, fsm_output[0]);
  assign mux_1604_nl = MUX_s_1_2_2(nand_320_nl, mux_1603_nl, fsm_output[4]);
  assign or_1506_nl = (operator_64_false_acc_cse_sva[3:0]!=4'b0111) | (fsm_output[4])
      | (fsm_output[0]) | (~ (fsm_output[5])) | (~ (fsm_output[6])) | (~ (fsm_output[3]))
      | (fsm_output[2]);
  assign mux_1605_nl = MUX_s_1_2_2(mux_1604_nl, or_1506_nl, fsm_output[1]);
  assign mux_1609_nl = MUX_s_1_2_2(mux_1608_nl, mux_1605_nl, fsm_output[9]);
  assign mux_1617_nl = MUX_s_1_2_2(mux_1616_nl, mux_1609_nl, fsm_output[8]);
  assign or_1505_nl = (COMP_LOOP_acc_7_psp_sva[2:0]!=3'b011) | (~ (STAGE_VEC_LOOP_j_sva_9_0[0]))
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[5])
      | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign or_1503_nl = (operator_64_false_acc_cse_3_sva[3:0]!=4'b0111) | (fsm_output[5])
      | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign mux_1598_nl = MUX_s_1_2_2(or_1505_nl, or_1503_nl, fsm_output[0]);
  assign or_1501_nl = (~(operator_64_false_slc_operator_64_false_acc_1_60_itm & (COMP_LOOP_acc_cse_4_sva[3:0]==4'b0111)
      & (fsm_output[0]) & (fsm_output[5]) & (~ (fsm_output[6])))) | nand_442_cse;
  assign mux_1599_nl = MUX_s_1_2_2(mux_1598_nl, or_1501_nl, fsm_output[4]);
  assign nand_467_nl = ~((STAGE_VEC_LOOP_j_sva_9_0[1:0]==2'b11) & (COMP_LOOP_acc_8_psp_sva[1:0]==2'b01)
      & COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm & (fsm_output[5])
      & (fsm_output[6]) & (~ (fsm_output[3])) & (fsm_output[2]));
  assign nand_323_nl = ~((STAGE_VEC_LOOP_j_sva_9_0[1:0]==2'b11) & (COMP_LOOP_acc_8_psp_sva[1:0]==2'b01)
      & COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm);
  assign mux_1595_nl = MUX_s_1_2_2(nand_tmp_19, or_tmp_669, nand_323_nl);
  assign and_546_nl = (operator_64_false_acc_cse_4_sva[3:0]==4'b0111);
  assign mux_1596_nl = MUX_s_1_2_2(nand_467_nl, mux_1595_nl, and_546_nl);
  assign nand_463_nl = ~((operator_64_false_acc_cse_5_sva[3:0]==4'b0111) & (fsm_output[5])
      & (fsm_output[6]) & (~ (fsm_output[3])) & (fsm_output[2]));
  assign mux_1597_nl = MUX_s_1_2_2(mux_1596_nl, nand_463_nl, fsm_output[0]);
  assign nand_62_nl = ~((fsm_output[4]) & (~ mux_1597_nl));
  assign mux_1600_nl = MUX_s_1_2_2(mux_1599_nl, nand_62_nl, fsm_output[1]);
  assign or_1494_nl = (~ operator_64_false_slc_operator_64_false_acc_1_60_itm) |
      (~ (fsm_output[0])) | (COMP_LOOP_acc_cse_12_sva[3:0]!=4'b0111) | (fsm_output[5])
      | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign or_1492_nl = (operator_64_false_acc_cse_14_sva[3:0]!=4'b0111) | (fsm_output[0])
      | (~ (fsm_output[5])) | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign mux_1593_nl = MUX_s_1_2_2(or_1494_nl, or_1492_nl, fsm_output[4]);
  assign or_1491_nl = (operator_64_false_acc_cse_12_sva[3:0]!=4'b0111) | (fsm_output[0])
      | (fsm_output[5]) | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign or_1489_nl = (~((COMP_LOOP_acc_12_psp_sva[1:0]==2'b01) & (STAGE_VEC_LOOP_j_sva_9_0[1:0]==2'b11)
      & COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm & (fsm_output[6:5]==2'b01)))
      | nand_442_cse;
  assign or_1487_nl = (operator_64_false_acc_cse_13_sva[3:0]!=4'b0111) | (fsm_output[6:5]!=2'b01)
      | nand_442_cse;
  assign and_547_nl = (operator_64_false_acc_cse_13_sva[3:0]==4'b0111);
  assign mux_1589_nl = MUX_s_1_2_2(nand_437_cse, mux_1112_cse, and_547_nl);
  assign and_548_nl = (COMP_LOOP_acc_cse_14_sva[3:0]==4'b0111);
  assign mux_1590_nl = MUX_s_1_2_2(or_1487_nl, mux_1589_nl, and_548_nl);
  assign mux_1591_nl = MUX_s_1_2_2(or_1489_nl, mux_1590_nl, fsm_output[0]);
  assign mux_1592_nl = MUX_s_1_2_2(or_1491_nl, mux_1591_nl, fsm_output[4]);
  assign mux_1594_nl = MUX_s_1_2_2(mux_1593_nl, mux_1592_nl, fsm_output[1]);
  assign mux_1601_nl = MUX_s_1_2_2(mux_1600_nl, mux_1594_nl, fsm_output[9]);
  assign or_1479_nl = (COMP_LOOP_acc_cse_8_sva[3:0]!=4'b0111) | (fsm_output[4]) |
      (~ operator_64_false_slc_operator_64_false_acc_1_60_itm) | (~ (fsm_output[0]))
      | (~ (fsm_output[5])) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign or_1478_nl = (operator_64_false_acc_cse_8_sva[3:0]!=4'b0111) | (fsm_output[0])
      | (~ (fsm_output[5])) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign or_1477_nl = (STAGE_VEC_LOOP_j_sva_9_0[2:0]!=3'b111) | (COMP_LOOP_acc_10_psp_sva[0])
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[5])
      | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign or_1476_nl = (operator_64_false_acc_cse_9_sva[3:0]!=4'b0111) | (fsm_output[5])
      | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign mux_1584_nl = MUX_s_1_2_2(or_1477_nl, or_1476_nl, fsm_output[0]);
  assign mux_1585_nl = MUX_s_1_2_2(or_1478_nl, mux_1584_nl, fsm_output[4]);
  assign mux_1586_nl = MUX_s_1_2_2(or_1479_nl, mux_1585_nl, fsm_output[1]);
  assign or_1480_nl = (fsm_output[9]) | mux_1586_nl;
  assign mux_1602_nl = MUX_s_1_2_2(mux_1601_nl, or_1480_nl, fsm_output[8]);
  assign mux_1618_nl = MUX_s_1_2_2(mux_1617_nl, mux_1602_nl, fsm_output[7]);
  assign vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d = ~ mux_1618_nl;
  assign nor_669_nl = ~((operator_64_false_acc_cse_1_sva[3:0]!=4'b1000) | (fsm_output[2])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]));
  assign nor_670_nl = ~((COMP_LOOP_acc_cse_2_sva[3:0]!=4'b1000) | (fsm_output[2])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]));
  assign mux_1647_nl = MUX_s_1_2_2(nor_669_nl, nor_670_nl, fsm_output[4]);
  assign nor_671_nl = ~((operator_64_false_acc_cse_5_sva[3:0]!=4'b1000) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5])));
  assign nor_672_nl = ~((COMP_LOOP_acc_cse_6_sva[3:0]!=4'b1000) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5])));
  assign mux_1646_nl = MUX_s_1_2_2(nor_671_nl, nor_672_nl, fsm_output[4]);
  assign mux_1648_nl = MUX_s_1_2_2(mux_1647_nl, mux_1646_nl, fsm_output[8]);
  assign nand_66_nl = ~((fsm_output[1]) & mux_1648_nl);
  assign nor_673_nl = ~((operator_64_false_acc_cse_15_sva[3:0]!=4'b1000) | (fsm_output[2])
      | not_tmp_311);
  assign nor_674_nl = ~((COMP_LOOP_acc_cse_sva[3:0]!=4'b1000) | (fsm_output[2]) |
      not_tmp_311);
  assign mux_1644_nl = MUX_s_1_2_2(nor_673_nl, nor_674_nl, fsm_output[4]);
  assign nand_65_nl = ~((fsm_output[8]) & mux_1644_nl);
  assign or_1571_nl = (COMP_LOOP_acc_cse_10_sva[3:0]!=4'b1000) | (fsm_output[2])
      | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign or_1569_nl = (operator_64_false_acc_cse_9_sva[3:0]!=4'b1000) | (fsm_output[2])
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1642_nl = MUX_s_1_2_2(or_1571_nl, or_1569_nl, fsm_output[4]);
  assign or_1568_nl = (fsm_output[4]) | (COMP_LOOP_acc_cse_14_sva[3:0]!=4'b1000)
      | (~ (fsm_output[2])) | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1643_nl = MUX_s_1_2_2(mux_1642_nl, or_1568_nl, fsm_output[8]);
  assign mux_1645_nl = MUX_s_1_2_2(nand_65_nl, mux_1643_nl, fsm_output[1]);
  assign mux_1649_nl = MUX_s_1_2_2(nand_66_nl, mux_1645_nl, fsm_output[9]);
  assign or_1566_nl = (COMP_LOOP_acc_cse_4_sva[3:0]!=4'b1000) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]);
  assign or_1565_nl = (operator_64_false_acc_cse_3_sva[3:0]!=4'b1000) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign mux_1639_nl = MUX_s_1_2_2(or_1566_nl, or_1565_nl, fsm_output[4]);
  assign or_1563_nl = (operator_64_false_acc_cse_7_sva[3:0]!=4'b1000) | (fsm_output[2])
      | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign or_1561_nl = (COMP_LOOP_acc_cse_8_sva[3:0]!=4'b1000) | (fsm_output[2]) |
      (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign mux_1638_nl = MUX_s_1_2_2(or_1563_nl, or_1561_nl, fsm_output[4]);
  assign mux_1640_nl = MUX_s_1_2_2(mux_1639_nl, mux_1638_nl, fsm_output[8]);
  assign or_1567_nl = (fsm_output[1]) | mux_1640_nl;
  assign or_1558_nl = (operator_64_false_acc_cse_11_sva[3:0]!=4'b1000) | (~ (fsm_output[2]))
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign or_1557_nl = (COMP_LOOP_acc_cse_12_sva[3:0]!=4'b1000) | (~ (fsm_output[2]))
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1636_nl = MUX_s_1_2_2(or_1558_nl, or_1557_nl, fsm_output[4]);
  assign or_1559_nl = (fsm_output[8]) | mux_1636_nl;
  assign or_1556_nl = (operator_64_false_acc_cse_13_sva[3:0]!=4'b1000) | (fsm_output[8])
      | (~ (fsm_output[4])) | (~ (fsm_output[2])) | (fsm_output[3]) | not_tmp_312;
  assign mux_1637_nl = MUX_s_1_2_2(or_1559_nl, or_1556_nl, fsm_output[1]);
  assign mux_1641_nl = MUX_s_1_2_2(or_1567_nl, mux_1637_nl, fsm_output[9]);
  assign mux_1650_nl = MUX_s_1_2_2(mux_1649_nl, mux_1641_nl, fsm_output[7]);
  assign or_1554_nl = (~ (fsm_output[8])) | (COMP_LOOP_acc_8_psp_sva[1:0]!=2'b10)
      | (fsm_output[4]) | (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b00) | (~ (fsm_output[2]))
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1632_nl = MUX_s_1_2_2(or_1554_nl, nand_tmp_64, fsm_output[1]);
  assign or_1551_nl = (COMP_LOOP_acc_8_psp_sva[1:0]!=2'b10) | (fsm_output[4]) | (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b00)
      | (~ (fsm_output[2])) | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1630_nl = MUX_s_1_2_2(or_694_cse, or_1551_nl, fsm_output[8]);
  assign mux_1631_nl = MUX_s_1_2_2(mux_1630_nl, nand_tmp_64, fsm_output[1]);
  assign mux_1633_nl = MUX_s_1_2_2(mux_1632_nl, mux_1631_nl, STAGE_VEC_LOOP_j_sva_9_0[3]);
  assign nor_675_nl = ~((operator_64_false_acc_cse_10_sva[3:0]!=4'b1000) | (fsm_output[2])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]));
  assign nor_676_nl = ~((COMP_LOOP_acc_11_psp_sva[2:0]!=3'b100) | (STAGE_VEC_LOOP_j_sva_9_0[0])
      | (fsm_output[2]) | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]));
  assign mux_1627_nl = MUX_s_1_2_2(nor_675_nl, nor_676_nl, fsm_output[4]);
  assign nor_677_nl = ~((operator_64_false_acc_cse_14_sva[3:0]!=4'b1000) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5])));
  assign nor_678_nl = ~((COMP_LOOP_acc_13_psp_sva[2:0]!=3'b100) | (STAGE_VEC_LOOP_j_sva_9_0[0])
      | (~ (fsm_output[2])) | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5])));
  assign mux_1626_nl = MUX_s_1_2_2(nor_677_nl, nor_678_nl, fsm_output[4]);
  assign mux_1628_nl = MUX_s_1_2_2(mux_1627_nl, mux_1626_nl, fsm_output[8]);
  assign nand_63_nl = ~((fsm_output[1]) & mux_1628_nl);
  assign mux_1634_nl = MUX_s_1_2_2(mux_1633_nl, nand_63_nl, fsm_output[9]);
  assign or_1540_nl = (operator_64_false_acc_cse_4_sva[3:0]!=4'b1000) | (fsm_output[4:2]!=3'b101)
      | not_tmp_312;
  assign or_1538_nl = (STAGE_VEC_LOOP_j_sva_9_0[2:0]!=3'b000) | (~ (COMP_LOOP_acc_10_psp_sva[0]))
      | (fsm_output[2]) | not_tmp_311;
  assign or_1536_nl = (operator_64_false_acc_cse_8_sva[3:0]!=4'b1000) | (fsm_output[2])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]);
  assign mux_1622_nl = MUX_s_1_2_2(or_1538_nl, or_1536_nl, fsm_output[4]);
  assign mux_1623_nl = MUX_s_1_2_2(or_1540_nl, mux_1622_nl, fsm_output[8]);
  assign or_1534_nl = (operator_64_false_acc_cse_2_sva[3:0]!=4'b1000) | (fsm_output[2])
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign or_1533_nl = (COMP_LOOP_acc_7_psp_sva[2:0]!=3'b100) | (STAGE_VEC_LOOP_j_sva_9_0[0])
      | (fsm_output[2]) | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1621_nl = MUX_s_1_2_2(or_1534_nl, or_1533_nl, fsm_output[4]);
  assign or_1535_nl = (fsm_output[8]) | mux_1621_nl;
  assign mux_1624_nl = MUX_s_1_2_2(mux_1623_nl, or_1535_nl, fsm_output[1]);
  assign or_1531_nl = (COMP_LOOP_acc_12_psp_sva[1:0]!=2'b10) | (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b00)
      | (~ (fsm_output[2])) | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]);
  assign or_1530_nl = (operator_64_false_acc_cse_12_sva[3:0]!=4'b1000) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign mux_1619_nl = MUX_s_1_2_2(or_1531_nl, or_1530_nl, fsm_output[4]);
  assign or_1528_nl = (fsm_output[4]) | (operator_64_false_acc_cse_sva[3:0]!=4'b1000)
      | (fsm_output[2]) | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign mux_1620_nl = MUX_s_1_2_2(mux_1619_nl, or_1528_nl, fsm_output[8]);
  assign or_1532_nl = (fsm_output[1]) | mux_1620_nl;
  assign mux_1625_nl = MUX_s_1_2_2(mux_1624_nl, or_1532_nl, fsm_output[9]);
  assign mux_1635_nl = MUX_s_1_2_2(mux_1634_nl, mux_1625_nl, fsm_output[7]);
  assign mux_1651_nl = MUX_s_1_2_2(mux_1650_nl, mux_1635_nl, fsm_output[0]);
  assign vec_rsc_0_8_i_wea_d_pff = ~ mux_1651_nl;
  assign or_1635_nl = (operator_64_false_acc_cse_2_sva[3:0]!=4'b1000) | (fsm_output[4])
      | (fsm_output[0]) | (fsm_output[5]) | not_tmp_322;
  assign or_1633_nl = (COMP_LOOP_acc_cse_2_sva[3:0]!=4'b1000) | (~ (fsm_output[0]))
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[5])
      | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign or_1632_nl = (COMP_LOOP_1_operator_64_false_acc_tmp[3:0]!=4'b1000) | (fsm_output[5])
      | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign or_1631_nl = (STAGE_VEC_LOOP_j_sva_9_0[3:0]!=4'b1000) | (fsm_output[5])
      | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign mux_1681_nl = MUX_s_1_2_2(or_1632_nl, or_1631_nl, fsm_output[0]);
  assign mux_1682_nl = MUX_s_1_2_2(or_1633_nl, mux_1681_nl, fsm_output[4]);
  assign mux_1683_nl = MUX_s_1_2_2(or_1635_nl, mux_1682_nl, fsm_output[1]);
  assign or_1630_nl = (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b100) | (STAGE_VEC_LOOP_j_sva_9_0[0])
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[5])
      | not_tmp_322;
  assign or_1628_nl = (operator_64_false_acc_cse_11_sva[3:0]!=4'b1000) | (fsm_output[5])
      | not_tmp_322;
  assign mux_1678_nl = MUX_s_1_2_2(or_1630_nl, or_1628_nl, fsm_output[0]);
  assign or_1626_nl = (fsm_output[0]) | (operator_64_false_acc_cse_10_sva[3:0]!=4'b1000)
      | (fsm_output[5]) | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign mux_1679_nl = MUX_s_1_2_2(mux_1678_nl, or_1626_nl, fsm_output[4]);
  assign or_1624_nl = (~ (fsm_output[4])) | (~ (fsm_output[0])) | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      | (COMP_LOOP_acc_cse_10_sva[3:0]!=4'b1000) | (fsm_output[5]) | (fsm_output[6])
      | (fsm_output[3]) | (fsm_output[2]);
  assign mux_1680_nl = MUX_s_1_2_2(mux_1679_nl, or_1624_nl, fsm_output[1]);
  assign mux_1684_nl = MUX_s_1_2_2(mux_1683_nl, mux_1680_nl, fsm_output[9]);
  assign or_1623_nl = (COMP_LOOP_acc_9_psp_sva[2:0]!=3'b100) | (STAGE_VEC_LOOP_j_sva_9_0[0])
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (~
      (fsm_output[5])) | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign or_1622_nl = (operator_64_false_acc_cse_7_sva[3:0]!=4'b1000) | (~ (fsm_output[5]))
      | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign mux_1674_nl = MUX_s_1_2_2(or_1623_nl, or_1622_nl, fsm_output[0]);
  assign or_1621_nl = (operator_64_false_acc_cse_6_sva[3:0]!=4'b1000) | (fsm_output[0])
      | (~ (fsm_output[5])) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign mux_1675_nl = MUX_s_1_2_2(mux_1674_nl, or_1621_nl, fsm_output[4]);
  assign or_1620_nl = (COMP_LOOP_acc_cse_6_sva[3:0]!=4'b1000) | (fsm_output[4]) |
      (~ (fsm_output[0])) | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      | (fsm_output[6:5]!=2'b01) | nand_442_cse;
  assign mux_1676_nl = MUX_s_1_2_2(mux_1675_nl, or_1620_nl, fsm_output[1]);
  assign or_1618_nl = (COMP_LOOP_acc_cse_sva[3:0]!=4'b1000) | (~ operator_64_false_slc_operator_64_false_acc_1_60_itm)
      | (~ (fsm_output[0])) | (~ (fsm_output[5])) | (~ (fsm_output[6])) | (~ (fsm_output[3]))
      | (fsm_output[2]);
  assign or_1617_nl = (COMP_LOOP_acc_13_psp_sva[2:0]!=3'b100) | (STAGE_VEC_LOOP_j_sva_9_0[0])
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (~
      (fsm_output[5])) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign or_1616_nl = (operator_64_false_acc_cse_15_sva[3:0]!=4'b1000) | (~ (fsm_output[5]))
      | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign mux_1671_nl = MUX_s_1_2_2(or_1617_nl, or_1616_nl, fsm_output[0]);
  assign mux_1672_nl = MUX_s_1_2_2(or_1618_nl, mux_1671_nl, fsm_output[4]);
  assign or_1615_nl = (operator_64_false_acc_cse_sva[3:0]!=4'b1000) | (fsm_output[4])
      | (fsm_output[0]) | (~ (fsm_output[5])) | (~ (fsm_output[6])) | (~ (fsm_output[3]))
      | (fsm_output[2]);
  assign mux_1673_nl = MUX_s_1_2_2(mux_1672_nl, or_1615_nl, fsm_output[1]);
  assign mux_1677_nl = MUX_s_1_2_2(mux_1676_nl, mux_1673_nl, fsm_output[9]);
  assign mux_1685_nl = MUX_s_1_2_2(mux_1684_nl, mux_1677_nl, fsm_output[8]);
  assign or_1614_nl = (COMP_LOOP_acc_7_psp_sva[2:0]!=3'b100) | (STAGE_VEC_LOOP_j_sva_9_0[0])
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[5])
      | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign or_1612_nl = (operator_64_false_acc_cse_3_sva[3:0]!=4'b1000) | (fsm_output[5])
      | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign mux_1666_nl = MUX_s_1_2_2(or_1614_nl, or_1612_nl, fsm_output[0]);
  assign or_1610_nl = (~ operator_64_false_slc_operator_64_false_acc_1_60_itm) |
      (COMP_LOOP_acc_cse_4_sva[3:0]!=4'b1000) | (~ (fsm_output[0])) | (~ (fsm_output[5]))
      | (fsm_output[6]) | nand_442_cse;
  assign mux_1667_nl = MUX_s_1_2_2(mux_1666_nl, or_1610_nl, fsm_output[4]);
  assign or_1608_nl = (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b00) | (COMP_LOOP_acc_8_psp_sva[1:0]!=2'b10)
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm);
  assign mux_1663_nl = MUX_s_1_2_2(nand_tmp_19, or_tmp_669, or_1608_nl);
  assign or_1607_nl = (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b00) | (COMP_LOOP_acc_8_psp_sva[1:0]!=2'b10)
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (~
      (fsm_output[5])) | (~ (fsm_output[6])) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign or_1605_nl = (operator_64_false_acc_cse_4_sva[3:0]!=4'b1000);
  assign mux_1664_nl = MUX_s_1_2_2(mux_1663_nl, or_1607_nl, or_1605_nl);
  assign or_1604_nl = (operator_64_false_acc_cse_5_sva[3:0]!=4'b1000) | (~ (fsm_output[5]))
      | (~ (fsm_output[6])) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign mux_1665_nl = MUX_s_1_2_2(mux_1664_nl, or_1604_nl, fsm_output[0]);
  assign nand_68_nl = ~((fsm_output[4]) & (~ mux_1665_nl));
  assign mux_1668_nl = MUX_s_1_2_2(mux_1667_nl, nand_68_nl, fsm_output[1]);
  assign or_1602_nl = (COMP_LOOP_acc_cse_12_sva[3:0]!=4'b1000) | (~ operator_64_false_slc_operator_64_false_acc_1_60_itm)
      | (~ (fsm_output[0])) | (fsm_output[5]) | (fsm_output[6]) | (fsm_output[3])
      | (~ (fsm_output[2]));
  assign or_1600_nl = (operator_64_false_acc_cse_14_sva[3:0]!=4'b1000) | (fsm_output[0])
      | (~ (fsm_output[5])) | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign mux_1661_nl = MUX_s_1_2_2(or_1602_nl, or_1600_nl, fsm_output[4]);
  assign or_1599_nl = (operator_64_false_acc_cse_12_sva[3:0]!=4'b1000) | (fsm_output[0])
      | (fsm_output[5]) | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign or_1597_nl = (COMP_LOOP_acc_12_psp_sva[1:0]!=2'b10) | (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b00)
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[6:5]!=2'b01)
      | nand_442_cse;
  assign or_1590_nl = (operator_64_false_acc_cse_13_sva[3:0]!=4'b1000);
  assign mux_1657_nl = MUX_s_1_2_2(mux_1112_cse, nand_437_cse, or_1590_nl);
  assign or_1589_nl = (operator_64_false_acc_cse_13_sva[3:0]!=4'b1000) | (fsm_output[6:5]!=2'b01)
      | nand_442_cse;
  assign or_1587_nl = (COMP_LOOP_acc_cse_14_sva[3:0]!=4'b1000);
  assign mux_1658_nl = MUX_s_1_2_2(mux_1657_nl, or_1589_nl, or_1587_nl);
  assign mux_1659_nl = MUX_s_1_2_2(or_1597_nl, mux_1658_nl, fsm_output[0]);
  assign mux_1660_nl = MUX_s_1_2_2(or_1599_nl, mux_1659_nl, fsm_output[4]);
  assign mux_1662_nl = MUX_s_1_2_2(mux_1661_nl, mux_1660_nl, fsm_output[1]);
  assign mux_1669_nl = MUX_s_1_2_2(mux_1668_nl, mux_1662_nl, fsm_output[9]);
  assign or_1585_nl = (COMP_LOOP_acc_cse_8_sva[3:0]!=4'b1000) | (fsm_output[4]) |
      (~ operator_64_false_slc_operator_64_false_acc_1_60_itm) | (~ (fsm_output[0]))
      | (~ (fsm_output[5])) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign or_1584_nl = (operator_64_false_acc_cse_8_sva[3:0]!=4'b1000) | (fsm_output[0])
      | (~ (fsm_output[5])) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign or_1583_nl = (STAGE_VEC_LOOP_j_sva_9_0[2:0]!=3'b000) | (~ (COMP_LOOP_acc_10_psp_sva[0]))
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[5])
      | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign or_1582_nl = (operator_64_false_acc_cse_9_sva[3:0]!=4'b1000) | (fsm_output[5])
      | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign mux_1652_nl = MUX_s_1_2_2(or_1583_nl, or_1582_nl, fsm_output[0]);
  assign mux_1653_nl = MUX_s_1_2_2(or_1584_nl, mux_1652_nl, fsm_output[4]);
  assign mux_1654_nl = MUX_s_1_2_2(or_1585_nl, mux_1653_nl, fsm_output[1]);
  assign or_1586_nl = (fsm_output[9]) | mux_1654_nl;
  assign mux_1670_nl = MUX_s_1_2_2(mux_1669_nl, or_1586_nl, fsm_output[8]);
  assign mux_1686_nl = MUX_s_1_2_2(mux_1685_nl, mux_1670_nl, fsm_output[7]);
  assign vec_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d = ~ mux_1686_nl;
  assign nor_657_nl = ~((operator_64_false_acc_cse_1_sva[3:0]!=4'b1001) | (fsm_output[2])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]));
  assign nor_658_nl = ~((COMP_LOOP_acc_cse_2_sva[3:0]!=4'b1001) | (fsm_output[2])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]));
  assign mux_1715_nl = MUX_s_1_2_2(nor_657_nl, nor_658_nl, fsm_output[4]);
  assign nor_659_nl = ~((operator_64_false_acc_cse_5_sva[3:0]!=4'b1001) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5])));
  assign nor_660_nl = ~((COMP_LOOP_acc_cse_6_sva[3:0]!=4'b1001) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5])));
  assign mux_1714_nl = MUX_s_1_2_2(nor_659_nl, nor_660_nl, fsm_output[4]);
  assign mux_1716_nl = MUX_s_1_2_2(mux_1715_nl, mux_1714_nl, fsm_output[8]);
  assign nand_72_nl = ~((fsm_output[1]) & mux_1716_nl);
  assign nor_661_nl = ~((operator_64_false_acc_cse_15_sva[3:0]!=4'b1001) | (fsm_output[2])
      | not_tmp_311);
  assign nor_662_nl = ~((COMP_LOOP_acc_cse_sva[3:0]!=4'b1001) | (fsm_output[2]) |
      not_tmp_311);
  assign mux_1712_nl = MUX_s_1_2_2(nor_661_nl, nor_662_nl, fsm_output[4]);
  assign nand_71_nl = ~((fsm_output[8]) & mux_1712_nl);
  assign or_1680_nl = (COMP_LOOP_acc_cse_10_sva[3:0]!=4'b1001) | (fsm_output[2])
      | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign or_1678_nl = (operator_64_false_acc_cse_9_sva[3:0]!=4'b1001) | (fsm_output[2])
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1710_nl = MUX_s_1_2_2(or_1680_nl, or_1678_nl, fsm_output[4]);
  assign or_1677_nl = (fsm_output[4]) | (COMP_LOOP_acc_cse_14_sva[3:0]!=4'b1001)
      | (~ (fsm_output[2])) | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1711_nl = MUX_s_1_2_2(mux_1710_nl, or_1677_nl, fsm_output[8]);
  assign mux_1713_nl = MUX_s_1_2_2(nand_71_nl, mux_1711_nl, fsm_output[1]);
  assign mux_1717_nl = MUX_s_1_2_2(nand_72_nl, mux_1713_nl, fsm_output[9]);
  assign or_1675_nl = (COMP_LOOP_acc_cse_4_sva[3:0]!=4'b1001) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]);
  assign or_1674_nl = (operator_64_false_acc_cse_3_sva[3:0]!=4'b1001) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign mux_1707_nl = MUX_s_1_2_2(or_1675_nl, or_1674_nl, fsm_output[4]);
  assign or_1672_nl = (operator_64_false_acc_cse_7_sva[3:0]!=4'b1001) | (fsm_output[2])
      | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign or_1670_nl = (COMP_LOOP_acc_cse_8_sva[3:0]!=4'b1001) | (fsm_output[2]) |
      (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign mux_1706_nl = MUX_s_1_2_2(or_1672_nl, or_1670_nl, fsm_output[4]);
  assign mux_1708_nl = MUX_s_1_2_2(mux_1707_nl, mux_1706_nl, fsm_output[8]);
  assign or_1676_nl = (fsm_output[1]) | mux_1708_nl;
  assign or_1667_nl = (operator_64_false_acc_cse_11_sva[3:0]!=4'b1001) | (~ (fsm_output[2]))
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign or_1666_nl = (COMP_LOOP_acc_cse_12_sva[3:0]!=4'b1001) | (~ (fsm_output[2]))
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1704_nl = MUX_s_1_2_2(or_1667_nl, or_1666_nl, fsm_output[4]);
  assign or_1668_nl = (fsm_output[8]) | mux_1704_nl;
  assign or_1665_nl = (operator_64_false_acc_cse_13_sva[3:0]!=4'b1001) | (fsm_output[8])
      | (~ (fsm_output[4])) | (~ (fsm_output[2])) | (fsm_output[3]) | not_tmp_312;
  assign mux_1705_nl = MUX_s_1_2_2(or_1668_nl, or_1665_nl, fsm_output[1]);
  assign mux_1709_nl = MUX_s_1_2_2(or_1676_nl, mux_1705_nl, fsm_output[9]);
  assign mux_1718_nl = MUX_s_1_2_2(mux_1717_nl, mux_1709_nl, fsm_output[7]);
  assign or_1663_nl = (~ (fsm_output[8])) | (COMP_LOOP_acc_8_psp_sva[1:0]!=2'b10)
      | (fsm_output[4]) | (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b01) | (~ (fsm_output[2]))
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1700_nl = MUX_s_1_2_2(or_1663_nl, nand_tmp_70, fsm_output[1]);
  assign or_1660_nl = (COMP_LOOP_acc_8_psp_sva[1:0]!=2'b10) | (fsm_output[4]) | (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b01)
      | (~ (fsm_output[2])) | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1698_nl = MUX_s_1_2_2(or_803_cse, or_1660_nl, fsm_output[8]);
  assign mux_1699_nl = MUX_s_1_2_2(mux_1698_nl, nand_tmp_70, fsm_output[1]);
  assign mux_1701_nl = MUX_s_1_2_2(mux_1700_nl, mux_1699_nl, STAGE_VEC_LOOP_j_sva_9_0[3]);
  assign nor_663_nl = ~((operator_64_false_acc_cse_10_sva[3:0]!=4'b1001) | (fsm_output[2])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]));
  assign nor_664_nl = ~((COMP_LOOP_acc_11_psp_sva[2:0]!=3'b100) | (~ (STAGE_VEC_LOOP_j_sva_9_0[0]))
      | (fsm_output[2]) | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]));
  assign mux_1695_nl = MUX_s_1_2_2(nor_663_nl, nor_664_nl, fsm_output[4]);
  assign nor_665_nl = ~((operator_64_false_acc_cse_14_sva[3:0]!=4'b1001) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5])));
  assign nor_666_nl = ~((COMP_LOOP_acc_13_psp_sva[2:0]!=3'b100) | (~ (STAGE_VEC_LOOP_j_sva_9_0[0]))
      | (~ (fsm_output[2])) | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5])));
  assign mux_1694_nl = MUX_s_1_2_2(nor_665_nl, nor_666_nl, fsm_output[4]);
  assign mux_1696_nl = MUX_s_1_2_2(mux_1695_nl, mux_1694_nl, fsm_output[8]);
  assign nand_69_nl = ~((fsm_output[1]) & mux_1696_nl);
  assign mux_1702_nl = MUX_s_1_2_2(mux_1701_nl, nand_69_nl, fsm_output[9]);
  assign or_1649_nl = (operator_64_false_acc_cse_4_sva[3:0]!=4'b1001) | (fsm_output[4:2]!=3'b101)
      | not_tmp_312;
  assign or_1647_nl = (STAGE_VEC_LOOP_j_sva_9_0[2:0]!=3'b001) | (~ (COMP_LOOP_acc_10_psp_sva[0]))
      | (fsm_output[2]) | not_tmp_311;
  assign or_1645_nl = (operator_64_false_acc_cse_8_sva[3:0]!=4'b1001) | (fsm_output[2])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]);
  assign mux_1690_nl = MUX_s_1_2_2(or_1647_nl, or_1645_nl, fsm_output[4]);
  assign mux_1691_nl = MUX_s_1_2_2(or_1649_nl, mux_1690_nl, fsm_output[8]);
  assign or_1643_nl = (operator_64_false_acc_cse_2_sva[3:0]!=4'b1001) | (fsm_output[2])
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign or_1642_nl = (COMP_LOOP_acc_7_psp_sva[2:0]!=3'b100) | (~ (STAGE_VEC_LOOP_j_sva_9_0[0]))
      | (fsm_output[2]) | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1689_nl = MUX_s_1_2_2(or_1643_nl, or_1642_nl, fsm_output[4]);
  assign or_1644_nl = (fsm_output[8]) | mux_1689_nl;
  assign mux_1692_nl = MUX_s_1_2_2(mux_1691_nl, or_1644_nl, fsm_output[1]);
  assign or_1640_nl = (COMP_LOOP_acc_12_psp_sva[1:0]!=2'b10) | (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b01)
      | (~ (fsm_output[2])) | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]);
  assign or_1639_nl = (operator_64_false_acc_cse_12_sva[3:0]!=4'b1001) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign mux_1687_nl = MUX_s_1_2_2(or_1640_nl, or_1639_nl, fsm_output[4]);
  assign or_1637_nl = (fsm_output[4]) | (operator_64_false_acc_cse_sva[3:0]!=4'b1001)
      | (fsm_output[2]) | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign mux_1688_nl = MUX_s_1_2_2(mux_1687_nl, or_1637_nl, fsm_output[8]);
  assign or_1641_nl = (fsm_output[1]) | mux_1688_nl;
  assign mux_1693_nl = MUX_s_1_2_2(mux_1692_nl, or_1641_nl, fsm_output[9]);
  assign mux_1703_nl = MUX_s_1_2_2(mux_1702_nl, mux_1693_nl, fsm_output[7]);
  assign mux_1719_nl = MUX_s_1_2_2(mux_1718_nl, mux_1703_nl, fsm_output[0]);
  assign vec_rsc_0_9_i_wea_d_pff = ~ mux_1719_nl;
  assign or_1741_nl = (operator_64_false_acc_cse_2_sva[3:0]!=4'b1001) | (fsm_output[4])
      | (fsm_output[0]) | (fsm_output[5]) | not_tmp_322;
  assign or_1739_nl = (COMP_LOOP_acc_cse_2_sva[3:0]!=4'b1001) | (~ (fsm_output[0]))
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[5])
      | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign or_1738_nl = (COMP_LOOP_1_operator_64_false_acc_tmp[3:0]!=4'b1001) | (fsm_output[5])
      | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign or_1737_nl = (STAGE_VEC_LOOP_j_sva_9_0[3:0]!=4'b1001) | (fsm_output[5])
      | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign mux_1749_nl = MUX_s_1_2_2(or_1738_nl, or_1737_nl, fsm_output[0]);
  assign mux_1750_nl = MUX_s_1_2_2(or_1739_nl, mux_1749_nl, fsm_output[4]);
  assign mux_1751_nl = MUX_s_1_2_2(or_1741_nl, mux_1750_nl, fsm_output[1]);
  assign or_1736_nl = (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b100) | (~ (STAGE_VEC_LOOP_j_sva_9_0[0]))
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[5])
      | not_tmp_322;
  assign or_1734_nl = (operator_64_false_acc_cse_11_sva[3:0]!=4'b1001) | (fsm_output[5])
      | not_tmp_322;
  assign mux_1746_nl = MUX_s_1_2_2(or_1736_nl, or_1734_nl, fsm_output[0]);
  assign or_1732_nl = (fsm_output[0]) | (operator_64_false_acc_cse_10_sva[3:0]!=4'b1001)
      | (fsm_output[5]) | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign mux_1747_nl = MUX_s_1_2_2(mux_1746_nl, or_1732_nl, fsm_output[4]);
  assign or_1730_nl = (COMP_LOOP_acc_cse_10_sva[3:0]!=4'b1001) | (~ (fsm_output[4]))
      | (~ (fsm_output[0])) | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      | (fsm_output[5]) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign mux_1748_nl = MUX_s_1_2_2(mux_1747_nl, or_1730_nl, fsm_output[1]);
  assign mux_1752_nl = MUX_s_1_2_2(mux_1751_nl, mux_1748_nl, fsm_output[9]);
  assign or_1729_nl = (COMP_LOOP_acc_9_psp_sva[2:0]!=3'b100) | (~ (STAGE_VEC_LOOP_j_sva_9_0[0]))
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (~
      (fsm_output[5])) | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign or_1728_nl = (operator_64_false_acc_cse_7_sva[3:0]!=4'b1001) | (~ (fsm_output[5]))
      | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign mux_1742_nl = MUX_s_1_2_2(or_1729_nl, or_1728_nl, fsm_output[0]);
  assign or_1727_nl = (operator_64_false_acc_cse_6_sva[3:0]!=4'b1001) | (fsm_output[0])
      | (~ (fsm_output[5])) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign mux_1743_nl = MUX_s_1_2_2(mux_1742_nl, or_1727_nl, fsm_output[4]);
  assign or_1726_nl = (COMP_LOOP_acc_cse_6_sva[3:0]!=4'b1001) | (fsm_output[4]) |
      (~ (fsm_output[0])) | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      | (fsm_output[6:5]!=2'b01) | nand_442_cse;
  assign mux_1744_nl = MUX_s_1_2_2(mux_1743_nl, or_1726_nl, fsm_output[1]);
  assign nand_306_nl = ~((COMP_LOOP_acc_cse_sva[3:0]==4'b1001) & operator_64_false_slc_operator_64_false_acc_1_60_itm
      & (fsm_output[0]) & (fsm_output[5]) & (fsm_output[6]) & (fsm_output[3]) & (~
      (fsm_output[2])));
  assign or_1723_nl = (COMP_LOOP_acc_13_psp_sva[2:0]!=3'b100) | (~ (STAGE_VEC_LOOP_j_sva_9_0[0]))
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (~
      (fsm_output[5])) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign or_1722_nl = (operator_64_false_acc_cse_15_sva[3:0]!=4'b1001) | (~ (fsm_output[5]))
      | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign mux_1739_nl = MUX_s_1_2_2(or_1723_nl, or_1722_nl, fsm_output[0]);
  assign mux_1740_nl = MUX_s_1_2_2(nand_306_nl, mux_1739_nl, fsm_output[4]);
  assign or_1721_nl = (operator_64_false_acc_cse_sva[3:0]!=4'b1001) | (fsm_output[4])
      | (fsm_output[0]) | (~ (fsm_output[5])) | (~ (fsm_output[6])) | (~ (fsm_output[3]))
      | (fsm_output[2]);
  assign mux_1741_nl = MUX_s_1_2_2(mux_1740_nl, or_1721_nl, fsm_output[1]);
  assign mux_1745_nl = MUX_s_1_2_2(mux_1744_nl, mux_1741_nl, fsm_output[9]);
  assign mux_1753_nl = MUX_s_1_2_2(mux_1752_nl, mux_1745_nl, fsm_output[8]);
  assign or_1720_nl = (COMP_LOOP_acc_7_psp_sva[2:0]!=3'b100) | (~ (STAGE_VEC_LOOP_j_sva_9_0[0]))
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[5])
      | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign or_1718_nl = (operator_64_false_acc_cse_3_sva[3:0]!=4'b1001) | (fsm_output[5])
      | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign mux_1734_nl = MUX_s_1_2_2(or_1720_nl, or_1718_nl, fsm_output[0]);
  assign or_1716_nl = (~ operator_64_false_slc_operator_64_false_acc_1_60_itm) |
      (COMP_LOOP_acc_cse_4_sva[3:0]!=4'b1001) | (~ (fsm_output[0])) | (~ (fsm_output[5]))
      | (fsm_output[6]) | nand_442_cse;
  assign mux_1735_nl = MUX_s_1_2_2(mux_1734_nl, or_1716_nl, fsm_output[4]);
  assign or_1714_nl = (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b01) | (COMP_LOOP_acc_8_psp_sva[1:0]!=2'b10)
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (~
      (fsm_output[5])) | (~ (fsm_output[6])) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign or_1712_nl = (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b01) | (COMP_LOOP_acc_8_psp_sva[1:0]!=2'b10)
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm);
  assign mux_1731_nl = MUX_s_1_2_2(nand_tmp_19, or_tmp_669, or_1712_nl);
  assign nor_321_nl = ~((operator_64_false_acc_cse_4_sva[3:0]!=4'b1001));
  assign mux_1732_nl = MUX_s_1_2_2(or_1714_nl, mux_1731_nl, nor_321_nl);
  assign or_1711_nl = (operator_64_false_acc_cse_5_sva[3:0]!=4'b1001) | (~ (fsm_output[5]))
      | (~ (fsm_output[6])) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign mux_1733_nl = MUX_s_1_2_2(mux_1732_nl, or_1711_nl, fsm_output[0]);
  assign nand_74_nl = ~((fsm_output[4]) & (~ mux_1733_nl));
  assign mux_1736_nl = MUX_s_1_2_2(mux_1735_nl, nand_74_nl, fsm_output[1]);
  assign or_1709_nl = (COMP_LOOP_acc_cse_12_sva[3:0]!=4'b1001) | (~ operator_64_false_slc_operator_64_false_acc_1_60_itm)
      | (~ (fsm_output[0])) | (fsm_output[5]) | (fsm_output[6]) | (fsm_output[3])
      | (~ (fsm_output[2]));
  assign or_1707_nl = (operator_64_false_acc_cse_14_sva[3:0]!=4'b1001) | (fsm_output[0])
      | (~ (fsm_output[5])) | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign mux_1729_nl = MUX_s_1_2_2(or_1709_nl, or_1707_nl, fsm_output[4]);
  assign or_1706_nl = (operator_64_false_acc_cse_12_sva[3:0]!=4'b1001) | (fsm_output[0])
      | (fsm_output[5]) | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign or_1704_nl = (COMP_LOOP_acc_12_psp_sva[1:0]!=2'b10) | (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b01)
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[6:5]!=2'b01)
      | nand_442_cse;
  assign or_1702_nl = (operator_64_false_acc_cse_13_sva[3:0]!=4'b1001) | (fsm_output[6:5]!=2'b01)
      | nand_442_cse;
  assign nor_319_nl = ~((operator_64_false_acc_cse_13_sva[3:0]!=4'b1001));
  assign mux_1725_nl = MUX_s_1_2_2(nand_437_cse, mux_1112_cse, nor_319_nl);
  assign nor_318_nl = ~((COMP_LOOP_acc_cse_14_sva[3:0]!=4'b1001));
  assign mux_1726_nl = MUX_s_1_2_2(or_1702_nl, mux_1725_nl, nor_318_nl);
  assign mux_1727_nl = MUX_s_1_2_2(or_1704_nl, mux_1726_nl, fsm_output[0]);
  assign mux_1728_nl = MUX_s_1_2_2(or_1706_nl, mux_1727_nl, fsm_output[4]);
  assign mux_1730_nl = MUX_s_1_2_2(mux_1729_nl, mux_1728_nl, fsm_output[1]);
  assign mux_1737_nl = MUX_s_1_2_2(mux_1736_nl, mux_1730_nl, fsm_output[9]);
  assign or_1694_nl = (COMP_LOOP_acc_cse_8_sva[3:0]!=4'b1001) | (fsm_output[4]) |
      (~ operator_64_false_slc_operator_64_false_acc_1_60_itm) | (~ (fsm_output[0]))
      | (~ (fsm_output[5])) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign or_1693_nl = (operator_64_false_acc_cse_8_sva[3:0]!=4'b1001) | (fsm_output[0])
      | (~ (fsm_output[5])) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign or_1692_nl = (STAGE_VEC_LOOP_j_sva_9_0[2:0]!=3'b001) | (~ (COMP_LOOP_acc_10_psp_sva[0]))
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[5])
      | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign or_1691_nl = (operator_64_false_acc_cse_9_sva[3:0]!=4'b1001) | (fsm_output[5])
      | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign mux_1720_nl = MUX_s_1_2_2(or_1692_nl, or_1691_nl, fsm_output[0]);
  assign mux_1721_nl = MUX_s_1_2_2(or_1693_nl, mux_1720_nl, fsm_output[4]);
  assign mux_1722_nl = MUX_s_1_2_2(or_1694_nl, mux_1721_nl, fsm_output[1]);
  assign or_1695_nl = (fsm_output[9]) | mux_1722_nl;
  assign mux_1738_nl = MUX_s_1_2_2(mux_1737_nl, or_1695_nl, fsm_output[8]);
  assign mux_1754_nl = MUX_s_1_2_2(mux_1753_nl, mux_1738_nl, fsm_output[7]);
  assign vec_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d = ~ mux_1754_nl;
  assign nor_645_nl = ~((operator_64_false_acc_cse_1_sva[3:0]!=4'b1010) | (fsm_output[2])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]));
  assign nor_646_nl = ~((COMP_LOOP_acc_cse_2_sva[3:0]!=4'b1010) | (fsm_output[2])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]));
  assign mux_1783_nl = MUX_s_1_2_2(nor_645_nl, nor_646_nl, fsm_output[4]);
  assign nor_647_nl = ~((operator_64_false_acc_cse_5_sva[3:0]!=4'b1010) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5])));
  assign nor_648_nl = ~((COMP_LOOP_acc_cse_6_sva[3:0]!=4'b1010) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5])));
  assign mux_1782_nl = MUX_s_1_2_2(nor_647_nl, nor_648_nl, fsm_output[4]);
  assign mux_1784_nl = MUX_s_1_2_2(mux_1783_nl, mux_1782_nl, fsm_output[8]);
  assign nand_78_nl = ~((fsm_output[1]) & mux_1784_nl);
  assign nor_649_nl = ~((operator_64_false_acc_cse_15_sva[3:0]!=4'b1010) | (fsm_output[2])
      | not_tmp_311);
  assign nor_650_nl = ~((COMP_LOOP_acc_cse_sva[3:0]!=4'b1010) | (fsm_output[2]) |
      not_tmp_311);
  assign mux_1780_nl = MUX_s_1_2_2(nor_649_nl, nor_650_nl, fsm_output[4]);
  assign nand_77_nl = ~((fsm_output[8]) & mux_1780_nl);
  assign or_1786_nl = (COMP_LOOP_acc_cse_10_sva[3:0]!=4'b1010) | (fsm_output[2])
      | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign or_1784_nl = (operator_64_false_acc_cse_9_sva[3:0]!=4'b1010) | (fsm_output[2])
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1778_nl = MUX_s_1_2_2(or_1786_nl, or_1784_nl, fsm_output[4]);
  assign or_1783_nl = (fsm_output[4]) | (COMP_LOOP_acc_cse_14_sva[3:0]!=4'b1010)
      | (~ (fsm_output[2])) | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1779_nl = MUX_s_1_2_2(mux_1778_nl, or_1783_nl, fsm_output[8]);
  assign mux_1781_nl = MUX_s_1_2_2(nand_77_nl, mux_1779_nl, fsm_output[1]);
  assign mux_1785_nl = MUX_s_1_2_2(nand_78_nl, mux_1781_nl, fsm_output[9]);
  assign or_1781_nl = (COMP_LOOP_acc_cse_4_sva[3:0]!=4'b1010) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]);
  assign or_1780_nl = (operator_64_false_acc_cse_3_sva[3:0]!=4'b1010) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign mux_1775_nl = MUX_s_1_2_2(or_1781_nl, or_1780_nl, fsm_output[4]);
  assign or_1778_nl = (operator_64_false_acc_cse_7_sva[3:0]!=4'b1010) | (fsm_output[2])
      | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign or_1776_nl = (COMP_LOOP_acc_cse_8_sva[3:0]!=4'b1010) | (fsm_output[2]) |
      (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign mux_1774_nl = MUX_s_1_2_2(or_1778_nl, or_1776_nl, fsm_output[4]);
  assign mux_1776_nl = MUX_s_1_2_2(mux_1775_nl, mux_1774_nl, fsm_output[8]);
  assign or_1782_nl = (fsm_output[1]) | mux_1776_nl;
  assign or_1773_nl = (operator_64_false_acc_cse_11_sva[3:0]!=4'b1010) | (~ (fsm_output[2]))
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign or_1772_nl = (COMP_LOOP_acc_cse_12_sva[3:0]!=4'b1010) | (~ (fsm_output[2]))
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1772_nl = MUX_s_1_2_2(or_1773_nl, or_1772_nl, fsm_output[4]);
  assign or_1774_nl = (fsm_output[8]) | mux_1772_nl;
  assign or_1771_nl = (operator_64_false_acc_cse_13_sva[3:0]!=4'b1010) | (fsm_output[8])
      | (~ (fsm_output[4])) | (~ (fsm_output[2])) | (fsm_output[3]) | not_tmp_312;
  assign mux_1773_nl = MUX_s_1_2_2(or_1774_nl, or_1771_nl, fsm_output[1]);
  assign mux_1777_nl = MUX_s_1_2_2(or_1782_nl, mux_1773_nl, fsm_output[9]);
  assign mux_1786_nl = MUX_s_1_2_2(mux_1785_nl, mux_1777_nl, fsm_output[7]);
  assign or_1769_nl = (~ (fsm_output[8])) | (COMP_LOOP_acc_8_psp_sva[1:0]!=2'b10)
      | (fsm_output[4]) | (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b10) | (~ (fsm_output[2]))
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1768_nl = MUX_s_1_2_2(or_1769_nl, nand_tmp_76, fsm_output[1]);
  assign or_1766_nl = (COMP_LOOP_acc_8_psp_sva[1:0]!=2'b10) | (fsm_output[4]) | (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b10)
      | (~ (fsm_output[2])) | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1766_nl = MUX_s_1_2_2(or_909_cse, or_1766_nl, fsm_output[8]);
  assign mux_1767_nl = MUX_s_1_2_2(mux_1766_nl, nand_tmp_76, fsm_output[1]);
  assign mux_1769_nl = MUX_s_1_2_2(mux_1768_nl, mux_1767_nl, STAGE_VEC_LOOP_j_sva_9_0[3]);
  assign nor_651_nl = ~((operator_64_false_acc_cse_10_sva[3:0]!=4'b1010) | (fsm_output[2])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]));
  assign nor_652_nl = ~((COMP_LOOP_acc_11_psp_sva[2:0]!=3'b101) | (STAGE_VEC_LOOP_j_sva_9_0[0])
      | (fsm_output[2]) | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]));
  assign mux_1763_nl = MUX_s_1_2_2(nor_651_nl, nor_652_nl, fsm_output[4]);
  assign nor_653_nl = ~((operator_64_false_acc_cse_14_sva[3:0]!=4'b1010) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5])));
  assign nor_654_nl = ~((COMP_LOOP_acc_13_psp_sva[2:0]!=3'b101) | (STAGE_VEC_LOOP_j_sva_9_0[0])
      | (~ (fsm_output[2])) | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5])));
  assign mux_1762_nl = MUX_s_1_2_2(nor_653_nl, nor_654_nl, fsm_output[4]);
  assign mux_1764_nl = MUX_s_1_2_2(mux_1763_nl, mux_1762_nl, fsm_output[8]);
  assign nand_75_nl = ~((fsm_output[1]) & mux_1764_nl);
  assign mux_1770_nl = MUX_s_1_2_2(mux_1769_nl, nand_75_nl, fsm_output[9]);
  assign or_1755_nl = (operator_64_false_acc_cse_4_sva[3:0]!=4'b1010) | (fsm_output[4:2]!=3'b101)
      | not_tmp_312;
  assign or_1753_nl = (STAGE_VEC_LOOP_j_sva_9_0[2:0]!=3'b010) | (~ (COMP_LOOP_acc_10_psp_sva[0]))
      | (fsm_output[2]) | not_tmp_311;
  assign or_1751_nl = (operator_64_false_acc_cse_8_sva[3:0]!=4'b1010) | (fsm_output[2])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]);
  assign mux_1758_nl = MUX_s_1_2_2(or_1753_nl, or_1751_nl, fsm_output[4]);
  assign mux_1759_nl = MUX_s_1_2_2(or_1755_nl, mux_1758_nl, fsm_output[8]);
  assign or_1749_nl = (operator_64_false_acc_cse_2_sva[3:0]!=4'b1010) | (fsm_output[2])
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign or_1748_nl = (COMP_LOOP_acc_7_psp_sva[2:0]!=3'b101) | (STAGE_VEC_LOOP_j_sva_9_0[0])
      | (fsm_output[2]) | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1757_nl = MUX_s_1_2_2(or_1749_nl, or_1748_nl, fsm_output[4]);
  assign or_1750_nl = (fsm_output[8]) | mux_1757_nl;
  assign mux_1760_nl = MUX_s_1_2_2(mux_1759_nl, or_1750_nl, fsm_output[1]);
  assign or_1746_nl = (COMP_LOOP_acc_12_psp_sva[1:0]!=2'b10) | (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b10)
      | (~ (fsm_output[2])) | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]);
  assign or_1745_nl = (operator_64_false_acc_cse_12_sva[3:0]!=4'b1010) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign mux_1755_nl = MUX_s_1_2_2(or_1746_nl, or_1745_nl, fsm_output[4]);
  assign or_1743_nl = (fsm_output[4]) | (operator_64_false_acc_cse_sva[3:0]!=4'b1010)
      | (fsm_output[2]) | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign mux_1756_nl = MUX_s_1_2_2(mux_1755_nl, or_1743_nl, fsm_output[8]);
  assign or_1747_nl = (fsm_output[1]) | mux_1756_nl;
  assign mux_1761_nl = MUX_s_1_2_2(mux_1760_nl, or_1747_nl, fsm_output[9]);
  assign mux_1771_nl = MUX_s_1_2_2(mux_1770_nl, mux_1761_nl, fsm_output[7]);
  assign mux_1787_nl = MUX_s_1_2_2(mux_1786_nl, mux_1771_nl, fsm_output[0]);
  assign vec_rsc_0_10_i_wea_d_pff = ~ mux_1787_nl;
  assign or_1850_nl = (operator_64_false_acc_cse_2_sva[3:0]!=4'b1010) | (fsm_output[4])
      | (fsm_output[0]) | (fsm_output[5]) | not_tmp_322;
  assign or_1848_nl = (COMP_LOOP_acc_cse_2_sva[3:0]!=4'b1010) | (~ (fsm_output[0]))
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[5])
      | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign or_1847_nl = (COMP_LOOP_1_operator_64_false_acc_tmp[3:0]!=4'b1010) | (fsm_output[5])
      | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign or_1846_nl = (STAGE_VEC_LOOP_j_sva_9_0[3:0]!=4'b1010) | (fsm_output[5])
      | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign mux_1817_nl = MUX_s_1_2_2(or_1847_nl, or_1846_nl, fsm_output[0]);
  assign mux_1818_nl = MUX_s_1_2_2(or_1848_nl, mux_1817_nl, fsm_output[4]);
  assign mux_1819_nl = MUX_s_1_2_2(or_1850_nl, mux_1818_nl, fsm_output[1]);
  assign or_1845_nl = (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b101) | (STAGE_VEC_LOOP_j_sva_9_0[0])
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[5])
      | not_tmp_322;
  assign or_1843_nl = (operator_64_false_acc_cse_11_sva[3:0]!=4'b1010) | (fsm_output[5])
      | not_tmp_322;
  assign mux_1814_nl = MUX_s_1_2_2(or_1845_nl, or_1843_nl, fsm_output[0]);
  assign or_1841_nl = (fsm_output[0]) | (operator_64_false_acc_cse_10_sva[3:0]!=4'b1010)
      | (fsm_output[5]) | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign mux_1815_nl = MUX_s_1_2_2(mux_1814_nl, or_1841_nl, fsm_output[4]);
  assign or_1839_nl = (~ (fsm_output[4])) | (~ (fsm_output[0])) | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      | (COMP_LOOP_acc_cse_10_sva[3:0]!=4'b1010) | (fsm_output[5]) | (fsm_output[6])
      | (fsm_output[3]) | (fsm_output[2]);
  assign mux_1816_nl = MUX_s_1_2_2(mux_1815_nl, or_1839_nl, fsm_output[1]);
  assign mux_1820_nl = MUX_s_1_2_2(mux_1819_nl, mux_1816_nl, fsm_output[9]);
  assign or_1838_nl = (COMP_LOOP_acc_9_psp_sva[2:0]!=3'b101) | (STAGE_VEC_LOOP_j_sva_9_0[0])
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (~
      (fsm_output[5])) | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign or_1837_nl = (operator_64_false_acc_cse_7_sva[3:0]!=4'b1010) | (~ (fsm_output[5]))
      | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign mux_1810_nl = MUX_s_1_2_2(or_1838_nl, or_1837_nl, fsm_output[0]);
  assign or_1836_nl = (operator_64_false_acc_cse_6_sva[3:0]!=4'b1010) | (fsm_output[0])
      | (~ (fsm_output[5])) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign mux_1811_nl = MUX_s_1_2_2(mux_1810_nl, or_1836_nl, fsm_output[4]);
  assign or_1835_nl = (COMP_LOOP_acc_cse_6_sva[3:0]!=4'b1010) | (fsm_output[4]) |
      (~ (fsm_output[0])) | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      | (fsm_output[6:5]!=2'b01) | nand_442_cse;
  assign mux_1812_nl = MUX_s_1_2_2(mux_1811_nl, or_1835_nl, fsm_output[1]);
  assign nand_300_nl = ~(operator_64_false_slc_operator_64_false_acc_1_60_itm & (fsm_output[0])
      & (COMP_LOOP_acc_cse_sva[3:0]==4'b1010) & (fsm_output[5]) & (fsm_output[6])
      & (fsm_output[3]) & (~ (fsm_output[2])));
  assign or_1832_nl = (COMP_LOOP_acc_13_psp_sva[2:0]!=3'b101) | (STAGE_VEC_LOOP_j_sva_9_0[0])
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (~
      (fsm_output[5])) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign or_1831_nl = (operator_64_false_acc_cse_15_sva[3:0]!=4'b1010) | (~ (fsm_output[5]))
      | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign mux_1807_nl = MUX_s_1_2_2(or_1832_nl, or_1831_nl, fsm_output[0]);
  assign mux_1808_nl = MUX_s_1_2_2(nand_300_nl, mux_1807_nl, fsm_output[4]);
  assign or_1830_nl = (operator_64_false_acc_cse_sva[3:0]!=4'b1010) | (fsm_output[4])
      | (fsm_output[0]) | (~ (fsm_output[5])) | (~ (fsm_output[6])) | (~ (fsm_output[3]))
      | (fsm_output[2]);
  assign mux_1809_nl = MUX_s_1_2_2(mux_1808_nl, or_1830_nl, fsm_output[1]);
  assign mux_1813_nl = MUX_s_1_2_2(mux_1812_nl, mux_1809_nl, fsm_output[9]);
  assign mux_1821_nl = MUX_s_1_2_2(mux_1820_nl, mux_1813_nl, fsm_output[8]);
  assign or_1829_nl = (COMP_LOOP_acc_7_psp_sva[2:0]!=3'b101) | (STAGE_VEC_LOOP_j_sva_9_0[0])
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[5])
      | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign or_1827_nl = (operator_64_false_acc_cse_3_sva[3:0]!=4'b1010) | (fsm_output[5])
      | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign mux_1802_nl = MUX_s_1_2_2(or_1829_nl, or_1827_nl, fsm_output[0]);
  assign or_1825_nl = (~ operator_64_false_slc_operator_64_false_acc_1_60_itm) |
      (COMP_LOOP_acc_cse_4_sva[3:0]!=4'b1010) | (~ (fsm_output[0])) | (~ (fsm_output[5]))
      | (fsm_output[6]) | nand_442_cse;
  assign mux_1803_nl = MUX_s_1_2_2(mux_1802_nl, or_1825_nl, fsm_output[4]);
  assign or_1823_nl = (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b10) | (COMP_LOOP_acc_8_psp_sva[1:0]!=2'b10)
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm);
  assign mux_1799_nl = MUX_s_1_2_2(nand_tmp_19, or_tmp_669, or_1823_nl);
  assign or_1822_nl = (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b10) | (COMP_LOOP_acc_8_psp_sva[1:0]!=2'b10)
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (~
      (fsm_output[5])) | (~ (fsm_output[6])) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign or_1820_nl = (operator_64_false_acc_cse_4_sva[3:0]!=4'b1010);
  assign mux_1800_nl = MUX_s_1_2_2(mux_1799_nl, or_1822_nl, or_1820_nl);
  assign or_1819_nl = (operator_64_false_acc_cse_5_sva[3:0]!=4'b1010) | (~ (fsm_output[5]))
      | (~ (fsm_output[6])) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign mux_1801_nl = MUX_s_1_2_2(mux_1800_nl, or_1819_nl, fsm_output[0]);
  assign nand_80_nl = ~((fsm_output[4]) & (~ mux_1801_nl));
  assign mux_1804_nl = MUX_s_1_2_2(mux_1803_nl, nand_80_nl, fsm_output[1]);
  assign or_1817_nl = (~ operator_64_false_slc_operator_64_false_acc_1_60_itm) |
      (~ (fsm_output[0])) | (COMP_LOOP_acc_cse_12_sva[3:0]!=4'b1010) | (fsm_output[5])
      | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign or_1815_nl = (operator_64_false_acc_cse_14_sva[3:0]!=4'b1010) | (fsm_output[0])
      | (~ (fsm_output[5])) | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign mux_1797_nl = MUX_s_1_2_2(or_1817_nl, or_1815_nl, fsm_output[4]);
  assign or_1814_nl = (operator_64_false_acc_cse_12_sva[3:0]!=4'b1010) | (fsm_output[0])
      | (fsm_output[5]) | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign or_1812_nl = (COMP_LOOP_acc_12_psp_sva[1:0]!=2'b10) | (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b10)
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[6:5]!=2'b01)
      | nand_442_cse;
  assign or_1805_nl = (operator_64_false_acc_cse_13_sva[3:0]!=4'b1010);
  assign mux_1793_nl = MUX_s_1_2_2(mux_1112_cse, nand_437_cse, or_1805_nl);
  assign or_1804_nl = (operator_64_false_acc_cse_13_sva[3:0]!=4'b1010) | (fsm_output[6:5]!=2'b01)
      | nand_442_cse;
  assign or_1802_nl = (COMP_LOOP_acc_cse_14_sva[3:0]!=4'b1010);
  assign mux_1794_nl = MUX_s_1_2_2(mux_1793_nl, or_1804_nl, or_1802_nl);
  assign mux_1795_nl = MUX_s_1_2_2(or_1812_nl, mux_1794_nl, fsm_output[0]);
  assign mux_1796_nl = MUX_s_1_2_2(or_1814_nl, mux_1795_nl, fsm_output[4]);
  assign mux_1798_nl = MUX_s_1_2_2(mux_1797_nl, mux_1796_nl, fsm_output[1]);
  assign mux_1805_nl = MUX_s_1_2_2(mux_1804_nl, mux_1798_nl, fsm_output[9]);
  assign or_1800_nl = (COMP_LOOP_acc_cse_8_sva[3:0]!=4'b1010) | (fsm_output[4]) |
      (~ operator_64_false_slc_operator_64_false_acc_1_60_itm) | (~ (fsm_output[0]))
      | (~ (fsm_output[5])) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign or_1799_nl = (operator_64_false_acc_cse_8_sva[3:0]!=4'b1010) | (fsm_output[0])
      | (~ (fsm_output[5])) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign or_1798_nl = (STAGE_VEC_LOOP_j_sva_9_0[2:0]!=3'b010) | (~ (COMP_LOOP_acc_10_psp_sva[0]))
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[5])
      | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign or_1797_nl = (operator_64_false_acc_cse_9_sva[3:0]!=4'b1010) | (fsm_output[5])
      | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign mux_1788_nl = MUX_s_1_2_2(or_1798_nl, or_1797_nl, fsm_output[0]);
  assign mux_1789_nl = MUX_s_1_2_2(or_1799_nl, mux_1788_nl, fsm_output[4]);
  assign mux_1790_nl = MUX_s_1_2_2(or_1800_nl, mux_1789_nl, fsm_output[1]);
  assign or_1801_nl = (fsm_output[9]) | mux_1790_nl;
  assign mux_1806_nl = MUX_s_1_2_2(mux_1805_nl, or_1801_nl, fsm_output[8]);
  assign mux_1822_nl = MUX_s_1_2_2(mux_1821_nl, mux_1806_nl, fsm_output[7]);
  assign vec_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d = ~ mux_1822_nl;
  assign nor_633_nl = ~((operator_64_false_acc_cse_1_sva[3:0]!=4'b1011) | (fsm_output[2])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]));
  assign nor_634_nl = ~((COMP_LOOP_acc_cse_2_sva[3:0]!=4'b1011) | (fsm_output[2])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]));
  assign mux_1851_nl = MUX_s_1_2_2(nor_633_nl, nor_634_nl, fsm_output[4]);
  assign and_772_nl = (operator_64_false_acc_cse_5_sva[3:0]==4'b1011) & (fsm_output[2])
      & (fsm_output[3]) & (~ (fsm_output[6])) & (fsm_output[5]);
  assign and_778_nl = (COMP_LOOP_acc_cse_6_sva[3:0]==4'b1011) & (fsm_output[2]) &
      (fsm_output[3]) & (~ (fsm_output[6])) & (fsm_output[5]);
  assign mux_1850_nl = MUX_s_1_2_2(and_772_nl, and_778_nl, fsm_output[4]);
  assign mux_1852_nl = MUX_s_1_2_2(mux_1851_nl, mux_1850_nl, fsm_output[8]);
  assign nand_84_nl = ~((fsm_output[1]) & mux_1852_nl);
  assign nor_637_nl = ~((operator_64_false_acc_cse_15_sva[3:0]!=4'b1011) | (fsm_output[2])
      | not_tmp_311);
  assign nor_638_nl = ~((COMP_LOOP_acc_cse_sva[3:0]!=4'b1011) | (fsm_output[2]) |
      not_tmp_311);
  assign mux_1848_nl = MUX_s_1_2_2(nor_637_nl, nor_638_nl, fsm_output[4]);
  assign nand_83_nl = ~((fsm_output[8]) & mux_1848_nl);
  assign or_1895_nl = (COMP_LOOP_acc_cse_10_sva[3:0]!=4'b1011) | (fsm_output[2])
      | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign or_1893_nl = (operator_64_false_acc_cse_9_sva[3:0]!=4'b1011) | (fsm_output[2])
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1846_nl = MUX_s_1_2_2(or_1895_nl, or_1893_nl, fsm_output[4]);
  assign or_1892_nl = (fsm_output[4]) | (COMP_LOOP_acc_cse_14_sva[3:0]!=4'b1011)
      | (~ (fsm_output[2])) | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1847_nl = MUX_s_1_2_2(mux_1846_nl, or_1892_nl, fsm_output[8]);
  assign mux_1849_nl = MUX_s_1_2_2(nand_83_nl, mux_1847_nl, fsm_output[1]);
  assign mux_1853_nl = MUX_s_1_2_2(nand_84_nl, mux_1849_nl, fsm_output[9]);
  assign nand_291_nl = ~((COMP_LOOP_acc_cse_4_sva[3:0]==4'b1011) & (fsm_output[2])
      & (fsm_output[3]) & (fsm_output[6]) & (~ (fsm_output[5])));
  assign nand_471_nl = ~((operator_64_false_acc_cse_3_sva[3:0]==4'b1011) & (fsm_output[2])
      & (fsm_output[3]) & (~ (fsm_output[6])) & (fsm_output[5]));
  assign mux_1843_nl = MUX_s_1_2_2(nand_291_nl, nand_471_nl, fsm_output[4]);
  assign or_1887_nl = (operator_64_false_acc_cse_7_sva[3:0]!=4'b1011) | (fsm_output[2])
      | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign or_1885_nl = (COMP_LOOP_acc_cse_8_sva[3:0]!=4'b1011) | (fsm_output[2]) |
      (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign mux_1842_nl = MUX_s_1_2_2(or_1887_nl, or_1885_nl, fsm_output[4]);
  assign mux_1844_nl = MUX_s_1_2_2(mux_1843_nl, mux_1842_nl, fsm_output[8]);
  assign or_1891_nl = (fsm_output[1]) | mux_1844_nl;
  assign or_1882_nl = (operator_64_false_acc_cse_11_sva[3:0]!=4'b1011) | (~ (fsm_output[2]))
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign or_1881_nl = (COMP_LOOP_acc_cse_12_sva[3:0]!=4'b1011) | (~ (fsm_output[2]))
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1840_nl = MUX_s_1_2_2(or_1882_nl, or_1881_nl, fsm_output[4]);
  assign or_1883_nl = (fsm_output[8]) | mux_1840_nl;
  assign or_1880_nl = (operator_64_false_acc_cse_13_sva[3:0]!=4'b1011) | (fsm_output[8])
      | (~ (fsm_output[4])) | (~ (fsm_output[2])) | (fsm_output[3]) | not_tmp_312;
  assign mux_1841_nl = MUX_s_1_2_2(or_1883_nl, or_1880_nl, fsm_output[1]);
  assign mux_1845_nl = MUX_s_1_2_2(or_1891_nl, mux_1841_nl, fsm_output[9]);
  assign mux_1854_nl = MUX_s_1_2_2(mux_1853_nl, mux_1845_nl, fsm_output[7]);
  assign or_1878_nl = (~ (fsm_output[8])) | (COMP_LOOP_acc_8_psp_sva[1:0]!=2'b10)
      | (fsm_output[4]) | (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b11) | (~ (fsm_output[2]))
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1836_nl = MUX_s_1_2_2(or_1878_nl, nand_tmp_82, fsm_output[1]);
  assign or_1875_nl = (COMP_LOOP_acc_8_psp_sva[1:0]!=2'b10) | (fsm_output[4]) | (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b11)
      | (~ (fsm_output[2])) | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1834_nl = MUX_s_1_2_2(or_1018_cse, or_1875_nl, fsm_output[8]);
  assign mux_1835_nl = MUX_s_1_2_2(mux_1834_nl, nand_tmp_82, fsm_output[1]);
  assign mux_1837_nl = MUX_s_1_2_2(mux_1836_nl, mux_1835_nl, STAGE_VEC_LOOP_j_sva_9_0[3]);
  assign nor_639_nl = ~((operator_64_false_acc_cse_10_sva[3:0]!=4'b1011) | (fsm_output[2])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]));
  assign nor_640_nl = ~((COMP_LOOP_acc_11_psp_sva[2:0]!=3'b101) | (~ (STAGE_VEC_LOOP_j_sva_9_0[0]))
      | (fsm_output[2]) | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]));
  assign mux_1831_nl = MUX_s_1_2_2(nor_639_nl, nor_640_nl, fsm_output[4]);
  assign and_787_nl = (operator_64_false_acc_cse_14_sva[3:0]==4'b1011) & (fsm_output[2])
      & (fsm_output[3]) & (~ (fsm_output[6])) & (fsm_output[5]);
  assign and_788_nl = (COMP_LOOP_acc_13_psp_sva[2:0]==3'b101) & (STAGE_VEC_LOOP_j_sva_9_0[0])
      & (fsm_output[2]) & (fsm_output[3]) & (~ (fsm_output[6])) & (fsm_output[5]);
  assign mux_1830_nl = MUX_s_1_2_2(and_787_nl, and_788_nl, fsm_output[4]);
  assign mux_1832_nl = MUX_s_1_2_2(mux_1831_nl, mux_1830_nl, fsm_output[8]);
  assign nand_81_nl = ~((fsm_output[1]) & mux_1832_nl);
  assign mux_1838_nl = MUX_s_1_2_2(mux_1837_nl, nand_81_nl, fsm_output[9]);
  assign or_1864_nl = (~((operator_64_false_acc_cse_4_sva[3:0]==4'b1011) & (fsm_output[4:2]==3'b101)))
      | not_tmp_312;
  assign or_1862_nl = (STAGE_VEC_LOOP_j_sva_9_0[2:0]!=3'b011) | (~ (COMP_LOOP_acc_10_psp_sva[0]))
      | (fsm_output[2]) | not_tmp_311;
  assign or_1860_nl = (operator_64_false_acc_cse_8_sva[3:0]!=4'b1011) | (fsm_output[2])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]);
  assign mux_1826_nl = MUX_s_1_2_2(or_1862_nl, or_1860_nl, fsm_output[4]);
  assign mux_1827_nl = MUX_s_1_2_2(or_1864_nl, mux_1826_nl, fsm_output[8]);
  assign or_1858_nl = (operator_64_false_acc_cse_2_sva[3:0]!=4'b1011) | (fsm_output[2])
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign or_1857_nl = (COMP_LOOP_acc_7_psp_sva[2:0]!=3'b101) | (~ (STAGE_VEC_LOOP_j_sva_9_0[0]))
      | (fsm_output[2]) | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1825_nl = MUX_s_1_2_2(or_1858_nl, or_1857_nl, fsm_output[4]);
  assign or_1859_nl = (fsm_output[8]) | mux_1825_nl;
  assign mux_1828_nl = MUX_s_1_2_2(mux_1827_nl, or_1859_nl, fsm_output[1]);
  assign nand_296_nl = ~((COMP_LOOP_acc_12_psp_sva[1:0]==2'b10) & (STAGE_VEC_LOOP_j_sva_9_0[1:0]==2'b11)
      & (fsm_output[2]) & (fsm_output[3]) & (fsm_output[6]) & (~ (fsm_output[5])));
  assign nand_452_nl = ~((operator_64_false_acc_cse_12_sva[3:0]==4'b1011) & (fsm_output[2])
      & (fsm_output[3]) & (~ (fsm_output[6])) & (fsm_output[5]));
  assign mux_1823_nl = MUX_s_1_2_2(nand_296_nl, nand_452_nl, fsm_output[4]);
  assign or_1852_nl = (fsm_output[4]) | (operator_64_false_acc_cse_sva[3:0]!=4'b1011)
      | (fsm_output[2]) | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign mux_1824_nl = MUX_s_1_2_2(mux_1823_nl, or_1852_nl, fsm_output[8]);
  assign or_1856_nl = (fsm_output[1]) | mux_1824_nl;
  assign mux_1829_nl = MUX_s_1_2_2(mux_1828_nl, or_1856_nl, fsm_output[9]);
  assign mux_1839_nl = MUX_s_1_2_2(mux_1838_nl, mux_1829_nl, fsm_output[7]);
  assign mux_1855_nl = MUX_s_1_2_2(mux_1854_nl, mux_1839_nl, fsm_output[0]);
  assign vec_rsc_0_11_i_wea_d_pff = ~ mux_1855_nl;
  assign or_1956_nl = (operator_64_false_acc_cse_2_sva[3:0]!=4'b1011) | (fsm_output[4])
      | (fsm_output[0]) | (fsm_output[5]) | not_tmp_322;
  assign nand_277_nl = ~((COMP_LOOP_acc_cse_2_sva[3:0]==4'b1011) & (fsm_output[0])
      & COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm & (~ (fsm_output[5]))
      & (fsm_output[6]) & (fsm_output[3]) & (~ (fsm_output[2])));
  assign or_1953_nl = (COMP_LOOP_1_operator_64_false_acc_tmp[3:0]!=4'b1011) | (fsm_output[5])
      | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign or_1952_nl = (STAGE_VEC_LOOP_j_sva_9_0[3:0]!=4'b1011) | (fsm_output[5])
      | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign mux_1885_nl = MUX_s_1_2_2(or_1953_nl, or_1952_nl, fsm_output[0]);
  assign mux_1886_nl = MUX_s_1_2_2(nand_277_nl, mux_1885_nl, fsm_output[4]);
  assign mux_1887_nl = MUX_s_1_2_2(or_1956_nl, mux_1886_nl, fsm_output[1]);
  assign or_1951_nl = (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b101) | (~ (STAGE_VEC_LOOP_j_sva_9_0[0]))
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[5])
      | not_tmp_322;
  assign or_1949_nl = (operator_64_false_acc_cse_11_sva[3:0]!=4'b1011) | (fsm_output[5])
      | not_tmp_322;
  assign mux_1882_nl = MUX_s_1_2_2(or_1951_nl, or_1949_nl, fsm_output[0]);
  assign or_1947_nl = (fsm_output[0]) | (operator_64_false_acc_cse_10_sva[3:0]!=4'b1011)
      | (fsm_output[5]) | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign mux_1883_nl = MUX_s_1_2_2(mux_1882_nl, or_1947_nl, fsm_output[4]);
  assign or_1945_nl = (COMP_LOOP_acc_cse_10_sva[3:0]!=4'b1011) | (~ (fsm_output[4]))
      | (~ (fsm_output[0])) | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      | (fsm_output[5]) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign mux_1884_nl = MUX_s_1_2_2(mux_1883_nl, or_1945_nl, fsm_output[1]);
  assign mux_1888_nl = MUX_s_1_2_2(mux_1887_nl, mux_1884_nl, fsm_output[9]);
  assign nand_278_nl = ~((COMP_LOOP_acc_9_psp_sva[2:0]==3'b101) & (STAGE_VEC_LOOP_j_sva_9_0[0])
      & COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm & (fsm_output[5])
      & (fsm_output[6]) & (fsm_output[3]) & (~ (fsm_output[2])));
  assign nand_279_nl = ~((operator_64_false_acc_cse_7_sva[3:0]==4'b1011) & (fsm_output[5])
      & (fsm_output[6]) & (fsm_output[3]) & (~ (fsm_output[2])));
  assign mux_1878_nl = MUX_s_1_2_2(nand_278_nl, nand_279_nl, fsm_output[0]);
  assign or_1942_nl = (operator_64_false_acc_cse_6_sva[3:0]!=4'b1011) | (fsm_output[0])
      | (~ (fsm_output[5])) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign mux_1879_nl = MUX_s_1_2_2(mux_1878_nl, or_1942_nl, fsm_output[4]);
  assign or_1941_nl = (COMP_LOOP_acc_cse_6_sva[3:0]!=4'b1011) | (fsm_output[4]) |
      (~ (fsm_output[0])) | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      | (fsm_output[6:5]!=2'b01) | nand_442_cse;
  assign mux_1880_nl = MUX_s_1_2_2(mux_1879_nl, or_1941_nl, fsm_output[1]);
  assign nand_280_nl = ~(operator_64_false_slc_operator_64_false_acc_1_60_itm & (fsm_output[0])
      & (COMP_LOOP_acc_cse_sva[3:0]==4'b1011) & (fsm_output[5]) & (fsm_output[6])
      & (fsm_output[3]) & (~ (fsm_output[2])));
  assign or_1938_nl = (COMP_LOOP_acc_13_psp_sva[2:0]!=3'b101) | (~ (STAGE_VEC_LOOP_j_sva_9_0[0]))
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (~
      (fsm_output[5])) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign or_1937_nl = (operator_64_false_acc_cse_15_sva[3:0]!=4'b1011) | (~ (fsm_output[5]))
      | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign mux_1875_nl = MUX_s_1_2_2(or_1938_nl, or_1937_nl, fsm_output[0]);
  assign mux_1876_nl = MUX_s_1_2_2(nand_280_nl, mux_1875_nl, fsm_output[4]);
  assign or_1936_nl = (operator_64_false_acc_cse_sva[3:0]!=4'b1011) | (fsm_output[4])
      | (fsm_output[0]) | (~ (fsm_output[5])) | (~ (fsm_output[6])) | (~ (fsm_output[3]))
      | (fsm_output[2]);
  assign mux_1877_nl = MUX_s_1_2_2(mux_1876_nl, or_1936_nl, fsm_output[1]);
  assign mux_1881_nl = MUX_s_1_2_2(mux_1880_nl, mux_1877_nl, fsm_output[9]);
  assign mux_1889_nl = MUX_s_1_2_2(mux_1888_nl, mux_1881_nl, fsm_output[8]);
  assign or_1935_nl = (COMP_LOOP_acc_7_psp_sva[2:0]!=3'b101) | (~ (STAGE_VEC_LOOP_j_sva_9_0[0]))
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[5])
      | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign or_1933_nl = (operator_64_false_acc_cse_3_sva[3:0]!=4'b1011) | (fsm_output[5])
      | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign mux_1870_nl = MUX_s_1_2_2(or_1935_nl, or_1933_nl, fsm_output[0]);
  assign or_1931_nl = (~(operator_64_false_slc_operator_64_false_acc_1_60_itm & (COMP_LOOP_acc_cse_4_sva[3:0]==4'b1011)
      & (fsm_output[0]) & (fsm_output[5]) & (~ (fsm_output[6])))) | nand_442_cse;
  assign mux_1871_nl = MUX_s_1_2_2(mux_1870_nl, or_1931_nl, fsm_output[4]);
  assign nand_466_nl = ~((STAGE_VEC_LOOP_j_sva_9_0[1:0]==2'b11) & (COMP_LOOP_acc_8_psp_sva[1:0]==2'b10)
      & COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm & (fsm_output[5])
      & (fsm_output[6]) & (~ (fsm_output[3])) & (fsm_output[2]));
  assign nand_283_nl = ~((STAGE_VEC_LOOP_j_sva_9_0[1:0]==2'b11) & (COMP_LOOP_acc_8_psp_sva[1:0]==2'b10)
      & COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm);
  assign mux_1867_nl = MUX_s_1_2_2(nand_tmp_19, or_tmp_669, nand_283_nl);
  assign and_543_nl = (operator_64_false_acc_cse_4_sva[3:0]==4'b1011);
  assign mux_1868_nl = MUX_s_1_2_2(nand_466_nl, mux_1867_nl, and_543_nl);
  assign nand_462_nl = ~((operator_64_false_acc_cse_5_sva[3:0]==4'b1011) & (fsm_output[5])
      & (fsm_output[6]) & (~ (fsm_output[3])) & (fsm_output[2]));
  assign mux_1869_nl = MUX_s_1_2_2(mux_1868_nl, nand_462_nl, fsm_output[0]);
  assign nand_86_nl = ~((fsm_output[4]) & (~ mux_1869_nl));
  assign mux_1872_nl = MUX_s_1_2_2(mux_1871_nl, nand_86_nl, fsm_output[1]);
  assign or_1924_nl = (~ operator_64_false_slc_operator_64_false_acc_1_60_itm) |
      (~ (fsm_output[0])) | (COMP_LOOP_acc_cse_12_sva[3:0]!=4'b1011) | (fsm_output[5])
      | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign or_1922_nl = (operator_64_false_acc_cse_14_sva[3:0]!=4'b1011) | (fsm_output[0])
      | (~ (fsm_output[5])) | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign mux_1865_nl = MUX_s_1_2_2(or_1924_nl, or_1922_nl, fsm_output[4]);
  assign or_1921_nl = (operator_64_false_acc_cse_12_sva[3:0]!=4'b1011) | (fsm_output[0])
      | (fsm_output[5]) | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign or_1919_nl = (~((COMP_LOOP_acc_12_psp_sva[1:0]==2'b10) & (STAGE_VEC_LOOP_j_sva_9_0[1:0]==2'b11)
      & COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm & (fsm_output[6:5]==2'b01)))
      | nand_442_cse;
  assign or_1917_nl = (operator_64_false_acc_cse_13_sva[3:0]!=4'b1011) | (fsm_output[6:5]!=2'b01)
      | nand_442_cse;
  assign and_544_nl = (operator_64_false_acc_cse_13_sva[3:0]==4'b1011);
  assign mux_1861_nl = MUX_s_1_2_2(nand_437_cse, mux_1112_cse, and_544_nl);
  assign and_545_nl = (COMP_LOOP_acc_cse_14_sva[3:0]==4'b1011);
  assign mux_1862_nl = MUX_s_1_2_2(or_1917_nl, mux_1861_nl, and_545_nl);
  assign mux_1863_nl = MUX_s_1_2_2(or_1919_nl, mux_1862_nl, fsm_output[0]);
  assign mux_1864_nl = MUX_s_1_2_2(or_1921_nl, mux_1863_nl, fsm_output[4]);
  assign mux_1866_nl = MUX_s_1_2_2(mux_1865_nl, mux_1864_nl, fsm_output[1]);
  assign mux_1873_nl = MUX_s_1_2_2(mux_1872_nl, mux_1866_nl, fsm_output[9]);
  assign or_1909_nl = (COMP_LOOP_acc_cse_8_sva[3:0]!=4'b1011) | (fsm_output[4]) |
      (~ operator_64_false_slc_operator_64_false_acc_1_60_itm) | (~ (fsm_output[0]))
      | (~ (fsm_output[5])) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign or_1908_nl = (operator_64_false_acc_cse_8_sva[3:0]!=4'b1011) | (fsm_output[0])
      | (~ (fsm_output[5])) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign or_1907_nl = (STAGE_VEC_LOOP_j_sva_9_0[2:0]!=3'b011) | (~ (COMP_LOOP_acc_10_psp_sva[0]))
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[5])
      | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign or_1906_nl = (operator_64_false_acc_cse_9_sva[3:0]!=4'b1011) | (fsm_output[5])
      | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign mux_1856_nl = MUX_s_1_2_2(or_1907_nl, or_1906_nl, fsm_output[0]);
  assign mux_1857_nl = MUX_s_1_2_2(or_1908_nl, mux_1856_nl, fsm_output[4]);
  assign mux_1858_nl = MUX_s_1_2_2(or_1909_nl, mux_1857_nl, fsm_output[1]);
  assign or_1910_nl = (fsm_output[9]) | mux_1858_nl;
  assign mux_1874_nl = MUX_s_1_2_2(mux_1873_nl, or_1910_nl, fsm_output[8]);
  assign mux_1890_nl = MUX_s_1_2_2(mux_1889_nl, mux_1874_nl, fsm_output[7]);
  assign vec_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d = ~ mux_1890_nl;
  assign nor_621_nl = ~((operator_64_false_acc_cse_1_sva[3:0]!=4'b1100) | (fsm_output[2])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]));
  assign nor_622_nl = ~((COMP_LOOP_acc_cse_2_sva[3:0]!=4'b1100) | (fsm_output[2])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]));
  assign mux_1919_nl = MUX_s_1_2_2(nor_621_nl, nor_622_nl, fsm_output[4]);
  assign nor_623_nl = ~((operator_64_false_acc_cse_5_sva[3:0]!=4'b1100) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5])));
  assign nor_624_nl = ~((COMP_LOOP_acc_cse_6_sva[3:0]!=4'b1100) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5])));
  assign mux_1918_nl = MUX_s_1_2_2(nor_623_nl, nor_624_nl, fsm_output[4]);
  assign mux_1920_nl = MUX_s_1_2_2(mux_1919_nl, mux_1918_nl, fsm_output[8]);
  assign nand_90_nl = ~((fsm_output[1]) & mux_1920_nl);
  assign nor_625_nl = ~((operator_64_false_acc_cse_15_sva[3:0]!=4'b1100) | (fsm_output[2])
      | not_tmp_311);
  assign nor_626_nl = ~((COMP_LOOP_acc_cse_sva[3:0]!=4'b1100) | (fsm_output[2]) |
      not_tmp_311);
  assign mux_1916_nl = MUX_s_1_2_2(nor_625_nl, nor_626_nl, fsm_output[4]);
  assign nand_89_nl = ~((fsm_output[8]) & mux_1916_nl);
  assign or_2001_nl = (COMP_LOOP_acc_cse_10_sva[3:0]!=4'b1100) | (fsm_output[2])
      | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign or_1999_nl = (operator_64_false_acc_cse_9_sva[3:0]!=4'b1100) | (fsm_output[2])
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1914_nl = MUX_s_1_2_2(or_2001_nl, or_1999_nl, fsm_output[4]);
  assign or_1998_nl = (fsm_output[4]) | (COMP_LOOP_acc_cse_14_sva[3:0]!=4'b1100)
      | (~ (fsm_output[2])) | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1915_nl = MUX_s_1_2_2(mux_1914_nl, or_1998_nl, fsm_output[8]);
  assign mux_1917_nl = MUX_s_1_2_2(nand_89_nl, mux_1915_nl, fsm_output[1]);
  assign mux_1921_nl = MUX_s_1_2_2(nand_90_nl, mux_1917_nl, fsm_output[9]);
  assign or_1996_nl = (COMP_LOOP_acc_cse_4_sva[3:0]!=4'b1100) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]);
  assign or_1995_nl = (operator_64_false_acc_cse_3_sva[3:0]!=4'b1100) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign mux_1911_nl = MUX_s_1_2_2(or_1996_nl, or_1995_nl, fsm_output[4]);
  assign or_1993_nl = (operator_64_false_acc_cse_7_sva[3:0]!=4'b1100) | (fsm_output[2])
      | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign or_1991_nl = (COMP_LOOP_acc_cse_8_sva[3:0]!=4'b1100) | (fsm_output[2]) |
      (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign mux_1910_nl = MUX_s_1_2_2(or_1993_nl, or_1991_nl, fsm_output[4]);
  assign mux_1912_nl = MUX_s_1_2_2(mux_1911_nl, mux_1910_nl, fsm_output[8]);
  assign or_1997_nl = (fsm_output[1]) | mux_1912_nl;
  assign or_1988_nl = (operator_64_false_acc_cse_11_sva[3:0]!=4'b1100) | (~ (fsm_output[2]))
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign or_1987_nl = (COMP_LOOP_acc_cse_12_sva[3:0]!=4'b1100) | (~ (fsm_output[2]))
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1908_nl = MUX_s_1_2_2(or_1988_nl, or_1987_nl, fsm_output[4]);
  assign or_1989_nl = (fsm_output[8]) | mux_1908_nl;
  assign or_1986_nl = (operator_64_false_acc_cse_13_sva[3:0]!=4'b1100) | (fsm_output[8])
      | (~ (fsm_output[4])) | (~ (fsm_output[2])) | (fsm_output[3]) | not_tmp_312;
  assign mux_1909_nl = MUX_s_1_2_2(or_1989_nl, or_1986_nl, fsm_output[1]);
  assign mux_1913_nl = MUX_s_1_2_2(or_1997_nl, mux_1909_nl, fsm_output[9]);
  assign mux_1922_nl = MUX_s_1_2_2(mux_1921_nl, mux_1913_nl, fsm_output[7]);
  assign or_1984_nl = (~ (fsm_output[8])) | (COMP_LOOP_acc_8_psp_sva[1:0]!=2'b11)
      | (fsm_output[4]) | (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b00) | (~ (fsm_output[2]))
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1904_nl = MUX_s_1_2_2(or_1984_nl, nand_tmp_88, fsm_output[1]);
  assign or_1981_nl = (COMP_LOOP_acc_8_psp_sva[1:0]!=2'b11) | (fsm_output[4]) | (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b00)
      | (~ (fsm_output[2])) | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1902_nl = MUX_s_1_2_2(or_1124_cse, or_1981_nl, fsm_output[8]);
  assign mux_1903_nl = MUX_s_1_2_2(mux_1902_nl, nand_tmp_88, fsm_output[1]);
  assign mux_1905_nl = MUX_s_1_2_2(mux_1904_nl, mux_1903_nl, STAGE_VEC_LOOP_j_sva_9_0[3]);
  assign nor_627_nl = ~((operator_64_false_acc_cse_10_sva[3:0]!=4'b1100) | (fsm_output[2])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]));
  assign nor_628_nl = ~((COMP_LOOP_acc_11_psp_sva[2:0]!=3'b110) | (STAGE_VEC_LOOP_j_sva_9_0[0])
      | (fsm_output[2]) | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]));
  assign mux_1899_nl = MUX_s_1_2_2(nor_627_nl, nor_628_nl, fsm_output[4]);
  assign nor_629_nl = ~((operator_64_false_acc_cse_14_sva[3:0]!=4'b1100) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5])));
  assign nor_630_nl = ~((COMP_LOOP_acc_13_psp_sva[2:0]!=3'b110) | (STAGE_VEC_LOOP_j_sva_9_0[0])
      | (~ (fsm_output[2])) | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5])));
  assign mux_1898_nl = MUX_s_1_2_2(nor_629_nl, nor_630_nl, fsm_output[4]);
  assign mux_1900_nl = MUX_s_1_2_2(mux_1899_nl, mux_1898_nl, fsm_output[8]);
  assign nand_87_nl = ~((fsm_output[1]) & mux_1900_nl);
  assign mux_1906_nl = MUX_s_1_2_2(mux_1905_nl, nand_87_nl, fsm_output[9]);
  assign or_1970_nl = (operator_64_false_acc_cse_4_sva[3:0]!=4'b1100) | (fsm_output[4:2]!=3'b101)
      | not_tmp_312;
  assign or_1968_nl = (STAGE_VEC_LOOP_j_sva_9_0[2:0]!=3'b100) | (~ (COMP_LOOP_acc_10_psp_sva[0]))
      | (fsm_output[2]) | not_tmp_311;
  assign or_1966_nl = (operator_64_false_acc_cse_8_sva[3:0]!=4'b1100) | (fsm_output[2])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]);
  assign mux_1894_nl = MUX_s_1_2_2(or_1968_nl, or_1966_nl, fsm_output[4]);
  assign mux_1895_nl = MUX_s_1_2_2(or_1970_nl, mux_1894_nl, fsm_output[8]);
  assign or_1964_nl = (operator_64_false_acc_cse_2_sva[3:0]!=4'b1100) | (fsm_output[2])
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign or_1963_nl = (COMP_LOOP_acc_7_psp_sva[2:0]!=3'b110) | (STAGE_VEC_LOOP_j_sva_9_0[0])
      | (fsm_output[2]) | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1893_nl = MUX_s_1_2_2(or_1964_nl, or_1963_nl, fsm_output[4]);
  assign or_1965_nl = (fsm_output[8]) | mux_1893_nl;
  assign mux_1896_nl = MUX_s_1_2_2(mux_1895_nl, or_1965_nl, fsm_output[1]);
  assign or_1961_nl = (COMP_LOOP_acc_12_psp_sva[1:0]!=2'b11) | (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b00)
      | (~ (fsm_output[2])) | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]);
  assign or_1960_nl = (operator_64_false_acc_cse_12_sva[3:0]!=4'b1100) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign mux_1891_nl = MUX_s_1_2_2(or_1961_nl, or_1960_nl, fsm_output[4]);
  assign or_1958_nl = (fsm_output[4]) | (operator_64_false_acc_cse_sva[3:0]!=4'b1100)
      | (fsm_output[2]) | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign mux_1892_nl = MUX_s_1_2_2(mux_1891_nl, or_1958_nl, fsm_output[8]);
  assign or_1962_nl = (fsm_output[1]) | mux_1892_nl;
  assign mux_1897_nl = MUX_s_1_2_2(mux_1896_nl, or_1962_nl, fsm_output[9]);
  assign mux_1907_nl = MUX_s_1_2_2(mux_1906_nl, mux_1897_nl, fsm_output[7]);
  assign mux_1923_nl = MUX_s_1_2_2(mux_1922_nl, mux_1907_nl, fsm_output[0]);
  assign vec_rsc_0_12_i_wea_d_pff = ~ mux_1923_nl;
  assign or_2065_nl = (operator_64_false_acc_cse_2_sva[3:0]!=4'b1100) | (fsm_output[4])
      | (fsm_output[0]) | (fsm_output[5]) | not_tmp_322;
  assign or_2063_nl = (COMP_LOOP_acc_cse_2_sva[3:0]!=4'b1100) | (~ (fsm_output[0]))
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[5])
      | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign or_2062_nl = (COMP_LOOP_1_operator_64_false_acc_tmp[3:0]!=4'b1100) | (fsm_output[5])
      | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign or_2061_nl = (STAGE_VEC_LOOP_j_sva_9_0[3:0]!=4'b1100) | (fsm_output[5])
      | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign mux_1953_nl = MUX_s_1_2_2(or_2062_nl, or_2061_nl, fsm_output[0]);
  assign mux_1954_nl = MUX_s_1_2_2(or_2063_nl, mux_1953_nl, fsm_output[4]);
  assign mux_1955_nl = MUX_s_1_2_2(or_2065_nl, mux_1954_nl, fsm_output[1]);
  assign or_2060_nl = (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b110) | (STAGE_VEC_LOOP_j_sva_9_0[0])
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[5])
      | not_tmp_322;
  assign or_2058_nl = (operator_64_false_acc_cse_11_sva[3:0]!=4'b1100) | (fsm_output[5])
      | not_tmp_322;
  assign mux_1950_nl = MUX_s_1_2_2(or_2060_nl, or_2058_nl, fsm_output[0]);
  assign or_2056_nl = (fsm_output[0]) | (operator_64_false_acc_cse_10_sva[3:0]!=4'b1100)
      | (fsm_output[5]) | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign mux_1951_nl = MUX_s_1_2_2(mux_1950_nl, or_2056_nl, fsm_output[4]);
  assign or_2054_nl = (~ (fsm_output[4])) | (~ (fsm_output[0])) | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      | (COMP_LOOP_acc_cse_10_sva[3:0]!=4'b1100) | (fsm_output[5]) | (fsm_output[6])
      | (fsm_output[3]) | (fsm_output[2]);
  assign mux_1952_nl = MUX_s_1_2_2(mux_1951_nl, or_2054_nl, fsm_output[1]);
  assign mux_1956_nl = MUX_s_1_2_2(mux_1955_nl, mux_1952_nl, fsm_output[9]);
  assign or_2053_nl = (COMP_LOOP_acc_9_psp_sva[2:0]!=3'b110) | (STAGE_VEC_LOOP_j_sva_9_0[0])
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (~
      (fsm_output[5])) | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign or_2052_nl = (operator_64_false_acc_cse_7_sva[3:0]!=4'b1100) | (~ (fsm_output[5]))
      | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign mux_1946_nl = MUX_s_1_2_2(or_2053_nl, or_2052_nl, fsm_output[0]);
  assign or_2051_nl = (operator_64_false_acc_cse_6_sva[3:0]!=4'b1100) | (fsm_output[0])
      | (~ (fsm_output[5])) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign mux_1947_nl = MUX_s_1_2_2(mux_1946_nl, or_2051_nl, fsm_output[4]);
  assign or_2050_nl = (COMP_LOOP_acc_cse_6_sva[3:0]!=4'b1100) | (fsm_output[4]) |
      (~ (fsm_output[0])) | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      | (fsm_output[6:5]!=2'b01) | nand_442_cse;
  assign mux_1948_nl = MUX_s_1_2_2(mux_1947_nl, or_2050_nl, fsm_output[1]);
  assign nand_271_nl = ~((COMP_LOOP_acc_cse_sva[3:0]==4'b1100) & operator_64_false_slc_operator_64_false_acc_1_60_itm
      & (fsm_output[0]) & (fsm_output[5]) & (fsm_output[6]) & (fsm_output[3]) & (~
      (fsm_output[2])));
  assign or_2047_nl = (COMP_LOOP_acc_13_psp_sva[2:0]!=3'b110) | (STAGE_VEC_LOOP_j_sva_9_0[0])
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (~
      (fsm_output[5])) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign or_2046_nl = (operator_64_false_acc_cse_15_sva[3:0]!=4'b1100) | (~ (fsm_output[5]))
      | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign mux_1943_nl = MUX_s_1_2_2(or_2047_nl, or_2046_nl, fsm_output[0]);
  assign mux_1944_nl = MUX_s_1_2_2(nand_271_nl, mux_1943_nl, fsm_output[4]);
  assign or_2045_nl = (operator_64_false_acc_cse_sva[3:0]!=4'b1100) | (fsm_output[4])
      | (fsm_output[0]) | (~ (fsm_output[5])) | (~ (fsm_output[6])) | (~ (fsm_output[3]))
      | (fsm_output[2]);
  assign mux_1945_nl = MUX_s_1_2_2(mux_1944_nl, or_2045_nl, fsm_output[1]);
  assign mux_1949_nl = MUX_s_1_2_2(mux_1948_nl, mux_1945_nl, fsm_output[9]);
  assign mux_1957_nl = MUX_s_1_2_2(mux_1956_nl, mux_1949_nl, fsm_output[8]);
  assign or_2044_nl = (COMP_LOOP_acc_7_psp_sva[2:0]!=3'b110) | (STAGE_VEC_LOOP_j_sva_9_0[0])
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[5])
      | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign or_2042_nl = (operator_64_false_acc_cse_3_sva[3:0]!=4'b1100) | (fsm_output[5])
      | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign mux_1938_nl = MUX_s_1_2_2(or_2044_nl, or_2042_nl, fsm_output[0]);
  assign or_2040_nl = (~ operator_64_false_slc_operator_64_false_acc_1_60_itm) |
      (COMP_LOOP_acc_cse_4_sva[3:0]!=4'b1100) | (~ (fsm_output[0])) | (~ (fsm_output[5]))
      | (fsm_output[6]) | nand_442_cse;
  assign mux_1939_nl = MUX_s_1_2_2(mux_1938_nl, or_2040_nl, fsm_output[4]);
  assign or_2038_nl = (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b00) | (COMP_LOOP_acc_8_psp_sva[1:0]!=2'b11)
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm);
  assign mux_1935_nl = MUX_s_1_2_2(nand_tmp_19, or_tmp_669, or_2038_nl);
  assign or_2037_nl = (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b00) | (COMP_LOOP_acc_8_psp_sva[1:0]!=2'b11)
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (~
      (fsm_output[5])) | (~ (fsm_output[6])) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign or_2035_nl = (operator_64_false_acc_cse_4_sva[3:0]!=4'b1100);
  assign mux_1936_nl = MUX_s_1_2_2(mux_1935_nl, or_2037_nl, or_2035_nl);
  assign or_2034_nl = (operator_64_false_acc_cse_5_sva[3:0]!=4'b1100) | (~ (fsm_output[5]))
      | (~ (fsm_output[6])) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign mux_1937_nl = MUX_s_1_2_2(mux_1936_nl, or_2034_nl, fsm_output[0]);
  assign nand_92_nl = ~((fsm_output[4]) & (~ mux_1937_nl));
  assign mux_1940_nl = MUX_s_1_2_2(mux_1939_nl, nand_92_nl, fsm_output[1]);
  assign or_2032_nl = (COMP_LOOP_acc_cse_12_sva[3:0]!=4'b1100) | (~ operator_64_false_slc_operator_64_false_acc_1_60_itm)
      | (~ (fsm_output[0])) | (fsm_output[5]) | (fsm_output[6]) | (fsm_output[3])
      | (~ (fsm_output[2]));
  assign or_2030_nl = (operator_64_false_acc_cse_14_sva[3:0]!=4'b1100) | (fsm_output[0])
      | (~ (fsm_output[5])) | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign mux_1933_nl = MUX_s_1_2_2(or_2032_nl, or_2030_nl, fsm_output[4]);
  assign or_2029_nl = (operator_64_false_acc_cse_12_sva[3:0]!=4'b1100) | (fsm_output[0])
      | (fsm_output[5]) | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign or_2027_nl = (COMP_LOOP_acc_12_psp_sva[1:0]!=2'b11) | (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b00)
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[6:5]!=2'b01)
      | nand_442_cse;
  assign or_2020_nl = (operator_64_false_acc_cse_13_sva[3:0]!=4'b1100);
  assign mux_1929_nl = MUX_s_1_2_2(mux_1112_cse, nand_437_cse, or_2020_nl);
  assign or_2019_nl = (operator_64_false_acc_cse_13_sva[3:0]!=4'b1100) | (fsm_output[6:5]!=2'b01)
      | nand_442_cse;
  assign or_2017_nl = (COMP_LOOP_acc_cse_14_sva[3:0]!=4'b1100);
  assign mux_1930_nl = MUX_s_1_2_2(mux_1929_nl, or_2019_nl, or_2017_nl);
  assign mux_1931_nl = MUX_s_1_2_2(or_2027_nl, mux_1930_nl, fsm_output[0]);
  assign mux_1932_nl = MUX_s_1_2_2(or_2029_nl, mux_1931_nl, fsm_output[4]);
  assign mux_1934_nl = MUX_s_1_2_2(mux_1933_nl, mux_1932_nl, fsm_output[1]);
  assign mux_1941_nl = MUX_s_1_2_2(mux_1940_nl, mux_1934_nl, fsm_output[9]);
  assign or_2015_nl = (COMP_LOOP_acc_cse_8_sva[3:0]!=4'b1100) | (fsm_output[4]) |
      (~ operator_64_false_slc_operator_64_false_acc_1_60_itm) | (~ (fsm_output[0]))
      | (~ (fsm_output[5])) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign or_2014_nl = (operator_64_false_acc_cse_8_sva[3:0]!=4'b1100) | (fsm_output[0])
      | (~ (fsm_output[5])) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign or_2013_nl = (STAGE_VEC_LOOP_j_sva_9_0[2:0]!=3'b100) | (~ (COMP_LOOP_acc_10_psp_sva[0]))
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[5])
      | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign or_2012_nl = (operator_64_false_acc_cse_9_sva[3:0]!=4'b1100) | (fsm_output[5])
      | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign mux_1924_nl = MUX_s_1_2_2(or_2013_nl, or_2012_nl, fsm_output[0]);
  assign mux_1925_nl = MUX_s_1_2_2(or_2014_nl, mux_1924_nl, fsm_output[4]);
  assign mux_1926_nl = MUX_s_1_2_2(or_2015_nl, mux_1925_nl, fsm_output[1]);
  assign or_2016_nl = (fsm_output[9]) | mux_1926_nl;
  assign mux_1942_nl = MUX_s_1_2_2(mux_1941_nl, or_2016_nl, fsm_output[8]);
  assign mux_1958_nl = MUX_s_1_2_2(mux_1957_nl, mux_1942_nl, fsm_output[7]);
  assign vec_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d = ~ mux_1958_nl;
  assign nor_609_nl = ~((operator_64_false_acc_cse_1_sva[3:0]!=4'b1101) | (fsm_output[2])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]));
  assign nor_610_nl = ~((COMP_LOOP_acc_cse_2_sva[3:0]!=4'b1101) | (fsm_output[2])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]));
  assign mux_1987_nl = MUX_s_1_2_2(nor_609_nl, nor_610_nl, fsm_output[4]);
  assign and_771_nl = (operator_64_false_acc_cse_5_sva[3:0]==4'b1101) & (fsm_output[2])
      & (fsm_output[3]) & (~ (fsm_output[6])) & (fsm_output[5]);
  assign and_777_nl = (COMP_LOOP_acc_cse_6_sva[3:0]==4'b1101) & (fsm_output[2]) &
      (fsm_output[3]) & (~ (fsm_output[6])) & (fsm_output[5]);
  assign mux_1986_nl = MUX_s_1_2_2(and_771_nl, and_777_nl, fsm_output[4]);
  assign mux_1988_nl = MUX_s_1_2_2(mux_1987_nl, mux_1986_nl, fsm_output[8]);
  assign nand_96_nl = ~((fsm_output[1]) & mux_1988_nl);
  assign nor_613_nl = ~((operator_64_false_acc_cse_15_sva[3:0]!=4'b1101) | (fsm_output[2])
      | not_tmp_311);
  assign nor_614_nl = ~((COMP_LOOP_acc_cse_sva[3:0]!=4'b1101) | (fsm_output[2]) |
      not_tmp_311);
  assign mux_1984_nl = MUX_s_1_2_2(nor_613_nl, nor_614_nl, fsm_output[4]);
  assign nand_95_nl = ~((fsm_output[8]) & mux_1984_nl);
  assign or_2110_nl = (COMP_LOOP_acc_cse_10_sva[3:0]!=4'b1101) | (fsm_output[2])
      | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign or_2108_nl = (operator_64_false_acc_cse_9_sva[3:0]!=4'b1101) | (fsm_output[2])
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1982_nl = MUX_s_1_2_2(or_2110_nl, or_2108_nl, fsm_output[4]);
  assign or_2107_nl = (fsm_output[4]) | (COMP_LOOP_acc_cse_14_sva[3:0]!=4'b1101)
      | (~ (fsm_output[2])) | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1983_nl = MUX_s_1_2_2(mux_1982_nl, or_2107_nl, fsm_output[8]);
  assign mux_1985_nl = MUX_s_1_2_2(nand_95_nl, mux_1983_nl, fsm_output[1]);
  assign mux_1989_nl = MUX_s_1_2_2(nand_96_nl, mux_1985_nl, fsm_output[9]);
  assign nand_262_nl = ~((COMP_LOOP_acc_cse_4_sva[3:0]==4'b1101) & (fsm_output[2])
      & (fsm_output[3]) & (fsm_output[6]) & (~ (fsm_output[5])));
  assign nand_470_nl = ~((operator_64_false_acc_cse_3_sva[3:0]==4'b1101) & (fsm_output[2])
      & (fsm_output[3]) & (~ (fsm_output[6])) & (fsm_output[5]));
  assign mux_1979_nl = MUX_s_1_2_2(nand_262_nl, nand_470_nl, fsm_output[4]);
  assign or_2102_nl = (operator_64_false_acc_cse_7_sva[3:0]!=4'b1101) | (fsm_output[2])
      | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign or_2100_nl = (COMP_LOOP_acc_cse_8_sva[3:0]!=4'b1101) | (fsm_output[2]) |
      (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign mux_1978_nl = MUX_s_1_2_2(or_2102_nl, or_2100_nl, fsm_output[4]);
  assign mux_1980_nl = MUX_s_1_2_2(mux_1979_nl, mux_1978_nl, fsm_output[8]);
  assign or_2106_nl = (fsm_output[1]) | mux_1980_nl;
  assign or_2097_nl = (operator_64_false_acc_cse_11_sva[3:0]!=4'b1101) | (~ (fsm_output[2]))
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign or_2096_nl = (COMP_LOOP_acc_cse_12_sva[3:0]!=4'b1101) | (~ (fsm_output[2]))
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1976_nl = MUX_s_1_2_2(or_2097_nl, or_2096_nl, fsm_output[4]);
  assign or_2098_nl = (fsm_output[8]) | mux_1976_nl;
  assign or_2095_nl = (operator_64_false_acc_cse_13_sva[3:0]!=4'b1101) | (fsm_output[8])
      | (~ (fsm_output[4])) | (~ (fsm_output[2])) | (fsm_output[3]) | not_tmp_312;
  assign mux_1977_nl = MUX_s_1_2_2(or_2098_nl, or_2095_nl, fsm_output[1]);
  assign mux_1981_nl = MUX_s_1_2_2(or_2106_nl, mux_1977_nl, fsm_output[9]);
  assign mux_1990_nl = MUX_s_1_2_2(mux_1989_nl, mux_1981_nl, fsm_output[7]);
  assign or_2093_nl = (~ (fsm_output[8])) | (COMP_LOOP_acc_8_psp_sva[1:0]!=2'b11)
      | (fsm_output[4]) | (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b01) | (~ (fsm_output[2]))
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1972_nl = MUX_s_1_2_2(or_2093_nl, nand_tmp_94, fsm_output[1]);
  assign or_2090_nl = (COMP_LOOP_acc_8_psp_sva[1:0]!=2'b11) | (fsm_output[4]) | (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b01)
      | (~ (fsm_output[2])) | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1970_nl = MUX_s_1_2_2(or_1233_cse, or_2090_nl, fsm_output[8]);
  assign mux_1971_nl = MUX_s_1_2_2(mux_1970_nl, nand_tmp_94, fsm_output[1]);
  assign mux_1973_nl = MUX_s_1_2_2(mux_1972_nl, mux_1971_nl, STAGE_VEC_LOOP_j_sva_9_0[3]);
  assign nor_615_nl = ~((operator_64_false_acc_cse_10_sva[3:0]!=4'b1101) | (fsm_output[2])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]));
  assign nor_616_nl = ~((COMP_LOOP_acc_11_psp_sva[2:0]!=3'b110) | (~ (STAGE_VEC_LOOP_j_sva_9_0[0]))
      | (fsm_output[2]) | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]));
  assign mux_1967_nl = MUX_s_1_2_2(nor_615_nl, nor_616_nl, fsm_output[4]);
  assign and_785_nl = (operator_64_false_acc_cse_14_sva[3:0]==4'b1101) & (fsm_output[2])
      & (fsm_output[3]) & (~ (fsm_output[6])) & (fsm_output[5]);
  assign and_786_nl = (COMP_LOOP_acc_13_psp_sva[2:0]==3'b110) & (STAGE_VEC_LOOP_j_sva_9_0[0])
      & (fsm_output[2]) & (fsm_output[3]) & (~ (fsm_output[6])) & (fsm_output[5]);
  assign mux_1966_nl = MUX_s_1_2_2(and_785_nl, and_786_nl, fsm_output[4]);
  assign mux_1968_nl = MUX_s_1_2_2(mux_1967_nl, mux_1966_nl, fsm_output[8]);
  assign nand_93_nl = ~((fsm_output[1]) & mux_1968_nl);
  assign mux_1974_nl = MUX_s_1_2_2(mux_1973_nl, nand_93_nl, fsm_output[9]);
  assign or_2079_nl = (~((operator_64_false_acc_cse_4_sva[3:0]==4'b1101) & (fsm_output[4:2]==3'b101)))
      | not_tmp_312;
  assign or_2077_nl = (STAGE_VEC_LOOP_j_sva_9_0[2:0]!=3'b101) | (~ (COMP_LOOP_acc_10_psp_sva[0]))
      | (fsm_output[2]) | not_tmp_311;
  assign or_2075_nl = (operator_64_false_acc_cse_8_sva[3:0]!=4'b1101) | (fsm_output[2])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]);
  assign mux_1962_nl = MUX_s_1_2_2(or_2077_nl, or_2075_nl, fsm_output[4]);
  assign mux_1963_nl = MUX_s_1_2_2(or_2079_nl, mux_1962_nl, fsm_output[8]);
  assign or_2073_nl = (operator_64_false_acc_cse_2_sva[3:0]!=4'b1101) | (fsm_output[2])
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign or_2072_nl = (COMP_LOOP_acc_7_psp_sva[2:0]!=3'b110) | (~ (STAGE_VEC_LOOP_j_sva_9_0[0]))
      | (fsm_output[2]) | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1961_nl = MUX_s_1_2_2(or_2073_nl, or_2072_nl, fsm_output[4]);
  assign or_2074_nl = (fsm_output[8]) | mux_1961_nl;
  assign mux_1964_nl = MUX_s_1_2_2(mux_1963_nl, or_2074_nl, fsm_output[1]);
  assign nand_267_nl = ~((COMP_LOOP_acc_12_psp_sva[1:0]==2'b11) & (STAGE_VEC_LOOP_j_sva_9_0[1:0]==2'b01)
      & (fsm_output[2]) & (fsm_output[3]) & (fsm_output[6]) & (~ (fsm_output[5])));
  assign nand_451_nl = ~((operator_64_false_acc_cse_12_sva[3:0]==4'b1101) & (fsm_output[2])
      & (fsm_output[3]) & (~ (fsm_output[6])) & (fsm_output[5]));
  assign mux_1959_nl = MUX_s_1_2_2(nand_267_nl, nand_451_nl, fsm_output[4]);
  assign or_2067_nl = (fsm_output[4]) | (operator_64_false_acc_cse_sva[3:0]!=4'b1101)
      | (fsm_output[2]) | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign mux_1960_nl = MUX_s_1_2_2(mux_1959_nl, or_2067_nl, fsm_output[8]);
  assign or_2071_nl = (fsm_output[1]) | mux_1960_nl;
  assign mux_1965_nl = MUX_s_1_2_2(mux_1964_nl, or_2071_nl, fsm_output[9]);
  assign mux_1975_nl = MUX_s_1_2_2(mux_1974_nl, mux_1965_nl, fsm_output[7]);
  assign mux_1991_nl = MUX_s_1_2_2(mux_1990_nl, mux_1975_nl, fsm_output[0]);
  assign vec_rsc_0_13_i_wea_d_pff = ~ mux_1991_nl;
  assign or_2171_nl = (operator_64_false_acc_cse_2_sva[3:0]!=4'b1101) | (fsm_output[4])
      | (fsm_output[0]) | (fsm_output[5]) | not_tmp_322;
  assign nand_248_nl = ~((COMP_LOOP_acc_cse_2_sva[3:0]==4'b1101) & (fsm_output[0])
      & COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm & (~ (fsm_output[5]))
      & (fsm_output[6]) & (fsm_output[3]) & (~ (fsm_output[2])));
  assign or_2168_nl = (COMP_LOOP_1_operator_64_false_acc_tmp[3:0]!=4'b1101) | (fsm_output[5])
      | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign or_2167_nl = (STAGE_VEC_LOOP_j_sva_9_0[3:0]!=4'b1101) | (fsm_output[5])
      | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign mux_2021_nl = MUX_s_1_2_2(or_2168_nl, or_2167_nl, fsm_output[0]);
  assign mux_2022_nl = MUX_s_1_2_2(nand_248_nl, mux_2021_nl, fsm_output[4]);
  assign mux_2023_nl = MUX_s_1_2_2(or_2171_nl, mux_2022_nl, fsm_output[1]);
  assign or_2166_nl = (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b110) | (~ (STAGE_VEC_LOOP_j_sva_9_0[0]))
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[5])
      | not_tmp_322;
  assign or_2164_nl = (operator_64_false_acc_cse_11_sva[3:0]!=4'b1101) | (fsm_output[5])
      | not_tmp_322;
  assign mux_2018_nl = MUX_s_1_2_2(or_2166_nl, or_2164_nl, fsm_output[0]);
  assign or_2162_nl = (fsm_output[0]) | (operator_64_false_acc_cse_10_sva[3:0]!=4'b1101)
      | (fsm_output[5]) | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign mux_2019_nl = MUX_s_1_2_2(mux_2018_nl, or_2162_nl, fsm_output[4]);
  assign or_2160_nl = (COMP_LOOP_acc_cse_10_sva[3:0]!=4'b1101) | (~ (fsm_output[4]))
      | (~ (fsm_output[0])) | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      | (fsm_output[5]) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign mux_2020_nl = MUX_s_1_2_2(mux_2019_nl, or_2160_nl, fsm_output[1]);
  assign mux_2024_nl = MUX_s_1_2_2(mux_2023_nl, mux_2020_nl, fsm_output[9]);
  assign nand_249_nl = ~((COMP_LOOP_acc_9_psp_sva[2:0]==3'b110) & (STAGE_VEC_LOOP_j_sva_9_0[0])
      & COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm & (fsm_output[5])
      & (fsm_output[6]) & (fsm_output[3]) & (~ (fsm_output[2])));
  assign nand_250_nl = ~((operator_64_false_acc_cse_7_sva[3:0]==4'b1101) & (fsm_output[5])
      & (fsm_output[6]) & (fsm_output[3]) & (~ (fsm_output[2])));
  assign mux_2014_nl = MUX_s_1_2_2(nand_249_nl, nand_250_nl, fsm_output[0]);
  assign or_2157_nl = (operator_64_false_acc_cse_6_sva[3:0]!=4'b1101) | (fsm_output[0])
      | (~ (fsm_output[5])) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign mux_2015_nl = MUX_s_1_2_2(mux_2014_nl, or_2157_nl, fsm_output[4]);
  assign or_2156_nl = (COMP_LOOP_acc_cse_6_sva[3:0]!=4'b1101) | (fsm_output[4]) |
      (~ (fsm_output[0])) | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      | (fsm_output[6:5]!=2'b01) | nand_442_cse;
  assign mux_2016_nl = MUX_s_1_2_2(mux_2015_nl, or_2156_nl, fsm_output[1]);
  assign nand_251_nl = ~((COMP_LOOP_acc_cse_sva[3:0]==4'b1101) & operator_64_false_slc_operator_64_false_acc_1_60_itm
      & (fsm_output[0]) & (fsm_output[5]) & (fsm_output[6]) & (fsm_output[3]) & (~
      (fsm_output[2])));
  assign or_2153_nl = (COMP_LOOP_acc_13_psp_sva[2:0]!=3'b110) | (~ (STAGE_VEC_LOOP_j_sva_9_0[0]))
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (~
      (fsm_output[5])) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign or_2152_nl = (operator_64_false_acc_cse_15_sva[3:0]!=4'b1101) | (~ (fsm_output[5]))
      | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign mux_2011_nl = MUX_s_1_2_2(or_2153_nl, or_2152_nl, fsm_output[0]);
  assign mux_2012_nl = MUX_s_1_2_2(nand_251_nl, mux_2011_nl, fsm_output[4]);
  assign or_2151_nl = (operator_64_false_acc_cse_sva[3:0]!=4'b1101) | (fsm_output[4])
      | (fsm_output[0]) | (~ (fsm_output[5])) | (~ (fsm_output[6])) | (~ (fsm_output[3]))
      | (fsm_output[2]);
  assign mux_2013_nl = MUX_s_1_2_2(mux_2012_nl, or_2151_nl, fsm_output[1]);
  assign mux_2017_nl = MUX_s_1_2_2(mux_2016_nl, mux_2013_nl, fsm_output[9]);
  assign mux_2025_nl = MUX_s_1_2_2(mux_2024_nl, mux_2017_nl, fsm_output[8]);
  assign or_2150_nl = (COMP_LOOP_acc_7_psp_sva[2:0]!=3'b110) | (~ (STAGE_VEC_LOOP_j_sva_9_0[0]))
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[5])
      | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign or_2148_nl = (operator_64_false_acc_cse_3_sva[3:0]!=4'b1101) | (fsm_output[5])
      | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign mux_2006_nl = MUX_s_1_2_2(or_2150_nl, or_2148_nl, fsm_output[0]);
  assign or_2146_nl = (~(operator_64_false_slc_operator_64_false_acc_1_60_itm & (COMP_LOOP_acc_cse_4_sva[3:0]==4'b1101)
      & (fsm_output[0]) & (fsm_output[5]) & (~ (fsm_output[6])))) | nand_442_cse;
  assign mux_2007_nl = MUX_s_1_2_2(mux_2006_nl, or_2146_nl, fsm_output[4]);
  assign nand_465_nl = ~((STAGE_VEC_LOOP_j_sva_9_0[1:0]==2'b01) & (COMP_LOOP_acc_8_psp_sva[1:0]==2'b11)
      & COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm & (fsm_output[5])
      & (fsm_output[6]) & (~ (fsm_output[3])) & (fsm_output[2]));
  assign nand_254_nl = ~((STAGE_VEC_LOOP_j_sva_9_0[1:0]==2'b01) & (COMP_LOOP_acc_8_psp_sva[1:0]==2'b11)
      & COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm);
  assign mux_2003_nl = MUX_s_1_2_2(nand_tmp_19, or_tmp_669, nand_254_nl);
  assign and_540_nl = (operator_64_false_acc_cse_4_sva[3:0]==4'b1101);
  assign mux_2004_nl = MUX_s_1_2_2(nand_465_nl, mux_2003_nl, and_540_nl);
  assign nand_461_nl = ~((operator_64_false_acc_cse_5_sva[3:0]==4'b1101) & (fsm_output[5])
      & (fsm_output[6]) & (~ (fsm_output[3])) & (fsm_output[2]));
  assign mux_2005_nl = MUX_s_1_2_2(mux_2004_nl, nand_461_nl, fsm_output[0]);
  assign nand_98_nl = ~((fsm_output[4]) & (~ mux_2005_nl));
  assign mux_2008_nl = MUX_s_1_2_2(mux_2007_nl, nand_98_nl, fsm_output[1]);
  assign or_2139_nl = (COMP_LOOP_acc_cse_12_sva[3:0]!=4'b1101) | (~ operator_64_false_slc_operator_64_false_acc_1_60_itm)
      | (~ (fsm_output[0])) | (fsm_output[5]) | (fsm_output[6]) | (fsm_output[3])
      | (~ (fsm_output[2]));
  assign or_2137_nl = (operator_64_false_acc_cse_14_sva[3:0]!=4'b1101) | (fsm_output[0])
      | (~ (fsm_output[5])) | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign mux_2001_nl = MUX_s_1_2_2(or_2139_nl, or_2137_nl, fsm_output[4]);
  assign or_2136_nl = (operator_64_false_acc_cse_12_sva[3:0]!=4'b1101) | (fsm_output[0])
      | (fsm_output[5]) | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign or_2134_nl = (~((COMP_LOOP_acc_12_psp_sva[1:0]==2'b11) & (STAGE_VEC_LOOP_j_sva_9_0[1:0]==2'b01)
      & COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm & (fsm_output[6:5]==2'b01)))
      | nand_442_cse;
  assign or_2132_nl = (operator_64_false_acc_cse_13_sva[3:0]!=4'b1101) | (fsm_output[6:5]!=2'b01)
      | nand_442_cse;
  assign and_541_nl = (operator_64_false_acc_cse_13_sva[3:0]==4'b1101);
  assign mux_1997_nl = MUX_s_1_2_2(nand_437_cse, mux_1112_cse, and_541_nl);
  assign and_542_nl = (COMP_LOOP_acc_cse_14_sva[3:0]==4'b1101);
  assign mux_1998_nl = MUX_s_1_2_2(or_2132_nl, mux_1997_nl, and_542_nl);
  assign mux_1999_nl = MUX_s_1_2_2(or_2134_nl, mux_1998_nl, fsm_output[0]);
  assign mux_2000_nl = MUX_s_1_2_2(or_2136_nl, mux_1999_nl, fsm_output[4]);
  assign mux_2002_nl = MUX_s_1_2_2(mux_2001_nl, mux_2000_nl, fsm_output[1]);
  assign mux_2009_nl = MUX_s_1_2_2(mux_2008_nl, mux_2002_nl, fsm_output[9]);
  assign or_2124_nl = (COMP_LOOP_acc_cse_8_sva[3:0]!=4'b1101) | (fsm_output[4]) |
      (~ operator_64_false_slc_operator_64_false_acc_1_60_itm) | (~ (fsm_output[0]))
      | (~ (fsm_output[5])) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign or_2123_nl = (operator_64_false_acc_cse_8_sva[3:0]!=4'b1101) | (fsm_output[0])
      | (~ (fsm_output[5])) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign or_2122_nl = (STAGE_VEC_LOOP_j_sva_9_0[2:0]!=3'b101) | (~ (COMP_LOOP_acc_10_psp_sva[0]))
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[5])
      | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign or_2121_nl = (operator_64_false_acc_cse_9_sva[3:0]!=4'b1101) | (fsm_output[5])
      | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign mux_1992_nl = MUX_s_1_2_2(or_2122_nl, or_2121_nl, fsm_output[0]);
  assign mux_1993_nl = MUX_s_1_2_2(or_2123_nl, mux_1992_nl, fsm_output[4]);
  assign mux_1994_nl = MUX_s_1_2_2(or_2124_nl, mux_1993_nl, fsm_output[1]);
  assign or_2125_nl = (fsm_output[9]) | mux_1994_nl;
  assign mux_2010_nl = MUX_s_1_2_2(mux_2009_nl, or_2125_nl, fsm_output[8]);
  assign mux_2026_nl = MUX_s_1_2_2(mux_2025_nl, mux_2010_nl, fsm_output[7]);
  assign vec_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d = ~ mux_2026_nl;
  assign nor_597_nl = ~((operator_64_false_acc_cse_1_sva[3:0]!=4'b1110) | (fsm_output[2])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]));
  assign nor_598_nl = ~((COMP_LOOP_acc_cse_2_sva[3:0]!=4'b1110) | (fsm_output[2])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]));
  assign mux_2055_nl = MUX_s_1_2_2(nor_597_nl, nor_598_nl, fsm_output[4]);
  assign and_770_nl = (operator_64_false_acc_cse_5_sva[3:0]==4'b1110) & (fsm_output[2])
      & (fsm_output[3]) & (~ (fsm_output[6])) & (fsm_output[5]);
  assign and_776_nl = (COMP_LOOP_acc_cse_6_sva[3:0]==4'b1110) & (fsm_output[2]) &
      (fsm_output[3]) & (~ (fsm_output[6])) & (fsm_output[5]);
  assign mux_2054_nl = MUX_s_1_2_2(and_770_nl, and_776_nl, fsm_output[4]);
  assign mux_2056_nl = MUX_s_1_2_2(mux_2055_nl, mux_2054_nl, fsm_output[8]);
  assign nand_102_nl = ~((fsm_output[1]) & mux_2056_nl);
  assign nor_601_nl = ~((operator_64_false_acc_cse_15_sva[3:0]!=4'b1110) | (fsm_output[2])
      | not_tmp_311);
  assign nor_602_nl = ~((COMP_LOOP_acc_cse_sva[3:0]!=4'b1110) | (fsm_output[2]) |
      not_tmp_311);
  assign mux_2052_nl = MUX_s_1_2_2(nor_601_nl, nor_602_nl, fsm_output[4]);
  assign nand_101_nl = ~((fsm_output[8]) & mux_2052_nl);
  assign or_2216_nl = (COMP_LOOP_acc_cse_10_sva[3:0]!=4'b1110) | (fsm_output[2])
      | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign or_2214_nl = (operator_64_false_acc_cse_9_sva[3:0]!=4'b1110) | (fsm_output[2])
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_2050_nl = MUX_s_1_2_2(or_2216_nl, or_2214_nl, fsm_output[4]);
  assign or_2213_nl = (fsm_output[4]) | (COMP_LOOP_acc_cse_14_sva[3:0]!=4'b1110)
      | (~ (fsm_output[2])) | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_2051_nl = MUX_s_1_2_2(mux_2050_nl, or_2213_nl, fsm_output[8]);
  assign mux_2053_nl = MUX_s_1_2_2(nand_101_nl, mux_2051_nl, fsm_output[1]);
  assign mux_2057_nl = MUX_s_1_2_2(nand_102_nl, mux_2053_nl, fsm_output[9]);
  assign nand_239_nl = ~((COMP_LOOP_acc_cse_4_sva[3:0]==4'b1110) & (fsm_output[2])
      & (fsm_output[3]) & (fsm_output[6]) & (~ (fsm_output[5])));
  assign nand_469_nl = ~((operator_64_false_acc_cse_3_sva[3:0]==4'b1110) & (fsm_output[2])
      & (fsm_output[3]) & (~ (fsm_output[6])) & (fsm_output[5]));
  assign mux_2047_nl = MUX_s_1_2_2(nand_239_nl, nand_469_nl, fsm_output[4]);
  assign or_2208_nl = (operator_64_false_acc_cse_7_sva[3:0]!=4'b1110) | (fsm_output[2])
      | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign or_2206_nl = (COMP_LOOP_acc_cse_8_sva[3:0]!=4'b1110) | (fsm_output[2]) |
      (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign mux_2046_nl = MUX_s_1_2_2(or_2208_nl, or_2206_nl, fsm_output[4]);
  assign mux_2048_nl = MUX_s_1_2_2(mux_2047_nl, mux_2046_nl, fsm_output[8]);
  assign or_2212_nl = (fsm_output[1]) | mux_2048_nl;
  assign or_2203_nl = (operator_64_false_acc_cse_11_sva[3:0]!=4'b1110) | (~ (fsm_output[2]))
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign or_2202_nl = (COMP_LOOP_acc_cse_12_sva[3:0]!=4'b1110) | (~ (fsm_output[2]))
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_2044_nl = MUX_s_1_2_2(or_2203_nl, or_2202_nl, fsm_output[4]);
  assign or_2204_nl = (fsm_output[8]) | mux_2044_nl;
  assign or_2201_nl = (operator_64_false_acc_cse_13_sva[3:0]!=4'b1110) | (fsm_output[8])
      | (~ (fsm_output[4])) | (~ (fsm_output[2])) | (fsm_output[3]) | not_tmp_312;
  assign mux_2045_nl = MUX_s_1_2_2(or_2204_nl, or_2201_nl, fsm_output[1]);
  assign mux_2049_nl = MUX_s_1_2_2(or_2212_nl, mux_2045_nl, fsm_output[9]);
  assign mux_2058_nl = MUX_s_1_2_2(mux_2057_nl, mux_2049_nl, fsm_output[7]);
  assign or_2199_nl = (~ (fsm_output[8])) | (COMP_LOOP_acc_8_psp_sva[1:0]!=2'b11)
      | (fsm_output[4]) | (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b10) | (~ (fsm_output[2]))
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_2040_nl = MUX_s_1_2_2(or_2199_nl, nand_tmp_100, fsm_output[1]);
  assign or_2196_nl = (COMP_LOOP_acc_8_psp_sva[1:0]!=2'b11) | (fsm_output[4]) | (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b10)
      | (~ (fsm_output[2])) | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_2038_nl = MUX_s_1_2_2(or_1339_cse, or_2196_nl, fsm_output[8]);
  assign mux_2039_nl = MUX_s_1_2_2(mux_2038_nl, nand_tmp_100, fsm_output[1]);
  assign mux_2041_nl = MUX_s_1_2_2(mux_2040_nl, mux_2039_nl, STAGE_VEC_LOOP_j_sva_9_0[3]);
  assign nor_603_nl = ~((operator_64_false_acc_cse_10_sva[3:0]!=4'b1110) | (fsm_output[2])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]));
  assign nor_604_nl = ~((COMP_LOOP_acc_11_psp_sva[2:0]!=3'b111) | (STAGE_VEC_LOOP_j_sva_9_0[0])
      | (fsm_output[2]) | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]));
  assign mux_2035_nl = MUX_s_1_2_2(nor_603_nl, nor_604_nl, fsm_output[4]);
  assign and_783_nl = (operator_64_false_acc_cse_14_sva[3:0]==4'b1110) & (fsm_output[2])
      & (fsm_output[3]) & (~ (fsm_output[6])) & (fsm_output[5]);
  assign and_784_nl = (COMP_LOOP_acc_13_psp_sva[2:0]==3'b111) & (~ (STAGE_VEC_LOOP_j_sva_9_0[0]))
      & (fsm_output[2]) & (fsm_output[3]) & (~ (fsm_output[6])) & (fsm_output[5]);
  assign mux_2034_nl = MUX_s_1_2_2(and_783_nl, and_784_nl, fsm_output[4]);
  assign mux_2036_nl = MUX_s_1_2_2(mux_2035_nl, mux_2034_nl, fsm_output[8]);
  assign nand_99_nl = ~((fsm_output[1]) & mux_2036_nl);
  assign mux_2042_nl = MUX_s_1_2_2(mux_2041_nl, nand_99_nl, fsm_output[9]);
  assign or_2185_nl = (~((operator_64_false_acc_cse_4_sva[3:0]==4'b1110) & (fsm_output[4:2]==3'b101)))
      | not_tmp_312;
  assign or_2183_nl = (STAGE_VEC_LOOP_j_sva_9_0[2:0]!=3'b110) | (~ (COMP_LOOP_acc_10_psp_sva[0]))
      | (fsm_output[2]) | not_tmp_311;
  assign or_2181_nl = (operator_64_false_acc_cse_8_sva[3:0]!=4'b1110) | (fsm_output[2])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[5]);
  assign mux_2030_nl = MUX_s_1_2_2(or_2183_nl, or_2181_nl, fsm_output[4]);
  assign mux_2031_nl = MUX_s_1_2_2(or_2185_nl, mux_2030_nl, fsm_output[8]);
  assign or_2179_nl = (operator_64_false_acc_cse_2_sva[3:0]!=4'b1110) | (fsm_output[2])
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign or_2178_nl = (COMP_LOOP_acc_7_psp_sva[2:0]!=3'b111) | (STAGE_VEC_LOOP_j_sva_9_0[0])
      | (fsm_output[2]) | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_2029_nl = MUX_s_1_2_2(or_2179_nl, or_2178_nl, fsm_output[4]);
  assign or_2180_nl = (fsm_output[8]) | mux_2029_nl;
  assign mux_2032_nl = MUX_s_1_2_2(mux_2031_nl, or_2180_nl, fsm_output[1]);
  assign nand_244_nl = ~((COMP_LOOP_acc_12_psp_sva[1:0]==2'b11) & (STAGE_VEC_LOOP_j_sva_9_0[1:0]==2'b10)
      & (fsm_output[2]) & (fsm_output[3]) & (fsm_output[6]) & (~ (fsm_output[5])));
  assign nand_450_nl = ~((operator_64_false_acc_cse_12_sva[3:0]==4'b1110) & (fsm_output[2])
      & (fsm_output[3]) & (~ (fsm_output[6])) & (fsm_output[5]));
  assign mux_2027_nl = MUX_s_1_2_2(nand_244_nl, nand_450_nl, fsm_output[4]);
  assign or_2173_nl = (fsm_output[4]) | (operator_64_false_acc_cse_sva[3:0]!=4'b1110)
      | (fsm_output[2]) | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign mux_2028_nl = MUX_s_1_2_2(mux_2027_nl, or_2173_nl, fsm_output[8]);
  assign or_2177_nl = (fsm_output[1]) | mux_2028_nl;
  assign mux_2033_nl = MUX_s_1_2_2(mux_2032_nl, or_2177_nl, fsm_output[9]);
  assign mux_2043_nl = MUX_s_1_2_2(mux_2042_nl, mux_2033_nl, fsm_output[7]);
  assign mux_2059_nl = MUX_s_1_2_2(mux_2058_nl, mux_2043_nl, fsm_output[0]);
  assign vec_rsc_0_14_i_wea_d_pff = ~ mux_2059_nl;
  assign or_2280_nl = (operator_64_false_acc_cse_2_sva[3:0]!=4'b1110) | (fsm_output[4])
      | (fsm_output[0]) | (fsm_output[5]) | not_tmp_322;
  assign nand_222_nl = ~((COMP_LOOP_acc_cse_2_sva[3:0]==4'b1110) & (fsm_output[0])
      & COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm & (~ (fsm_output[5]))
      & (fsm_output[6]) & (fsm_output[3]) & (~ (fsm_output[2])));
  assign or_2277_nl = (COMP_LOOP_1_operator_64_false_acc_tmp[3:0]!=4'b1110) | (fsm_output[5])
      | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign or_2276_nl = (STAGE_VEC_LOOP_j_sva_9_0[3:0]!=4'b1110) | (fsm_output[5])
      | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign mux_2089_nl = MUX_s_1_2_2(or_2277_nl, or_2276_nl, fsm_output[0]);
  assign mux_2090_nl = MUX_s_1_2_2(nand_222_nl, mux_2089_nl, fsm_output[4]);
  assign mux_2091_nl = MUX_s_1_2_2(or_2280_nl, mux_2090_nl, fsm_output[1]);
  assign or_2275_nl = (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b111) | (STAGE_VEC_LOOP_j_sva_9_0[0])
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[5])
      | not_tmp_322;
  assign or_2273_nl = (operator_64_false_acc_cse_11_sva[3:0]!=4'b1110) | (fsm_output[5])
      | not_tmp_322;
  assign mux_2086_nl = MUX_s_1_2_2(or_2275_nl, or_2273_nl, fsm_output[0]);
  assign or_2271_nl = (fsm_output[0]) | (operator_64_false_acc_cse_10_sva[3:0]!=4'b1110)
      | (fsm_output[5]) | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign mux_2087_nl = MUX_s_1_2_2(mux_2086_nl, or_2271_nl, fsm_output[4]);
  assign or_2269_nl = (~ (fsm_output[4])) | (~ (fsm_output[0])) | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      | (COMP_LOOP_acc_cse_10_sva[3:0]!=4'b1110) | (fsm_output[5]) | (fsm_output[6])
      | (fsm_output[3]) | (fsm_output[2]);
  assign mux_2088_nl = MUX_s_1_2_2(mux_2087_nl, or_2269_nl, fsm_output[1]);
  assign mux_2092_nl = MUX_s_1_2_2(mux_2091_nl, mux_2088_nl, fsm_output[9]);
  assign nand_223_nl = ~((COMP_LOOP_acc_9_psp_sva[2:0]==3'b111) & (~ (STAGE_VEC_LOOP_j_sva_9_0[0]))
      & COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm & (fsm_output[5])
      & (fsm_output[6]) & (fsm_output[3]) & (~ (fsm_output[2])));
  assign nand_224_nl = ~((operator_64_false_acc_cse_7_sva[3:0]==4'b1110) & (fsm_output[5])
      & (fsm_output[6]) & (fsm_output[3]) & (~ (fsm_output[2])));
  assign mux_2082_nl = MUX_s_1_2_2(nand_223_nl, nand_224_nl, fsm_output[0]);
  assign or_2266_nl = (operator_64_false_acc_cse_6_sva[3:0]!=4'b1110) | (fsm_output[0])
      | (~ (fsm_output[5])) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign mux_2083_nl = MUX_s_1_2_2(mux_2082_nl, or_2266_nl, fsm_output[4]);
  assign or_2265_nl = (COMP_LOOP_acc_cse_6_sva[3:0]!=4'b1110) | (fsm_output[4]) |
      (~ (fsm_output[0])) | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      | (fsm_output[6:5]!=2'b01) | nand_442_cse;
  assign mux_2084_nl = MUX_s_1_2_2(mux_2083_nl, or_2265_nl, fsm_output[1]);
  assign nand_225_nl = ~(operator_64_false_slc_operator_64_false_acc_1_60_itm & (fsm_output[0])
      & (COMP_LOOP_acc_cse_sva[3:0]==4'b1110) & (fsm_output[5]) & (fsm_output[6])
      & (fsm_output[3]) & (~ (fsm_output[2])));
  assign or_2262_nl = (COMP_LOOP_acc_13_psp_sva[2:0]!=3'b111) | (STAGE_VEC_LOOP_j_sva_9_0[0])
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (~
      (fsm_output[5])) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign or_2261_nl = (operator_64_false_acc_cse_15_sva[3:0]!=4'b1110) | (~ (fsm_output[5]))
      | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign mux_2079_nl = MUX_s_1_2_2(or_2262_nl, or_2261_nl, fsm_output[0]);
  assign mux_2080_nl = MUX_s_1_2_2(nand_225_nl, mux_2079_nl, fsm_output[4]);
  assign or_2260_nl = (operator_64_false_acc_cse_sva[3:0]!=4'b1110) | (fsm_output[4])
      | (fsm_output[0]) | (~ (fsm_output[5])) | (~ (fsm_output[6])) | (~ (fsm_output[3]))
      | (fsm_output[2]);
  assign mux_2081_nl = MUX_s_1_2_2(mux_2080_nl, or_2260_nl, fsm_output[1]);
  assign mux_2085_nl = MUX_s_1_2_2(mux_2084_nl, mux_2081_nl, fsm_output[9]);
  assign mux_2093_nl = MUX_s_1_2_2(mux_2092_nl, mux_2085_nl, fsm_output[8]);
  assign or_2259_nl = (COMP_LOOP_acc_7_psp_sva[2:0]!=3'b111) | (STAGE_VEC_LOOP_j_sva_9_0[0])
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[5])
      | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign or_2257_nl = (operator_64_false_acc_cse_3_sva[3:0]!=4'b1110) | (fsm_output[5])
      | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign mux_2074_nl = MUX_s_1_2_2(or_2259_nl, or_2257_nl, fsm_output[0]);
  assign or_2255_nl = (~(operator_64_false_slc_operator_64_false_acc_1_60_itm & (COMP_LOOP_acc_cse_4_sva[3:0]==4'b1110)
      & (fsm_output[0]) & (fsm_output[5]) & (~ (fsm_output[6])))) | nand_442_cse;
  assign mux_2075_nl = MUX_s_1_2_2(mux_2074_nl, or_2255_nl, fsm_output[4]);
  assign nand_227_nl = ~((STAGE_VEC_LOOP_j_sva_9_0[1:0]==2'b10) & (COMP_LOOP_acc_8_psp_sva[1:0]==2'b11)
      & COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm);
  assign mux_2071_nl = MUX_s_1_2_2(nand_tmp_19, or_tmp_669, nand_227_nl);
  assign nand_464_nl = ~((STAGE_VEC_LOOP_j_sva_9_0[1:0]==2'b10) & (COMP_LOOP_acc_8_psp_sva[1:0]==2'b11)
      & COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm & (fsm_output[5])
      & (fsm_output[6]) & (~ (fsm_output[3])) & (fsm_output[2]));
  assign nand_229_nl = ~((operator_64_false_acc_cse_4_sva[3:0]==4'b1110));
  assign mux_2072_nl = MUX_s_1_2_2(mux_2071_nl, nand_464_nl, nand_229_nl);
  assign nand_460_nl = ~((operator_64_false_acc_cse_5_sva[3:0]==4'b1110) & (fsm_output[5])
      & (fsm_output[6]) & (~ (fsm_output[3])) & (fsm_output[2]));
  assign mux_2073_nl = MUX_s_1_2_2(mux_2072_nl, nand_460_nl, fsm_output[0]);
  assign nand_104_nl = ~((fsm_output[4]) & (~ mux_2073_nl));
  assign mux_2076_nl = MUX_s_1_2_2(mux_2075_nl, nand_104_nl, fsm_output[1]);
  assign or_2247_nl = (~ operator_64_false_slc_operator_64_false_acc_1_60_itm) |
      (~ (fsm_output[0])) | (COMP_LOOP_acc_cse_12_sva[3:0]!=4'b1110) | (fsm_output[5])
      | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign or_2245_nl = (operator_64_false_acc_cse_14_sva[3:0]!=4'b1110) | (fsm_output[0])
      | (~ (fsm_output[5])) | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign mux_2069_nl = MUX_s_1_2_2(or_2247_nl, or_2245_nl, fsm_output[4]);
  assign or_2244_nl = (operator_64_false_acc_cse_12_sva[3:0]!=4'b1110) | (fsm_output[0])
      | (fsm_output[5]) | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign or_2242_nl = (~((COMP_LOOP_acc_12_psp_sva[1:0]==2'b11) & (STAGE_VEC_LOOP_j_sva_9_0[1:0]==2'b10)
      & COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm & (fsm_output[6:5]==2'b01)))
      | nand_442_cse;
  assign nand_233_nl = ~((operator_64_false_acc_cse_13_sva[3:0]==4'b1110));
  assign mux_2065_nl = MUX_s_1_2_2(mux_1112_cse, nand_437_cse, nand_233_nl);
  assign or_2234_nl = (operator_64_false_acc_cse_13_sva[3:0]!=4'b1110) | (fsm_output[6:5]!=2'b01)
      | nand_442_cse;
  assign nand_234_nl = ~((COMP_LOOP_acc_cse_14_sva[3:0]==4'b1110));
  assign mux_2066_nl = MUX_s_1_2_2(mux_2065_nl, or_2234_nl, nand_234_nl);
  assign mux_2067_nl = MUX_s_1_2_2(or_2242_nl, mux_2066_nl, fsm_output[0]);
  assign mux_2068_nl = MUX_s_1_2_2(or_2244_nl, mux_2067_nl, fsm_output[4]);
  assign mux_2070_nl = MUX_s_1_2_2(mux_2069_nl, mux_2068_nl, fsm_output[1]);
  assign mux_2077_nl = MUX_s_1_2_2(mux_2076_nl, mux_2070_nl, fsm_output[9]);
  assign or_2230_nl = (COMP_LOOP_acc_cse_8_sva[3:0]!=4'b1110) | (fsm_output[4]) |
      (~ operator_64_false_slc_operator_64_false_acc_1_60_itm) | (~ (fsm_output[0]))
      | (~ (fsm_output[5])) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign or_2229_nl = (operator_64_false_acc_cse_8_sva[3:0]!=4'b1110) | (fsm_output[0])
      | (~ (fsm_output[5])) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2]);
  assign or_2228_nl = (STAGE_VEC_LOOP_j_sva_9_0[2:0]!=3'b110) | (~ (COMP_LOOP_acc_10_psp_sva[0]))
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[5])
      | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign or_2227_nl = (operator_64_false_acc_cse_9_sva[3:0]!=4'b1110) | (fsm_output[5])
      | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[2]);
  assign mux_2060_nl = MUX_s_1_2_2(or_2228_nl, or_2227_nl, fsm_output[0]);
  assign mux_2061_nl = MUX_s_1_2_2(or_2229_nl, mux_2060_nl, fsm_output[4]);
  assign mux_2062_nl = MUX_s_1_2_2(or_2230_nl, mux_2061_nl, fsm_output[1]);
  assign or_2231_nl = (fsm_output[9]) | mux_2062_nl;
  assign mux_2078_nl = MUX_s_1_2_2(mux_2077_nl, or_2231_nl, fsm_output[8]);
  assign mux_2094_nl = MUX_s_1_2_2(mux_2093_nl, mux_2078_nl, fsm_output[7]);
  assign vec_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d = ~ mux_2094_nl;
  assign and_536_nl = (operator_64_false_acc_cse_1_sva[3:0]==4'b1111) & (~ (fsm_output[2]))
      & (fsm_output[3]) & (fsm_output[6]) & (~ (fsm_output[5]));
  assign and_537_nl = (COMP_LOOP_acc_cse_2_sva[3:0]==4'b1111) & (~ (fsm_output[2]))
      & (fsm_output[3]) & (fsm_output[6]) & (~ (fsm_output[5]));
  assign mux_2123_nl = MUX_s_1_2_2(and_536_nl, and_537_nl, fsm_output[4]);
  assign and_769_nl = (operator_64_false_acc_cse_5_sva[3:0]==4'b1111) & (fsm_output[2])
      & (fsm_output[3]) & (~ (fsm_output[6])) & (fsm_output[5]);
  assign and_775_nl = (COMP_LOOP_acc_cse_6_sva[3:0]==4'b1111) & (fsm_output[2]) &
      (fsm_output[3]) & (~ (fsm_output[6])) & (fsm_output[5]);
  assign mux_2122_nl = MUX_s_1_2_2(and_769_nl, and_775_nl, fsm_output[4]);
  assign mux_2124_nl = MUX_s_1_2_2(mux_2123_nl, mux_2122_nl, fsm_output[8]);
  assign nand_108_nl = ~((fsm_output[1]) & mux_2124_nl);
  assign nor_591_nl = ~((~((operator_64_false_acc_cse_15_sva[3:0]==4'b1111) & (~
      (fsm_output[2])))) | not_tmp_311);
  assign nor_592_nl = ~((~((COMP_LOOP_acc_cse_sva[3:0]==4'b1111) & (~ (fsm_output[2]))))
      | not_tmp_311);
  assign mux_2120_nl = MUX_s_1_2_2(nor_591_nl, nor_592_nl, fsm_output[4]);
  assign nand_107_nl = ~((fsm_output[8]) & mux_2120_nl);
  assign or_2325_nl = (COMP_LOOP_acc_cse_10_sva[3:0]!=4'b1111) | (fsm_output[2])
      | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign or_2323_nl = (operator_64_false_acc_cse_9_sva[3:0]!=4'b1111) | (fsm_output[2])
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_2118_nl = MUX_s_1_2_2(or_2325_nl, or_2323_nl, fsm_output[4]);
  assign or_2322_nl = (fsm_output[4]) | (COMP_LOOP_acc_cse_14_sva[3:0]!=4'b1111)
      | (~ (fsm_output[2])) | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_2119_nl = MUX_s_1_2_2(mux_2118_nl, or_2322_nl, fsm_output[8]);
  assign mux_2121_nl = MUX_s_1_2_2(nand_107_nl, mux_2119_nl, fsm_output[1]);
  assign mux_2125_nl = MUX_s_1_2_2(nand_108_nl, mux_2121_nl, fsm_output[9]);
  assign nand_208_nl = ~((COMP_LOOP_acc_cse_4_sva[3:0]==4'b1111) & (fsm_output[2])
      & (fsm_output[3]) & (fsm_output[6]) & (~ (fsm_output[5])));
  assign nand_468_nl = ~((operator_64_false_acc_cse_3_sva[3:0]==4'b1111) & (fsm_output[2])
      & (fsm_output[3]) & (~ (fsm_output[6])) & (fsm_output[5]));
  assign mux_2115_nl = MUX_s_1_2_2(nand_208_nl, nand_468_nl, fsm_output[4]);
  assign or_2317_nl = (operator_64_false_acc_cse_7_sva[3:0]!=4'b1111) | (fsm_output[2])
      | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign or_2315_nl = (COMP_LOOP_acc_cse_8_sva[3:0]!=4'b1111) | (fsm_output[2]) |
      (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign mux_2114_nl = MUX_s_1_2_2(or_2317_nl, or_2315_nl, fsm_output[4]);
  assign mux_2116_nl = MUX_s_1_2_2(mux_2115_nl, mux_2114_nl, fsm_output[8]);
  assign or_2321_nl = (fsm_output[1]) | mux_2116_nl;
  assign or_2312_nl = (operator_64_false_acc_cse_11_sva[3:0]!=4'b1111) | (~ (fsm_output[2]))
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign or_2311_nl = (COMP_LOOP_acc_cse_12_sva[3:0]!=4'b1111) | (~ (fsm_output[2]))
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_2112_nl = MUX_s_1_2_2(or_2312_nl, or_2311_nl, fsm_output[4]);
  assign or_2313_nl = (fsm_output[8]) | mux_2112_nl;
  assign or_2310_nl = (~((operator_64_false_acc_cse_13_sva[3:0]==4'b1111) & (~ (fsm_output[8]))
      & (fsm_output[4]) & (fsm_output[2]) & (~ (fsm_output[3])))) | not_tmp_312;
  assign mux_2113_nl = MUX_s_1_2_2(or_2313_nl, or_2310_nl, fsm_output[1]);
  assign mux_2117_nl = MUX_s_1_2_2(or_2321_nl, mux_2113_nl, fsm_output[9]);
  assign mux_2126_nl = MUX_s_1_2_2(mux_2125_nl, mux_2117_nl, fsm_output[7]);
  assign or_2308_nl = (~ (fsm_output[8])) | (COMP_LOOP_acc_8_psp_sva[1:0]!=2'b11)
      | (fsm_output[4]) | (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b11) | (~ (fsm_output[2]))
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_2108_nl = MUX_s_1_2_2(or_2308_nl, nand_tmp_106, fsm_output[1]);
  assign or_2305_nl = (COMP_LOOP_acc_8_psp_sva[1:0]!=2'b11) | (fsm_output[4]) | (STAGE_VEC_LOOP_j_sva_9_0[1:0]!=2'b11)
      | (~ (fsm_output[2])) | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_2106_nl = MUX_s_1_2_2(or_1448_cse, or_2305_nl, fsm_output[8]);
  assign mux_2107_nl = MUX_s_1_2_2(mux_2106_nl, nand_tmp_106, fsm_output[1]);
  assign mux_2109_nl = MUX_s_1_2_2(mux_2108_nl, mux_2107_nl, STAGE_VEC_LOOP_j_sva_9_0[3]);
  assign and_538_nl = (operator_64_false_acc_cse_10_sva[3:0]==4'b1111) & (~ (fsm_output[2]))
      & (fsm_output[3]) & (fsm_output[6]) & (~ (fsm_output[5]));
  assign and_539_nl = (COMP_LOOP_acc_11_psp_sva[2:0]==3'b111) & (STAGE_VEC_LOOP_j_sva_9_0[0])
      & (~ (fsm_output[2])) & (fsm_output[3]) & (fsm_output[6]) & (~ (fsm_output[5]));
  assign mux_2103_nl = MUX_s_1_2_2(and_538_nl, and_539_nl, fsm_output[4]);
  assign and_781_nl = (operator_64_false_acc_cse_14_sva[3:0]==4'b1111) & (fsm_output[2])
      & (fsm_output[3]) & (~ (fsm_output[6])) & (fsm_output[5]);
  assign and_782_nl = (COMP_LOOP_acc_13_psp_sva[2:0]==3'b111) & (STAGE_VEC_LOOP_j_sva_9_0[0])
      & (fsm_output[2]) & (fsm_output[3]) & (~ (fsm_output[6])) & (fsm_output[5]);
  assign mux_2102_nl = MUX_s_1_2_2(and_781_nl, and_782_nl, fsm_output[4]);
  assign mux_2104_nl = MUX_s_1_2_2(mux_2103_nl, mux_2102_nl, fsm_output[8]);
  assign nand_105_nl = ~((fsm_output[1]) & mux_2104_nl);
  assign mux_2110_nl = MUX_s_1_2_2(mux_2109_nl, nand_105_nl, fsm_output[9]);
  assign or_2294_nl = (~((operator_64_false_acc_cse_4_sva[3:0]==4'b1111) & (fsm_output[4:2]==3'b101)))
      | not_tmp_312;
  assign or_2292_nl = (~((STAGE_VEC_LOOP_j_sva_9_0[2:0]==3'b111) & (COMP_LOOP_acc_10_psp_sva[0])
      & (~ (fsm_output[2])))) | not_tmp_311;
  assign nand_215_nl = ~((operator_64_false_acc_cse_8_sva[3:0]==4'b1111) & (~ (fsm_output[2]))
      & (fsm_output[3]) & (fsm_output[6]) & (~ (fsm_output[5])));
  assign mux_2098_nl = MUX_s_1_2_2(or_2292_nl, nand_215_nl, fsm_output[4]);
  assign mux_2099_nl = MUX_s_1_2_2(or_2294_nl, mux_2098_nl, fsm_output[8]);
  assign or_2288_nl = (operator_64_false_acc_cse_2_sva[3:0]!=4'b1111) | (fsm_output[2])
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign or_2287_nl = (COMP_LOOP_acc_7_psp_sva[2:0]!=3'b111) | (~ (STAGE_VEC_LOOP_j_sva_9_0[0]))
      | (fsm_output[2]) | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_2097_nl = MUX_s_1_2_2(or_2288_nl, or_2287_nl, fsm_output[4]);
  assign or_2289_nl = (fsm_output[8]) | mux_2097_nl;
  assign mux_2100_nl = MUX_s_1_2_2(mux_2099_nl, or_2289_nl, fsm_output[1]);
  assign nand_216_nl = ~((COMP_LOOP_acc_12_psp_sva[1:0]==2'b11) & (STAGE_VEC_LOOP_j_sva_9_0[1:0]==2'b11)
      & (fsm_output[2]) & (fsm_output[3]) & (fsm_output[6]) & (~ (fsm_output[5])));
  assign nand_449_nl = ~((operator_64_false_acc_cse_12_sva[3:0]==4'b1111) & (fsm_output[2])
      & (fsm_output[3]) & (~ (fsm_output[6])) & (fsm_output[5]));
  assign mux_2095_nl = MUX_s_1_2_2(nand_216_nl, nand_449_nl, fsm_output[4]);
  assign or_2282_nl = (fsm_output[4]) | (operator_64_false_acc_cse_sva[3:0]!=4'b1111)
      | (fsm_output[2]) | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign mux_2096_nl = MUX_s_1_2_2(mux_2095_nl, or_2282_nl, fsm_output[8]);
  assign or_2286_nl = (fsm_output[1]) | mux_2096_nl;
  assign mux_2101_nl = MUX_s_1_2_2(mux_2100_nl, or_2286_nl, fsm_output[9]);
  assign mux_2111_nl = MUX_s_1_2_2(mux_2110_nl, mux_2101_nl, fsm_output[7]);
  assign mux_2127_nl = MUX_s_1_2_2(mux_2126_nl, mux_2111_nl, fsm_output[0]);
  assign vec_rsc_0_15_i_wea_d_pff = ~ mux_2127_nl;
  assign and_531_nl = (COMP_LOOP_acc_cse_2_sva[3:0]==4'b1111) & (fsm_output[0]) &
      COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm & (fsm_output[3])
      & (fsm_output[6]) & (~ (fsm_output[5]));
  assign nor_570_nl = ~((COMP_LOOP_1_operator_64_false_acc_tmp[3:0]!=4'b1111) | (fsm_output[3])
      | (fsm_output[6]) | (fsm_output[5]));
  assign nor_571_nl = ~((STAGE_VEC_LOOP_j_sva_9_0[3:0]!=4'b1111) | (fsm_output[3])
      | (fsm_output[6]) | (fsm_output[5]));
  assign mux_2155_nl = MUX_s_1_2_2(nor_570_nl, nor_571_nl, fsm_output[0]);
  assign mux_2156_nl = MUX_s_1_2_2(and_531_nl, mux_2155_nl, fsm_output[4]);
  assign and_530_nl = (fsm_output[1]) & mux_2156_nl;
  assign and_532_nl = (fsm_output[1]) & (fsm_output[4]) & (fsm_output[0]) & (COMP_LOOP_acc_cse_10_sva[3:0]==4'b1111)
      & COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm & (~ (fsm_output[3]))
      & (~ (fsm_output[6])) & (~ (fsm_output[5]));
  assign mux_2157_nl = MUX_s_1_2_2(and_530_nl, and_532_nl, fsm_output[9]);
  assign nor_572_nl = ~((~((operator_64_false_acc_cse_14_sva[3:0]==4'b1111) & (fsm_output[9])
      & (~ (fsm_output[1])) & (fsm_output[4]) & (~ (fsm_output[0])))) | not_tmp_311);
  assign mux_2158_nl = MUX_s_1_2_2(mux_2157_nl, nor_572_nl, fsm_output[7]);
  assign or_2835_nl = (~((COMP_LOOP_acc_9_psp_sva[2:0]==3'b111) & (STAGE_VEC_LOOP_j_sva_9_0[0])
      & COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)) | not_tmp_311;
  assign nand_188_nl = ~((operator_64_false_acc_cse_7_sva[3:0]==4'b1111) & (fsm_output[3])
      & (fsm_output[6]) & (fsm_output[5]));
  assign mux_2151_nl = MUX_s_1_2_2(or_2835_nl, nand_188_nl, fsm_output[0]);
  assign or_2377_nl = (operator_64_false_acc_cse_6_sva[3:0]!=4'b1111) | (fsm_output[0])
      | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign mux_2152_nl = MUX_s_1_2_2(mux_2151_nl, or_2377_nl, fsm_output[4]);
  assign nor_573_nl = ~((fsm_output[1]) | mux_2152_nl);
  assign and_533_nl = operator_64_false_slc_operator_64_false_acc_1_60_itm & (fsm_output[0])
      & (COMP_LOOP_acc_cse_sva[3:0]==4'b1111) & (fsm_output[3]) & (fsm_output[6])
      & (fsm_output[5]);
  assign and_766_nl = (COMP_LOOP_acc_13_psp_sva[2:0]==3'b111) & (STAGE_VEC_LOOP_j_sva_9_0[0])
      & COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm & (~ (fsm_output[3]))
      & (~ (fsm_output[6])) & (fsm_output[5]);
  assign and_767_nl = (operator_64_false_acc_cse_15_sva[3:0]==4'b1111) & (~ (fsm_output[3]))
      & (~ (fsm_output[6])) & (fsm_output[5]);
  assign mux_2148_nl = MUX_s_1_2_2(and_766_nl, and_767_nl, fsm_output[0]);
  assign mux_2149_nl = MUX_s_1_2_2(and_533_nl, mux_2148_nl, fsm_output[4]);
  assign nor_576_nl = ~((operator_64_false_acc_cse_sva[3:0]!=4'b1111) | (fsm_output[4])
      | (fsm_output[0]) | not_tmp_311);
  assign mux_2150_nl = MUX_s_1_2_2(mux_2149_nl, nor_576_nl, fsm_output[1]);
  assign mux_2153_nl = MUX_s_1_2_2(nor_573_nl, mux_2150_nl, fsm_output[9]);
  assign nand_459_nl = ~((COMP_LOOP_acc_cse_8_sva[3:0]==4'b1111) & (~ (fsm_output[4]))
      & operator_64_false_slc_operator_64_false_acc_1_60_itm & (fsm_output[0]) &
      (~ (fsm_output[3])) & (~ (fsm_output[6])) & (fsm_output[5]));
  assign or_2365_nl = (operator_64_false_acc_cse_8_sva[3:0]!=4'b1111) | (fsm_output[0])
      | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign nand_190_nl = ~((STAGE_VEC_LOOP_j_sva_9_0[2:1]==2'b11) & (COMP_LOOP_acc_10_psp_sva[0])
      & (STAGE_VEC_LOOP_j_sva_9_0[0]) & COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm
      & (fsm_output[3]) & (fsm_output[6]) & (~ (fsm_output[5])));
  assign nand_191_nl = ~((operator_64_false_acc_cse_9_sva[3:0]==4'b1111) & (fsm_output[3])
      & (fsm_output[6]) & (~ (fsm_output[5])));
  assign mux_2145_nl = MUX_s_1_2_2(nand_190_nl, nand_191_nl, fsm_output[0]);
  assign mux_2146_nl = MUX_s_1_2_2(or_2365_nl, mux_2145_nl, fsm_output[4]);
  assign mux_2147_nl = MUX_s_1_2_2(nand_459_nl, mux_2146_nl, fsm_output[1]);
  assign nor_577_nl = ~((fsm_output[9]) | mux_2147_nl);
  assign mux_2154_nl = MUX_s_1_2_2(mux_2153_nl, nor_577_nl, fsm_output[7]);
  assign mux_2159_nl = MUX_s_1_2_2(mux_2158_nl, mux_2154_nl, fsm_output[8]);
  assign nor_578_nl = ~((operator_64_false_acc_cse_2_sva[3:0]!=4'b1111) | (fsm_output[1])
      | (fsm_output[4]) | (fsm_output[0]) | (~ (fsm_output[3])) | (~ (fsm_output[6]))
      | (fsm_output[5]));
  assign nand_192_nl = ~((COMP_LOOP_acc_11_psp_sva[2:0]==3'b111) & (STAGE_VEC_LOOP_j_sva_9_0[0])
      & COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm & (fsm_output[3])
      & (fsm_output[6]) & (~ (fsm_output[5])));
  assign nand_193_nl = ~((operator_64_false_acc_cse_11_sva[3:0]==4'b1111) & (fsm_output[3])
      & (fsm_output[6]) & (~ (fsm_output[5])));
  assign mux_2140_nl = MUX_s_1_2_2(nand_192_nl, nand_193_nl, fsm_output[0]);
  assign or_2357_nl = (fsm_output[0]) | (operator_64_false_acc_cse_10_sva[3:0]!=4'b1111)
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_2141_nl = MUX_s_1_2_2(mux_2140_nl, or_2357_nl, fsm_output[4]);
  assign nor_579_nl = ~((fsm_output[1]) | mux_2141_nl);
  assign mux_2142_nl = MUX_s_1_2_2(nor_578_nl, nor_579_nl, fsm_output[9]);
  assign nor_580_nl = ~((COMP_LOOP_acc_7_psp_sva[2:0]!=3'b111) | (~ (STAGE_VEC_LOOP_j_sva_9_0[0]))
      | (~ COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) | (fsm_output[3])
      | (fsm_output[6]) | (fsm_output[5]));
  assign nor_581_nl = ~((operator_64_false_acc_cse_3_sva[3:0]!=4'b1111) | (fsm_output[3])
      | (fsm_output[6]) | (fsm_output[5]));
  assign mux_2136_nl = MUX_s_1_2_2(nor_580_nl, nor_581_nl, fsm_output[0]);
  assign and_768_nl = operator_64_false_slc_operator_64_false_acc_1_60_itm & (COMP_LOOP_acc_cse_4_sva[3:0]==4'b1111)
      & (fsm_output[0]) & (fsm_output[3]) & (~ (fsm_output[6])) & (fsm_output[5]);
  assign mux_2137_nl = MUX_s_1_2_2(mux_2136_nl, and_768_nl, fsm_output[4]);
  assign nand_448_nl = ~((operator_64_false_acc_cse_4_sva[3:0]==4'b1111) & (fsm_output[6:5]==2'b01));
  assign mux_2133_nl = MUX_s_1_2_2(not_tmp_312, nand_448_nl, fsm_output[3]);
  assign nand_422_nl = ~((fsm_output[3]) & (operator_64_false_acc_cse_4_sva[3:0]==4'b1111)
      & (fsm_output[6:5]==2'b01));
  assign nand_197_nl = ~((STAGE_VEC_LOOP_j_sva_9_0[1]) & (COMP_LOOP_acc_8_psp_sva[1:0]==2'b11)
      & (STAGE_VEC_LOOP_j_sva_9_0[0]) & COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm);
  assign mux_2134_nl = MUX_s_1_2_2(mux_2133_nl, nand_422_nl, nand_197_nl);
  assign or_2347_nl = (~((operator_64_false_acc_cse_5_sva[3:0]==4'b1111) & (~ (fsm_output[3]))))
      | not_tmp_312;
  assign mux_2135_nl = MUX_s_1_2_2(mux_2134_nl, or_2347_nl, fsm_output[0]);
  assign and_534_nl = (fsm_output[4]) & (~ mux_2135_nl);
  assign mux_2138_nl = MUX_s_1_2_2(mux_2137_nl, and_534_nl, fsm_output[1]);
  assign nor_583_nl = ~((fsm_output[4]) | (~ operator_64_false_slc_operator_64_false_acc_1_60_itm)
      | (~ (fsm_output[0])) | (COMP_LOOP_acc_cse_12_sva[3:0]!=4'b1111) | (fsm_output[3])
      | (fsm_output[6]) | (fsm_output[5]));
  assign nor_584_nl = ~((operator_64_false_acc_cse_12_sva[3:0]!=4'b1111) | (fsm_output[0])
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5]));
  assign and_774_nl = (COMP_LOOP_acc_12_psp_sva[1:0]==2'b11) & (STAGE_VEC_LOOP_j_sva_9_0[1:0]==2'b11)
      & COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm & (fsm_output[3])
      & (~ (fsm_output[6])) & (fsm_output[5]);
  assign and_780_nl = (fsm_output[3]) & (operator_64_false_acc_cse_13_sva[3:0]==4'b1111)
      & (fsm_output[6:5]==2'b01);
  assign and_535_nl = (COMP_LOOP_acc_cse_14_sva[3:0]==4'b1111) & (fsm_output[6:5]==2'b11);
  assign and_791_nl = (operator_64_false_acc_cse_13_sva[3:0]==4'b1111) & (fsm_output[6:5]==2'b01);
  assign mux_2128_nl = MUX_s_1_2_2(and_535_nl, and_791_nl, fsm_output[3]);
  assign mux_2129_nl = MUX_s_1_2_2(and_780_nl, mux_2128_nl, COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm);
  assign mux_2130_nl = MUX_s_1_2_2(and_774_nl, mux_2129_nl, fsm_output[0]);
  assign mux_2131_nl = MUX_s_1_2_2(nor_584_nl, mux_2130_nl, fsm_output[4]);
  assign mux_2132_nl = MUX_s_1_2_2(nor_583_nl, mux_2131_nl, fsm_output[1]);
  assign mux_2139_nl = MUX_s_1_2_2(mux_2138_nl, mux_2132_nl, fsm_output[9]);
  assign mux_2143_nl = MUX_s_1_2_2(mux_2142_nl, mux_2139_nl, fsm_output[7]);
  assign and_792_nl = (COMP_LOOP_acc_cse_6_sva[3:0]==4'b1111) & (~ (fsm_output[7]))
      & (~ (fsm_output[9])) & (fsm_output[1]) & (~ (fsm_output[4])) & (fsm_output[0])
      & COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm & (fsm_output[3])
      & (~ (fsm_output[6])) & (fsm_output[5]);
  assign mux_2144_nl = MUX_s_1_2_2(mux_2143_nl, and_792_nl, fsm_output[8]);
  assign vec_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_2159_nl,
      mux_2144_nl, fsm_output[2]);
  assign or_tmp_2740 = ~((fsm_output[5]) & (fsm_output[3]) & (~ (fsm_output[8]))
      & (fsm_output[2]));
  assign or_2912_nl = (~ (fsm_output[5])) | (fsm_output[3]) | (~ (fsm_output[8]))
      | (fsm_output[2]);
  assign mux_2799_nl = MUX_s_1_2_2(or_2912_nl, or_tmp_2740, fsm_output[4]);
  assign or_2913_nl = (fsm_output[7]) | mux_2799_nl;
  assign or_2999_nl = (fsm_output[5]) | (fsm_output[3]) | (~ (fsm_output[8])) | (fsm_output[2]);
  assign mux_nl = MUX_s_1_2_2(or_tmp_2740, or_2999_nl, fsm_output[4]);
  assign nand_481_nl = ~((fsm_output[7]) & (~ mux_nl));
  assign mux_2800_nl = MUX_s_1_2_2(or_2913_nl, nand_481_nl, fsm_output[1]);
  assign or_tmp_2743 = (fsm_output[6]) | mux_2800_nl;
  assign or_2918_nl = (~ (fsm_output[3])) | (~ (fsm_output[8])) | (fsm_output[2]);
  assign or_2917_nl = (fsm_output[3]) | (fsm_output[8]) | (~ (fsm_output[2]));
  assign mux_tmp_2749 = MUX_s_1_2_2(or_2918_nl, or_2917_nl, fsm_output[5]);
  assign nand_tmp_150 = (fsm_output[7]) | (~ (fsm_output[4])) | mux_tmp_2749;
  assign and_dcpl_402 = (fsm_output==10'b0000000101);
  assign or_2929_cse = (fsm_output[6]) | (fsm_output[3]) | (fsm_output[9]) | (~ and_697_cse);
  assign or_2938_cse = (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[9])) |
      (fsm_output[0]) | (~ (fsm_output[2]));
  assign and_dcpl_418 = (~ (fsm_output[2])) & (fsm_output[1]) & (fsm_output[8]) &
      (fsm_output[0]) & (fsm_output[7]) & and_dcpl_95 & (fsm_output[5]) & (fsm_output[9])
      & (~ (fsm_output[4]));
  assign and_dcpl_419 = ~((fsm_output[9]) | (fsm_output[4]));
  assign and_dcpl_421 = (fsm_output[3]) & (~ (fsm_output[6])) & (fsm_output[5]);
  assign and_dcpl_423 = (fsm_output[0]) & (~ (fsm_output[7]));
  assign and_dcpl_424 = (~ (fsm_output[8])) & (fsm_output[2]);
  assign and_dcpl_427 = and_dcpl_424 & (fsm_output[1]) & and_dcpl_423 & and_dcpl_421
      & and_dcpl_419;
  assign and_dcpl_429 = and_711_cse & (fsm_output[5]);
  assign and_dcpl_431 = ~((fsm_output[0]) | (fsm_output[7]));
  assign and_dcpl_432 = ~((fsm_output[8]) | (fsm_output[2]));
  assign and_dcpl_433 = and_dcpl_432 & (~ (fsm_output[1]));
  assign and_dcpl_434 = and_dcpl_433 & and_dcpl_431;
  assign and_dcpl_435 = and_dcpl_434 & and_dcpl_429 & and_dcpl_419;
  assign and_dcpl_436 = (~ (fsm_output[9])) & (fsm_output[4]);
  assign and_dcpl_437 = and_711_cse & (~ (fsm_output[5]));
  assign and_dcpl_439 = (~ (fsm_output[0])) & (fsm_output[7]);
  assign and_dcpl_440 = and_dcpl_432 & (fsm_output[1]);
  assign and_dcpl_441 = and_dcpl_440 & and_dcpl_439;
  assign and_dcpl_442 = and_dcpl_441 & and_dcpl_437 & and_dcpl_436;
  assign and_dcpl_444 = and_dcpl_95 & (~ (fsm_output[5]));
  assign and_dcpl_445 = and_dcpl_444 & and_dcpl_436;
  assign and_dcpl_449 = (fsm_output[8]) & (~ (fsm_output[2])) & (fsm_output[1]) &
      and_dcpl_423 & and_dcpl_445;
  assign and_dcpl_451 = (fsm_output[8]) & (fsm_output[2]);
  assign and_dcpl_452 = and_dcpl_451 & (~ (fsm_output[1]));
  assign and_dcpl_453 = and_dcpl_452 & and_dcpl_431;
  assign and_dcpl_454 = and_dcpl_453 & and_dcpl_437 & and_dcpl_419;
  assign and_dcpl_456 = and_dcpl_451 & (fsm_output[1]);
  assign and_dcpl_457 = and_dcpl_456 & and_dcpl_439;
  assign and_dcpl_458 = and_dcpl_457 & and_dcpl_421 & and_dcpl_436;
  assign and_dcpl_462 = (fsm_output[0]) & (fsm_output[7]);
  assign and_dcpl_464 = and_dcpl_456 & and_dcpl_462 & (~ (fsm_output[3])) & (fsm_output[6])
      & (fsm_output[5]) & and_dcpl_436;
  assign and_dcpl_465 = (fsm_output[9]) & (fsm_output[4]);
  assign and_dcpl_466 = and_dcpl_95 & (fsm_output[5]);
  assign and_dcpl_468 = and_dcpl_434 & and_dcpl_466 & and_dcpl_465;
  assign and_dcpl_469 = (fsm_output[9]) & (~ (fsm_output[4]));
  assign and_dcpl_470 = and_dcpl_466 & and_dcpl_469;
  assign and_dcpl_471 = and_dcpl_441 & and_dcpl_470;
  assign and_dcpl_474 = and_dcpl_440 & and_dcpl_462 & and_dcpl_437 & and_dcpl_465;
  assign and_dcpl_476 = and_dcpl_453 & and_dcpl_444 & and_dcpl_465;
  assign and_dcpl_478 = and_dcpl_440 & and_dcpl_431 & and_dcpl_445;
  assign and_dcpl_481 = and_dcpl_433 & and_dcpl_462 & and_dcpl_466 & and_dcpl_419;
  assign and_dcpl_483 = and_dcpl_433 & and_dcpl_423;
  assign and_dcpl_484 = and_dcpl_483 & and_dcpl_429 & and_dcpl_469;
  assign and_dcpl_487 = and_dcpl_452 & and_dcpl_423 & and_dcpl_437 & and_dcpl_469;
  assign or_2955_cse = (fsm_output[6]) | (fsm_output[3]) | (fsm_output[9]) | (~ (fsm_output[0]))
      | (fsm_output[2]);
  assign mux_2829_cse = MUX_s_1_2_2(or_2938_cse, or_2955_cse, fsm_output[1]);
  assign mux_2830_cse = MUX_s_1_2_2(or_2929_cse, or_2938_cse, fsm_output[1]);
  assign or_2960_cse = (fsm_output[1]) | nand_176_cse;
  assign nand_484_nl = ~((fsm_output[7]) & (fsm_output[1]) & (fsm_output[6]) & (fsm_output[3])
      & mux_2326_cse);
  assign mux_2832_nl = MUX_s_1_2_2(or_2960_cse, mux_2830_cse, fsm_output[7]);
  assign mux_2833_nl = MUX_s_1_2_2(nand_484_nl, mux_2832_nl, fsm_output[4]);
  assign or_2958_nl = (fsm_output[4]) | (fsm_output[7]) | mux_2829_cse;
  assign mux_2834_nl = MUX_s_1_2_2(mux_2833_nl, or_2958_nl, fsm_output[5]);
  assign or_2952_nl = (~ (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[0])
      | (fsm_output[2]);
  assign or_2950_nl = (fsm_output[0]) | (fsm_output[2]);
  assign or_2949_nl = (~ (fsm_output[0])) | (fsm_output[2]);
  assign mux_2825_nl = MUX_s_1_2_2(or_2950_nl, or_2949_nl, fsm_output[9]);
  assign or_2951_nl = (fsm_output[3]) | mux_2825_nl;
  assign mux_2826_nl = MUX_s_1_2_2(or_2952_nl, or_2951_nl, fsm_output[6]);
  assign mux_2827_nl = MUX_s_1_2_2(mux_2826_nl, or_2929_cse, fsm_output[1]);
  assign or_2953_nl = (fsm_output[4]) | (fsm_output[7]) | mux_2827_nl;
  assign nand_479_nl = ~((fsm_output[7]) & (fsm_output[1]) & (fsm_output[6]) & (fsm_output[3])
      & (~ (fsm_output[9])) & (fsm_output[0]) & (~ (fsm_output[2])));
  assign or_2944_nl = (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[9])
      | (~ (fsm_output[0])) | (fsm_output[2]);
  assign or_2943_nl = (~ (fsm_output[6])) | (~ (fsm_output[3])) | (~ (fsm_output[9]))
      | (fsm_output[0]) | (fsm_output[2]);
  assign mux_2822_nl = MUX_s_1_2_2(or_2944_nl, or_2943_nl, fsm_output[1]);
  assign or_2942_nl = (~ (fsm_output[1])) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[9])
      | (fsm_output[0]) | (fsm_output[2]);
  assign mux_2823_nl = MUX_s_1_2_2(mux_2822_nl, or_2942_nl, fsm_output[7]);
  assign mux_2824_nl = MUX_s_1_2_2(nand_479_nl, mux_2823_nl, fsm_output[4]);
  assign mux_2828_nl = MUX_s_1_2_2(or_2953_nl, mux_2824_nl, fsm_output[5]);
  assign mux_2835_cse = MUX_s_1_2_2(mux_2834_nl, mux_2828_nl, fsm_output[8]);
  assign and_dcpl_489 = and_dcpl_452 & and_dcpl_439 & and_dcpl_470;
  assign and_dcpl_490 = and_dcpl_444 & and_dcpl_419;
  assign and_dcpl_491 = and_dcpl_424 & (~ (fsm_output[1]));
  assign and_dcpl_493 = and_dcpl_491 & and_dcpl_431 & and_dcpl_490;
  assign and_dcpl_495 = and_dcpl_491 & and_dcpl_423 & and_dcpl_490;
  assign and_dcpl_496 = and_dcpl_483 & and_dcpl_445;
  assign and_dcpl_498 = and_dcpl_457 & and_dcpl_444 & and_dcpl_469;
  assign and_dcpl_505 = nor_554_cse & (~ (fsm_output[8]));
  assign and_dcpl_507 = and_dcpl_505 & and_dcpl_423 & and_dcpl_490;
  assign and_dcpl_508 = (fsm_output[2:1]==2'b10);
  assign and_dcpl_509 = and_dcpl_508 & (~ (fsm_output[8]));
  assign and_dcpl_510 = and_dcpl_509 & and_dcpl_423;
  assign and_dcpl_511 = and_dcpl_510 & and_dcpl_490;
  assign and_920_cse = and_dcpl_509 & and_dcpl_431 & and_dcpl_444 & and_dcpl_436;
  assign nand_477_nl = ~((fsm_output[7]) & (fsm_output[4]) & (fsm_output[1]) & (fsm_output[6])
      & (fsm_output[3]) & mux_2332_cse);
  assign mux_2860_nl = MUX_s_1_2_2(or_2960_cse, mux_2829_cse, fsm_output[4]);
  assign or_2996_nl = (fsm_output[4]) | mux_2830_cse;
  assign mux_2861_nl = MUX_s_1_2_2(mux_2860_nl, or_2996_nl, fsm_output[7]);
  assign mux_2862_nl = MUX_s_1_2_2(nand_477_nl, mux_2861_nl, fsm_output[8]);
  assign nand_476_nl = ~((fsm_output[6]) & (fsm_output[3]) & mux_2332_cse);
  assign or_2989_nl = (fsm_output[6]) | (~ (fsm_output[3])) | (fsm_output[9]) | (~
      and_697_cse);
  assign mux_2853_nl = MUX_s_1_2_2(nand_476_nl, or_2989_nl, fsm_output[1]);
  assign or_2987_nl = (fsm_output[1]) | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[9]))
      | (fsm_output[0]) | (fsm_output[2]);
  assign mux_2854_nl = MUX_s_1_2_2(mux_2853_nl, or_2987_nl, fsm_output[4]);
  assign or_2984_nl = (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[9])) | (fsm_output[0])
      | (fsm_output[2]);
  assign mux_2851_nl = MUX_s_1_2_2(or_2955_cse, or_2984_nl, fsm_output[1]);
  assign or_2986_nl = (fsm_output[4]) | mux_2851_nl;
  assign mux_2855_nl = MUX_s_1_2_2(mux_2854_nl, or_2986_nl, fsm_output[7]);
  assign nor_1007_nl = ~((~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[0])
      | (~ (fsm_output[2])));
  assign nor_1008_nl = ~((fsm_output[3]) | (fsm_output[9]) | (~ and_697_cse));
  assign mux_2850_nl = MUX_s_1_2_2(nor_1007_nl, nor_1008_nl, fsm_output[6]);
  assign nand_475_nl = ~((fsm_output[7]) & (fsm_output[4]) & (fsm_output[1]) & mux_2850_nl);
  assign mux_2856_nl = MUX_s_1_2_2(mux_2855_nl, nand_475_nl, fsm_output[8]);
  assign mux_2863_itm = MUX_s_1_2_2(mux_2862_nl, mux_2856_nl, fsm_output[5]);
  assign and_925_cse = and_dcpl_510 & and_dcpl_437 & and_dcpl_419;
  assign and_dcpl_523 = (fsm_output[2]) & (fsm_output[1]) & (~ (fsm_output[8]));
  assign and_dcpl_525 = and_dcpl_523 & and_dcpl_439 & and_dcpl_490;
  assign and_dcpl_530 = and_dcpl_523 & and_dcpl_462;
  assign and_936_cse = and_dcpl_530 & (fsm_output[3]) & (~ (fsm_output[6])) & (fsm_output[5])
      & and_dcpl_436;
  assign and_dcpl_534 = and_dcpl_505 & and_dcpl_439;
  assign and_940_cse = and_dcpl_534 & and_dcpl_429 & and_dcpl_436;
  assign and_945_cse = nor_554_cse & (fsm_output[8]) & and_dcpl_423 & and_dcpl_466
      & and_dcpl_436;
  assign and_dcpl_543 = (~ (fsm_output[2])) & (fsm_output[1]) & (fsm_output[8]);
  assign and_dcpl_544 = and_dcpl_543 & and_dcpl_431;
  assign and_950_cse = and_dcpl_544 & and_dcpl_429 & and_dcpl_419;
  assign and_953_cse = and_dcpl_543 & and_dcpl_462 & and_dcpl_466 & and_dcpl_419;
  assign and_957_cse = and_dcpl_508 & (fsm_output[8]) & and_dcpl_439 & and_dcpl_437
      & and_dcpl_436;
  assign and_960_cse = and_dcpl_510 & and_dcpl_444 & and_dcpl_465;
  assign and_964_cse = and_dcpl_523 & and_dcpl_431 & and_dcpl_437 & and_dcpl_469;
  assign and_966_cse = and_dcpl_530 & and_dcpl_444 & and_dcpl_469;
  assign and_970_cse = and_dcpl_534 & (~ (fsm_output[3])) & (fsm_output[6]) & (~
      (fsm_output[5])) & and_dcpl_469;
  assign and_973_cse = and_dcpl_505 & and_dcpl_462 & and_dcpl_429 & and_dcpl_465;
  assign and_975_cse = and_dcpl_544 & and_dcpl_466 & and_dcpl_465;
  assign and_978_cse = and_dcpl_543 & and_dcpl_423 & and_dcpl_429 & and_dcpl_469;
  assign and_dcpl_582 = and_dcpl_432 & (fsm_output[1]) & (~ (fsm_output[0])) & (~
      (fsm_output[7])) & nor_1039_cse & (~ (fsm_output[9])) & (fsm_output[4]);
  assign and_dcpl_584 = nor_1039_cse & (~ (fsm_output[9])) & (~ (fsm_output[4]));
  assign and_dcpl_589 = and_dcpl_451 & (~ (fsm_output[1])) & (fsm_output[0]) & (fsm_output[7])
      & and_dcpl_584;
  assign and_dcpl_593 = and_dcpl_432 & (~ (fsm_output[1])) & (fsm_output[0]) & (~
      (fsm_output[7])) & and_dcpl_584;
  assign and_dcpl_599 = and_dcpl_451 & (fsm_output[1]) & (~ (fsm_output[0])) & (fsm_output[7])
      & nor_1039_cse & (fsm_output[9]) & (~ (fsm_output[4]));
  assign and_dcpl_621 = and_dcpl_523 & and_dcpl_439 & and_dcpl_444 & and_dcpl_419;
  assign mux_tmp_2812 = MUX_s_1_2_2(and_694_cse, or_204_cse, fsm_output[3]);
  assign mux_tmp_2813 = MUX_s_1_2_2((~ or_204_cse), or_204_cse, fsm_output[3]);
  assign mux_tmp_2815 = MUX_s_1_2_2((~ or_204_cse), (fsm_output[6]), fsm_output[3]);
  assign mux_tmp_2823 = MUX_s_1_2_2((~ (fsm_output[6])), and_694_cse, fsm_output[3]);
  assign mux_tmp_2824 = MUX_s_1_2_2((~ and_694_cse), and_694_cse, fsm_output[3]);
  assign operator_64_false_or_120_itm = and_dcpl_427 | and_dcpl_435 | and_dcpl_442
      | and_dcpl_449 | and_dcpl_454 | and_dcpl_458 | and_dcpl_464 | and_dcpl_468
      | and_dcpl_471 | and_dcpl_474 | and_dcpl_476 | and_dcpl_496 | and_dcpl_498;
  assign operator_64_false_or_121_cse = (~ mux_2835_cse) | and_dcpl_495;
  assign operator_64_false_operator_64_false_or_1_cse = (~(and_dcpl_427 | and_dcpl_435
      | and_dcpl_442 | and_dcpl_449 | and_dcpl_454 | and_dcpl_458 | and_dcpl_464
      | and_dcpl_468 | and_dcpl_471 | and_dcpl_474 | and_dcpl_476 | and_dcpl_478
      | and_dcpl_481 | and_dcpl_484 | and_dcpl_487 | (~ mux_2835_cse) | and_dcpl_493
      | and_dcpl_495 | and_dcpl_496 | and_dcpl_498)) | and_dcpl_489;
  always @(posedge clk) begin
    if ( ~ not_tmp_266 ) begin
      p_sva <= p_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( ~ not_tmp_266 ) begin
      r_sva <= r_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_vec_rsc_triosy_0_15_obj_ld_cse <= 1'b0;
      reg_ensig_cgo_cse <= 1'b0;
      COMP_LOOP_COMP_LOOP_nor_1_itm <= 1'b0;
      COMP_LOOP_nor_12_itm <= 1'b0;
      COMP_LOOP_nor_14_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_19_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_20_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_21_itm <= 1'b0;
      COMP_LOOP_nor_17_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_23_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_24_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_25_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_26_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_27_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_28_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_29_itm <= 1'b0;
    end
    else begin
      reg_vec_rsc_triosy_0_15_obj_ld_cse <= and_dcpl_199 & and_dcpl_159 & (~ (fsm_output[0]))
          & (fsm_output[7]) & (fsm_output[8]) & (fsm_output[9]) & (z_out_2[4]);
      reg_ensig_cgo_cse <= ~ mux_2240_itm;
      COMP_LOOP_COMP_LOOP_nor_1_itm <= ~((COMP_LOOP_1_operator_64_false_acc_tmp[3:0]!=4'b0000));
      COMP_LOOP_nor_12_itm <= ~((COMP_LOOP_1_operator_64_false_acc_tmp[3]) | (COMP_LOOP_1_operator_64_false_acc_tmp[2])
          | (COMP_LOOP_1_operator_64_false_acc_tmp[0]));
      COMP_LOOP_nor_14_itm <= ~((COMP_LOOP_1_operator_64_false_acc_tmp[3]) | (COMP_LOOP_1_operator_64_false_acc_tmp[1])
          | (COMP_LOOP_1_operator_64_false_acc_tmp[0]));
      COMP_LOOP_COMP_LOOP_and_19_itm <= (COMP_LOOP_1_operator_64_false_acc_tmp[3:0]==4'b0101);
      COMP_LOOP_COMP_LOOP_and_20_itm <= (COMP_LOOP_1_operator_64_false_acc_tmp[3:0]==4'b0110);
      COMP_LOOP_COMP_LOOP_and_21_itm <= (COMP_LOOP_1_operator_64_false_acc_tmp[3:0]==4'b0111);
      COMP_LOOP_nor_17_itm <= ~((COMP_LOOP_1_operator_64_false_acc_tmp[2:0]!=3'b000));
      COMP_LOOP_COMP_LOOP_and_23_itm <= (COMP_LOOP_1_operator_64_false_acc_tmp[3:0]==4'b1001);
      COMP_LOOP_COMP_LOOP_and_24_itm <= (COMP_LOOP_1_operator_64_false_acc_tmp[3:0]==4'b1010);
      COMP_LOOP_COMP_LOOP_and_25_itm <= (COMP_LOOP_1_operator_64_false_acc_tmp[3:0]==4'b1011);
      COMP_LOOP_COMP_LOOP_and_26_itm <= (COMP_LOOP_1_operator_64_false_acc_tmp[3:0]==4'b1100);
      COMP_LOOP_COMP_LOOP_and_27_itm <= (COMP_LOOP_1_operator_64_false_acc_tmp[3:0]==4'b1101);
      COMP_LOOP_COMP_LOOP_and_28_itm <= (COMP_LOOP_1_operator_64_false_acc_tmp[3:0]==4'b1110);
      COMP_LOOP_COMP_LOOP_and_29_itm <= (COMP_LOOP_1_operator_64_false_acc_tmp[3:0]==4'b1111);
    end
  end
  always @(posedge clk) begin
    reg_COMP_LOOP_1_modulo_dev_cmp_m_rsc_dat_cse <= p_sva;
    modExp_dev_while_rem_cmp_a <= MUX_v_64_2_2(COMP_LOOP_10_modExp_dev_1_while_mul_mut,
        z_out, mux_2323_nl);
    STAGE_MAIN_LOOP_div_cmp_a <= MUX_v_64_2_2(z_out_3, COMP_LOOP_10_modExp_dev_1_while_mul_mut,
        and_dcpl_293);
    STAGE_MAIN_LOOP_div_cmp_b <= MUX_v_10_2_2(STAGE_MAIN_LOOP_lshift_psp_1_sva_mx0w0,
        STAGE_MAIN_LOOP_lshift_psp_1_sva, and_dcpl_293);
  end
  always @(posedge clk) begin
    if ( mux_2339_nl | and_dcpl_295 ) begin
      STAGE_MAIN_LOOP_acc_1_psp_sva <= MUX_v_4_2_2(4'b1010, (COMP_LOOP_slc_acc_3_12_1_slc[3:0]),
          and_dcpl_295);
    end
  end
  always @(posedge clk) begin
    if ( MUX_s_1_2_2(nor_548_nl, and_tmp_24, fsm_output[9]) ) begin
      STAGE_MAIN_LOOP_lshift_psp_1_sva <= STAGE_MAIN_LOOP_lshift_psp_1_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( and_dcpl_295 | and_dcpl_290 | not_tmp_597 | (~ mux_2336_itm) | COMP_LOOP_10_modExp_dev_1_while_mul_mut_mx0c4
        | COMP_LOOP_10_modExp_dev_1_while_mul_mut_mx0c5 ) begin
      COMP_LOOP_10_modExp_dev_1_while_mul_mut <= MUX1HOT_v_64_4_2(z_out_3, z_out,
          64'b0000000000000000000000000000000000000000000000000000000000000001, modExp_dev_while_rem_cmp_z,
          {and_dcpl_295 , operator_64_false_or_2_nl , not_tmp_597 , COMP_LOOP_10_modExp_dev_1_while_mul_mut_mx0c4});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      STAGE_VEC_LOOP_j_sva_9_0 <= 10'b0000000000;
    end
    else if ( (and_dcpl_95 & (~ (fsm_output[1])) & ((fsm_output[2]) ^ (fsm_output[4]))
        & (~ (fsm_output[5])) & (~ (fsm_output[0])) & (~ (fsm_output[7])) & and_dcpl)
        | STAGE_VEC_LOOP_j_sva_9_0_mx0c1 ) begin
      STAGE_VEC_LOOP_j_sva_9_0 <= MUX_v_10_2_2(10'b0000000000, (z_out_1[9:0]), STAGE_VEC_LOOP_j_sva_9_0_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( mux_2427_nl | and_330_rgt ) begin
      modExp_dev_result_sva <= MUX_v_64_2_2(64'b0000000000000000000000000000000000000000000000000000000000000001,
          modExp_dev_while_rem_cmp_z, and_330_rgt);
    end
  end
  always @(posedge clk) begin
    if ( MUX_s_1_2_2(mux_2475_nl, mux_2450_nl, fsm_output[9]) ) begin
      tmp_10_lpi_4_dfm <= MUX1HOT_v_64_18_2(STAGE_MAIN_LOOP_div_cmp_z, z_out_3, vec_rsc_0_0_i_qa_d,
          vec_rsc_0_1_i_qa_d, vec_rsc_0_2_i_qa_d, vec_rsc_0_3_i_qa_d, vec_rsc_0_4_i_qa_d,
          vec_rsc_0_5_i_qa_d, vec_rsc_0_6_i_qa_d, vec_rsc_0_7_i_qa_d, vec_rsc_0_8_i_qa_d,
          vec_rsc_0_9_i_qa_d, vec_rsc_0_10_i_qa_d, vec_rsc_0_11_i_qa_d, vec_rsc_0_12_i_qa_d,
          vec_rsc_0_13_i_qa_d, vec_rsc_0_14_i_qa_d, vec_rsc_0_15_i_qa_d, {and_331_nl
          , and_dcpl_290 , COMP_LOOP_or_2_nl , COMP_LOOP_or_3_nl , COMP_LOOP_or_4_nl
          , COMP_LOOP_or_5_nl , COMP_LOOP_or_6_nl , COMP_LOOP_or_7_nl , COMP_LOOP_or_8_nl
          , COMP_LOOP_or_9_nl , COMP_LOOP_or_10_nl , COMP_LOOP_or_11_nl , COMP_LOOP_or_12_nl
          , COMP_LOOP_or_13_nl , COMP_LOOP_or_14_nl , COMP_LOOP_or_15_nl , COMP_LOOP_or_16_nl
          , COMP_LOOP_or_17_nl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm <= 1'b0;
    end
    else if ( and_dcpl_290 | and_dcpl_98 | (~ mux_2336_itm) | COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c3
        | COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c4 |
        COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c5 | COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c6
        | COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c7 |
        COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c8 | COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c9
        | COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c10
        | COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c11
        | COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c12
        | COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c13
        | and_dcpl_345 ) begin
      COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm <= MUX1HOT_s_1_4_2((~
          (z_out_2[64])), COMP_LOOP_COMP_LOOP_and_17_nl, (z_out_2[63]), (~ (z_out_2[63])),
          {modExp_dev_while_or_nl , and_dcpl_98 , modExp_dev_while_or_1_nl , and_dcpl_345});
    end
  end
  always @(posedge clk) begin
    if ( mux_2864_nl & nor_1039_cse ) begin
      COMP_LOOP_k_9_4_sva_4_0 <= MUX_v_5_2_2(5'b00000, (COMP_LOOP_slc_acc_3_12_1_slc[4:0]),
          nand_486_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      operator_64_false_acc_cse_1_sva <= 10'b0000000000;
    end
    else if ( ~ or_dcpl_72 ) begin
      operator_64_false_acc_cse_1_sva <= COMP_LOOP_1_operator_64_false_acc_tmp;
    end
  end
  always @(posedge clk) begin
    if ( and_dcpl_98 | (~ mux_2545_itm) ) begin
      COMP_LOOP_acc_psp_sva <= MUX_v_6_2_2(({2'b00 , operator_64_false_or_2_nl_1}),
          (z_out_1[5:0]), mux_2545_itm);
    end
  end
  always @(posedge clk) begin
    if ( ~ or_dcpl_72 ) begin
      operator_64_false_1_slc_operator_64_false_1_acc_5_itm <= readslicef_6_1_5(operator_64_false_1_acc_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_nor_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_244_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_62_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_185_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_64_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_65_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_66_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_6_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_68_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_69_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_70_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_10_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_72_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_12_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_13_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_14_itm <= 1'b0;
    end
    else if ( mux_2586_itm ) begin
      COMP_LOOP_COMP_LOOP_nor_itm <= ~((STAGE_VEC_LOOP_j_sva_9_0[3:0]!=4'b0000));
      COMP_LOOP_COMP_LOOP_and_244_itm <= (COMP_LOOP_acc_8_psp_sva_1[0]) & (STAGE_VEC_LOOP_j_sva_9_0[0])
          & (~((COMP_LOOP_acc_8_psp_sva_1[1]) | (STAGE_VEC_LOOP_j_sva_9_0[1])));
      COMP_LOOP_COMP_LOOP_and_62_itm <= (COMP_LOOP_acc_cse_2_sva_1[3:0]==4'b0011);
      COMP_LOOP_COMP_LOOP_and_185_itm <= (COMP_LOOP_acc_cse_4_sva_1[3:0]==4'b0110);
      COMP_LOOP_COMP_LOOP_and_64_itm <= (COMP_LOOP_acc_cse_2_sva_1[3:0]==4'b0101);
      COMP_LOOP_COMP_LOOP_and_65_itm <= (COMP_LOOP_acc_cse_2_sva_1[3:0]==4'b0110);
      COMP_LOOP_COMP_LOOP_and_66_itm <= (COMP_LOOP_acc_cse_2_sva_1[3:0]==4'b0111);
      COMP_LOOP_COMP_LOOP_and_6_itm <= (STAGE_VEC_LOOP_j_sva_9_0[3:0]==4'b0111);
      COMP_LOOP_COMP_LOOP_and_68_itm <= (COMP_LOOP_acc_cse_2_sva_1[3:0]==4'b1001);
      COMP_LOOP_COMP_LOOP_and_69_itm <= (COMP_LOOP_acc_cse_2_sva_1[3:0]==4'b1010);
      COMP_LOOP_COMP_LOOP_and_70_itm <= (COMP_LOOP_acc_cse_2_sva_1[3:0]==4'b1011);
      COMP_LOOP_COMP_LOOP_and_10_itm <= (STAGE_VEC_LOOP_j_sva_9_0[3:0]==4'b1011);
      COMP_LOOP_COMP_LOOP_and_72_itm <= (COMP_LOOP_acc_cse_2_sva_1[3:0]==4'b1101);
      COMP_LOOP_COMP_LOOP_and_12_itm <= (STAGE_VEC_LOOP_j_sva_9_0[3:0]==4'b1101);
      COMP_LOOP_COMP_LOOP_and_13_itm <= (STAGE_VEC_LOOP_j_sva_9_0[3:0]==4'b1110);
      COMP_LOOP_COMP_LOOP_and_14_itm <= (STAGE_VEC_LOOP_j_sva_9_0[3:0]==4'b1111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_8_psp_sva <= 8'b00000000;
    end
    else if ( mux_2590_nl | (fsm_output[9]) ) begin
      COMP_LOOP_acc_8_psp_sva <= COMP_LOOP_acc_8_psp_sva_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_cse_4_sva <= 10'b0000000000;
    end
    else if ( ~(mux_2592_nl & and_dcpl) ) begin
      COMP_LOOP_acc_cse_4_sva <= COMP_LOOP_acc_cse_4_sva_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_cse_2_sva <= 10'b0000000000;
    end
    else if ( ~((~ mux_2599_nl) & nor_813_cse) ) begin
      COMP_LOOP_acc_cse_2_sva <= COMP_LOOP_acc_cse_2_sva_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      operator_64_false_acc_cse_2_sva <= 10'b0000000000;
    end
    else if ( ~(mux_2601_nl & and_dcpl) ) begin
      operator_64_false_acc_cse_2_sva <= operator_64_false_acc_cse_2_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_nor_5_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_354 ) begin
      COMP_LOOP_COMP_LOOP_nor_5_itm <= ~((operator_64_false_acc_cse_2_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_51_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_354 ) begin
      COMP_LOOP_nor_51_itm <= ~((operator_64_false_acc_cse_2_sva_mx0w0[3:1]!=3'b000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_52_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_354 ) begin
      COMP_LOOP_nor_52_itm <= ~((operator_64_false_acc_cse_2_sva_mx0w0[3]) | (operator_64_false_acc_cse_2_sva_mx0w0[2])
          | (operator_64_false_acc_cse_2_sva_mx0w0[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_77_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_354 ) begin
      COMP_LOOP_COMP_LOOP_and_77_itm <= (operator_64_false_acc_cse_2_sva_mx0w0[3:0]==4'b0011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_54_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_354 ) begin
      COMP_LOOP_nor_54_itm <= ~((operator_64_false_acc_cse_2_sva_mx0w0[3]) | (operator_64_false_acc_cse_2_sva_mx0w0[1])
          | (operator_64_false_acc_cse_2_sva_mx0w0[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_79_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_354 ) begin
      COMP_LOOP_COMP_LOOP_and_79_itm <= (operator_64_false_acc_cse_2_sva_mx0w0[3:0]==4'b0101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_80_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_354 ) begin
      COMP_LOOP_COMP_LOOP_and_80_itm <= (operator_64_false_acc_cse_2_sva_mx0w0[3:0]==4'b0110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_81_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_354 ) begin
      COMP_LOOP_COMP_LOOP_and_81_itm <= (operator_64_false_acc_cse_2_sva_mx0w0[3:0]==4'b0111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_57_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_354 ) begin
      COMP_LOOP_nor_57_itm <= ~((operator_64_false_acc_cse_2_sva_mx0w0[2:0]!=3'b000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_83_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_354 ) begin
      COMP_LOOP_COMP_LOOP_and_83_itm <= (operator_64_false_acc_cse_2_sva_mx0w0[3:0]==4'b1001);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_84_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_354 ) begin
      COMP_LOOP_COMP_LOOP_and_84_itm <= (operator_64_false_acc_cse_2_sva_mx0w0[3:0]==4'b1010);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_85_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_354 ) begin
      COMP_LOOP_COMP_LOOP_and_85_itm <= (operator_64_false_acc_cse_2_sva_mx0w0[3:0]==4'b1011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_86_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_354 ) begin
      COMP_LOOP_COMP_LOOP_and_86_itm <= (operator_64_false_acc_cse_2_sva_mx0w0[3:0]==4'b1100);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_87_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_354 ) begin
      COMP_LOOP_COMP_LOOP_and_87_itm <= (operator_64_false_acc_cse_2_sva_mx0w0[3:0]==4'b1101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_88_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_354 ) begin
      COMP_LOOP_COMP_LOOP_and_88_itm <= (operator_64_false_acc_cse_2_sva_mx0w0[3:0]==4'b1110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_89_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_354 ) begin
      COMP_LOOP_COMP_LOOP_and_89_itm <= (operator_64_false_acc_cse_2_sva_mx0w0[3:0]==4'b1111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_7_psp_sva <= 9'b000000000;
    end
    else if ( ~((mux_tmp_2538 ^ (fsm_output[7])) & and_dcpl) ) begin
      COMP_LOOP_acc_7_psp_sva <= nl_COMP_LOOP_acc_7_psp_sva[8:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      operator_64_false_acc_cse_3_sva <= 10'b0000000000;
    end
    else if ( ~(mux_2612_nl & and_dcpl) ) begin
      operator_64_false_acc_cse_3_sva <= operator_64_false_acc_cse_3_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_nor_9_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_357 ) begin
      COMP_LOOP_COMP_LOOP_nor_9_itm <= ~((operator_64_false_acc_cse_3_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_91_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_357 ) begin
      COMP_LOOP_nor_91_itm <= ~((operator_64_false_acc_cse_3_sva_mx0w0[3:1]!=3'b000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_92_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_357 ) begin
      COMP_LOOP_nor_92_itm <= ~((operator_64_false_acc_cse_3_sva_mx0w0[3]) | (operator_64_false_acc_cse_3_sva_mx0w0[2])
          | (operator_64_false_acc_cse_3_sva_mx0w0[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_137_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_357 ) begin
      COMP_LOOP_COMP_LOOP_and_137_itm <= (operator_64_false_acc_cse_3_sva_mx0w0[3:0]==4'b0011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_94_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_357 ) begin
      COMP_LOOP_nor_94_itm <= ~((operator_64_false_acc_cse_3_sva_mx0w0[3]) | (operator_64_false_acc_cse_3_sva_mx0w0[1])
          | (operator_64_false_acc_cse_3_sva_mx0w0[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_139_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_357 ) begin
      COMP_LOOP_COMP_LOOP_and_139_itm <= (operator_64_false_acc_cse_3_sva_mx0w0[3:0]==4'b0101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_140_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_357 ) begin
      COMP_LOOP_COMP_LOOP_and_140_itm <= (operator_64_false_acc_cse_3_sva_mx0w0[3:0]==4'b0110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_141_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_357 ) begin
      COMP_LOOP_COMP_LOOP_and_141_itm <= (operator_64_false_acc_cse_3_sva_mx0w0[3:0]==4'b0111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_97_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_357 ) begin
      COMP_LOOP_nor_97_itm <= ~((operator_64_false_acc_cse_3_sva_mx0w0[2:0]!=3'b000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_143_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_357 ) begin
      COMP_LOOP_COMP_LOOP_and_143_itm <= (operator_64_false_acc_cse_3_sva_mx0w0[3:0]==4'b1001);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_144_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_357 ) begin
      COMP_LOOP_COMP_LOOP_and_144_itm <= (operator_64_false_acc_cse_3_sva_mx0w0[3:0]==4'b1010);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_145_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_357 ) begin
      COMP_LOOP_COMP_LOOP_and_145_itm <= (operator_64_false_acc_cse_3_sva_mx0w0[3:0]==4'b1011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_146_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_357 ) begin
      COMP_LOOP_COMP_LOOP_and_146_itm <= (operator_64_false_acc_cse_3_sva_mx0w0[3:0]==4'b1100);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_147_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_357 ) begin
      COMP_LOOP_COMP_LOOP_and_147_itm <= (operator_64_false_acc_cse_3_sva_mx0w0[3:0]==4'b1101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_148_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_357 ) begin
      COMP_LOOP_COMP_LOOP_and_148_itm <= (operator_64_false_acc_cse_3_sva_mx0w0[3:0]==4'b1110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_149_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_357 ) begin
      COMP_LOOP_COMP_LOOP_and_149_itm <= (operator_64_false_acc_cse_3_sva_mx0w0[3:0]==4'b1111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      operator_64_false_acc_cse_4_sva <= 10'b0000000000;
    end
    else if ( ~(mux_2616_nl & and_dcpl) ) begin
      operator_64_false_acc_cse_4_sva <= operator_64_false_acc_cse_4_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_nor_13_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_359 ) begin
      COMP_LOOP_COMP_LOOP_nor_13_itm <= ~((operator_64_false_acc_cse_4_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_131_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_359 ) begin
      COMP_LOOP_nor_131_itm <= ~((operator_64_false_acc_cse_4_sva_mx0w0[3:1]!=3'b000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_132_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_359 ) begin
      COMP_LOOP_nor_132_itm <= ~((operator_64_false_acc_cse_4_sva_mx0w0[3]) | (operator_64_false_acc_cse_4_sva_mx0w0[2])
          | (operator_64_false_acc_cse_4_sva_mx0w0[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_197_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_359 ) begin
      COMP_LOOP_COMP_LOOP_and_197_itm <= (operator_64_false_acc_cse_4_sva_mx0w0[3:0]==4'b0011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_134_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_359 ) begin
      COMP_LOOP_nor_134_itm <= ~((operator_64_false_acc_cse_4_sva_mx0w0[3]) | (operator_64_false_acc_cse_4_sva_mx0w0[1])
          | (operator_64_false_acc_cse_4_sva_mx0w0[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_199_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_359 ) begin
      COMP_LOOP_COMP_LOOP_and_199_itm <= (operator_64_false_acc_cse_4_sva_mx0w0[3:0]==4'b0101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_200_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_359 ) begin
      COMP_LOOP_COMP_LOOP_and_200_itm <= (operator_64_false_acc_cse_4_sva_mx0w0[3:0]==4'b0110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_201_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_359 ) begin
      COMP_LOOP_COMP_LOOP_and_201_itm <= (operator_64_false_acc_cse_4_sva_mx0w0[3:0]==4'b0111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_137_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_359 ) begin
      COMP_LOOP_nor_137_itm <= ~((operator_64_false_acc_cse_4_sva_mx0w0[2:0]!=3'b000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_203_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_359 ) begin
      COMP_LOOP_COMP_LOOP_and_203_itm <= (operator_64_false_acc_cse_4_sva_mx0w0[3:0]==4'b1001);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_204_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_359 ) begin
      COMP_LOOP_COMP_LOOP_and_204_itm <= (operator_64_false_acc_cse_4_sva_mx0w0[3:0]==4'b1010);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_205_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_359 ) begin
      COMP_LOOP_COMP_LOOP_and_205_itm <= (operator_64_false_acc_cse_4_sva_mx0w0[3:0]==4'b1011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_206_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_359 ) begin
      COMP_LOOP_COMP_LOOP_and_206_itm <= (operator_64_false_acc_cse_4_sva_mx0w0[3:0]==4'b1100);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_207_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_359 ) begin
      COMP_LOOP_COMP_LOOP_and_207_itm <= (operator_64_false_acc_cse_4_sva_mx0w0[3:0]==4'b1101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_208_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_359 ) begin
      COMP_LOOP_COMP_LOOP_and_208_itm <= (operator_64_false_acc_cse_4_sva_mx0w0[3:0]==4'b1110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_209_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_359 ) begin
      COMP_LOOP_COMP_LOOP_and_209_itm <= (operator_64_false_acc_cse_4_sva_mx0w0[3:0]==4'b1111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      operator_64_false_acc_cse_5_sva <= 10'b0000000000;
    end
    else if ( mux_2621_nl | (fsm_output[9]) ) begin
      operator_64_false_acc_cse_5_sva <= operator_64_false_acc_cse_5_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_nor_17_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_361 ) begin
      COMP_LOOP_COMP_LOOP_nor_17_itm <= ~((operator_64_false_acc_cse_5_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_171_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_361 ) begin
      COMP_LOOP_nor_171_itm <= ~((operator_64_false_acc_cse_5_sva_mx0w0[3:1]!=3'b000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_172_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_361 ) begin
      COMP_LOOP_nor_172_itm <= ~((operator_64_false_acc_cse_5_sva_mx0w0[3]) | (operator_64_false_acc_cse_5_sva_mx0w0[2])
          | (operator_64_false_acc_cse_5_sva_mx0w0[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_257_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_361 ) begin
      COMP_LOOP_COMP_LOOP_and_257_itm <= (operator_64_false_acc_cse_5_sva_mx0w0[3:0]==4'b0011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_174_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_361 ) begin
      COMP_LOOP_nor_174_itm <= ~((operator_64_false_acc_cse_5_sva_mx0w0[3]) | (operator_64_false_acc_cse_5_sva_mx0w0[1])
          | (operator_64_false_acc_cse_5_sva_mx0w0[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_259_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_361 ) begin
      COMP_LOOP_COMP_LOOP_and_259_itm <= (operator_64_false_acc_cse_5_sva_mx0w0[3:0]==4'b0101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_260_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_361 ) begin
      COMP_LOOP_COMP_LOOP_and_260_itm <= (operator_64_false_acc_cse_5_sva_mx0w0[3:0]==4'b0110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_261_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_361 ) begin
      COMP_LOOP_COMP_LOOP_and_261_itm <= (operator_64_false_acc_cse_5_sva_mx0w0[3:0]==4'b0111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_177_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_361 ) begin
      COMP_LOOP_nor_177_itm <= ~((operator_64_false_acc_cse_5_sva_mx0w0[2:0]!=3'b000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_263_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_361 ) begin
      COMP_LOOP_COMP_LOOP_and_263_itm <= (operator_64_false_acc_cse_5_sva_mx0w0[3:0]==4'b1001);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_264_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_361 ) begin
      COMP_LOOP_COMP_LOOP_and_264_itm <= (operator_64_false_acc_cse_5_sva_mx0w0[3:0]==4'b1010);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_265_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_361 ) begin
      COMP_LOOP_COMP_LOOP_and_265_itm <= (operator_64_false_acc_cse_5_sva_mx0w0[3:0]==4'b1011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_266_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_361 ) begin
      COMP_LOOP_COMP_LOOP_and_266_itm <= (operator_64_false_acc_cse_5_sva_mx0w0[3:0]==4'b1100);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_267_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_361 ) begin
      COMP_LOOP_COMP_LOOP_and_267_itm <= (operator_64_false_acc_cse_5_sva_mx0w0[3:0]==4'b1101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_268_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_361 ) begin
      COMP_LOOP_COMP_LOOP_and_268_itm <= (operator_64_false_acc_cse_5_sva_mx0w0[3:0]==4'b1110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_269_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_361 ) begin
      COMP_LOOP_COMP_LOOP_and_269_itm <= (operator_64_false_acc_cse_5_sva_mx0w0[3:0]==4'b1111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_cse_6_sva <= 10'b0000000000;
    end
    else if ( mux_2624_nl | (fsm_output[9]) ) begin
      COMP_LOOP_acc_cse_6_sva <= COMP_LOOP_slc_acc_3_12_1_slc[9:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      operator_64_false_acc_cse_6_sva <= 10'b0000000000;
    end
    else if ( mux_2633_nl | (fsm_output[9]) ) begin
      operator_64_false_acc_cse_6_sva <= operator_64_false_acc_cse_6_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_nor_21_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_364 ) begin
      COMP_LOOP_COMP_LOOP_nor_21_itm <= ~((operator_64_false_acc_cse_6_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_211_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_364 ) begin
      COMP_LOOP_nor_211_itm <= ~((operator_64_false_acc_cse_6_sva_mx0w0[3:1]!=3'b000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_212_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_364 ) begin
      COMP_LOOP_nor_212_itm <= ~((operator_64_false_acc_cse_6_sva_mx0w0[3]) | (operator_64_false_acc_cse_6_sva_mx0w0[2])
          | (operator_64_false_acc_cse_6_sva_mx0w0[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_317_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_364 ) begin
      COMP_LOOP_COMP_LOOP_and_317_itm <= (operator_64_false_acc_cse_6_sva_mx0w0[3:0]==4'b0011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_214_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_364 ) begin
      COMP_LOOP_nor_214_itm <= ~((operator_64_false_acc_cse_6_sva_mx0w0[3]) | (operator_64_false_acc_cse_6_sva_mx0w0[1])
          | (operator_64_false_acc_cse_6_sva_mx0w0[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_319_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_364 ) begin
      COMP_LOOP_COMP_LOOP_and_319_itm <= (operator_64_false_acc_cse_6_sva_mx0w0[3:0]==4'b0101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_320_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_364 ) begin
      COMP_LOOP_COMP_LOOP_and_320_itm <= (operator_64_false_acc_cse_6_sva_mx0w0[3:0]==4'b0110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_321_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_364 ) begin
      COMP_LOOP_COMP_LOOP_and_321_itm <= (operator_64_false_acc_cse_6_sva_mx0w0[3:0]==4'b0111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_217_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_364 ) begin
      COMP_LOOP_nor_217_itm <= ~((operator_64_false_acc_cse_6_sva_mx0w0[2:0]!=3'b000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_323_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_364 ) begin
      COMP_LOOP_COMP_LOOP_and_323_itm <= (operator_64_false_acc_cse_6_sva_mx0w0[3:0]==4'b1001);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_324_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_364 ) begin
      COMP_LOOP_COMP_LOOP_and_324_itm <= (operator_64_false_acc_cse_6_sva_mx0w0[3:0]==4'b1010);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_325_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_364 ) begin
      COMP_LOOP_COMP_LOOP_and_325_itm <= (operator_64_false_acc_cse_6_sva_mx0w0[3:0]==4'b1011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_326_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_364 ) begin
      COMP_LOOP_COMP_LOOP_and_326_itm <= (operator_64_false_acc_cse_6_sva_mx0w0[3:0]==4'b1100);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_327_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_364 ) begin
      COMP_LOOP_COMP_LOOP_and_327_itm <= (operator_64_false_acc_cse_6_sva_mx0w0[3:0]==4'b1101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_328_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_364 ) begin
      COMP_LOOP_COMP_LOOP_and_328_itm <= (operator_64_false_acc_cse_6_sva_mx0w0[3:0]==4'b1110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_329_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_364 ) begin
      COMP_LOOP_COMP_LOOP_and_329_itm <= (operator_64_false_acc_cse_6_sva_mx0w0[3:0]==4'b1111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_9_psp_sva <= 9'b000000000;
    end
    else if ( mux_2640_nl | (fsm_output[9]) ) begin
      COMP_LOOP_acc_9_psp_sva <= nl_COMP_LOOP_acc_9_psp_sva[8:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      operator_64_false_acc_cse_7_sva <= 10'b0000000000;
    end
    else if ( mux_2641_nl | (fsm_output[9]) ) begin
      operator_64_false_acc_cse_7_sva <= operator_64_false_acc_cse_7_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_nor_25_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_367 ) begin
      COMP_LOOP_COMP_LOOP_nor_25_itm <= ~((operator_64_false_acc_cse_7_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_251_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_367 ) begin
      COMP_LOOP_nor_251_itm <= ~((operator_64_false_acc_cse_7_sva_mx0w0[3:1]!=3'b000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_252_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_367 ) begin
      COMP_LOOP_nor_252_itm <= ~((operator_64_false_acc_cse_7_sva_mx0w0[3]) | (operator_64_false_acc_cse_7_sva_mx0w0[2])
          | (operator_64_false_acc_cse_7_sva_mx0w0[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_377_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_367 ) begin
      COMP_LOOP_COMP_LOOP_and_377_itm <= (operator_64_false_acc_cse_7_sva_mx0w0[3:0]==4'b0011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_254_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_367 ) begin
      COMP_LOOP_nor_254_itm <= ~((operator_64_false_acc_cse_7_sva_mx0w0[3]) | (operator_64_false_acc_cse_7_sva_mx0w0[1])
          | (operator_64_false_acc_cse_7_sva_mx0w0[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_379_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_367 ) begin
      COMP_LOOP_COMP_LOOP_and_379_itm <= (operator_64_false_acc_cse_7_sva_mx0w0[3:0]==4'b0101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_380_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_367 ) begin
      COMP_LOOP_COMP_LOOP_and_380_itm <= (operator_64_false_acc_cse_7_sva_mx0w0[3:0]==4'b0110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_381_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_367 ) begin
      COMP_LOOP_COMP_LOOP_and_381_itm <= (operator_64_false_acc_cse_7_sva_mx0w0[3:0]==4'b0111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_257_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_367 ) begin
      COMP_LOOP_nor_257_itm <= ~((operator_64_false_acc_cse_7_sva_mx0w0[2:0]!=3'b000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_383_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_367 ) begin
      COMP_LOOP_COMP_LOOP_and_383_itm <= (operator_64_false_acc_cse_7_sva_mx0w0[3:0]==4'b1001);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_384_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_367 ) begin
      COMP_LOOP_COMP_LOOP_and_384_itm <= (operator_64_false_acc_cse_7_sva_mx0w0[3:0]==4'b1010);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_385_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_367 ) begin
      COMP_LOOP_COMP_LOOP_and_385_itm <= (operator_64_false_acc_cse_7_sva_mx0w0[3:0]==4'b1011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_386_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_367 ) begin
      COMP_LOOP_COMP_LOOP_and_386_itm <= (operator_64_false_acc_cse_7_sva_mx0w0[3:0]==4'b1100);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_387_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_367 ) begin
      COMP_LOOP_COMP_LOOP_and_387_itm <= (operator_64_false_acc_cse_7_sva_mx0w0[3:0]==4'b1101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_388_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_367 ) begin
      COMP_LOOP_COMP_LOOP_and_388_itm <= (operator_64_false_acc_cse_7_sva_mx0w0[3:0]==4'b1110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_389_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_367 ) begin
      COMP_LOOP_COMP_LOOP_and_389_itm <= (operator_64_false_acc_cse_7_sva_mx0w0[3:0]==4'b1111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_cse_8_sva <= 10'b0000000000;
    end
    else if ( mux_2645_nl | (fsm_output[9]) ) begin
      COMP_LOOP_acc_cse_8_sva <= nl_COMP_LOOP_acc_cse_8_sva[9:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      operator_64_false_acc_cse_8_sva <= 10'b0000000000;
    end
    else if ( mux_2649_nl | (fsm_output[9]) ) begin
      operator_64_false_acc_cse_8_sva <= operator_64_false_acc_cse_8_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_nor_29_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_370 ) begin
      COMP_LOOP_COMP_LOOP_nor_29_itm <= ~((operator_64_false_acc_cse_8_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_291_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_370 ) begin
      COMP_LOOP_nor_291_itm <= ~((operator_64_false_acc_cse_8_sva_mx0w0[3:1]!=3'b000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_292_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_370 ) begin
      COMP_LOOP_nor_292_itm <= ~((operator_64_false_acc_cse_8_sva_mx0w0[3]) | (operator_64_false_acc_cse_8_sva_mx0w0[2])
          | (operator_64_false_acc_cse_8_sva_mx0w0[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_437_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_370 ) begin
      COMP_LOOP_COMP_LOOP_and_437_itm <= (operator_64_false_acc_cse_8_sva_mx0w0[3:0]==4'b0011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_294_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_370 ) begin
      COMP_LOOP_nor_294_itm <= ~((operator_64_false_acc_cse_8_sva_mx0w0[3]) | (operator_64_false_acc_cse_8_sva_mx0w0[1])
          | (operator_64_false_acc_cse_8_sva_mx0w0[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_439_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_370 ) begin
      COMP_LOOP_COMP_LOOP_and_439_itm <= (operator_64_false_acc_cse_8_sva_mx0w0[3:0]==4'b0101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_440_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_370 ) begin
      COMP_LOOP_COMP_LOOP_and_440_itm <= (operator_64_false_acc_cse_8_sva_mx0w0[3:0]==4'b0110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_441_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_370 ) begin
      COMP_LOOP_COMP_LOOP_and_441_itm <= (operator_64_false_acc_cse_8_sva_mx0w0[3:0]==4'b0111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_297_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_370 ) begin
      COMP_LOOP_nor_297_itm <= ~((operator_64_false_acc_cse_8_sva_mx0w0[2:0]!=3'b000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_443_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_370 ) begin
      COMP_LOOP_COMP_LOOP_and_443_itm <= (operator_64_false_acc_cse_8_sva_mx0w0[3:0]==4'b1001);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_444_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_370 ) begin
      COMP_LOOP_COMP_LOOP_and_444_itm <= (operator_64_false_acc_cse_8_sva_mx0w0[3:0]==4'b1010);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_445_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_370 ) begin
      COMP_LOOP_COMP_LOOP_and_445_itm <= (operator_64_false_acc_cse_8_sva_mx0w0[3:0]==4'b1011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_446_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_370 ) begin
      COMP_LOOP_COMP_LOOP_and_446_itm <= (operator_64_false_acc_cse_8_sva_mx0w0[3:0]==4'b1100);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_447_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_370 ) begin
      COMP_LOOP_COMP_LOOP_and_447_itm <= (operator_64_false_acc_cse_8_sva_mx0w0[3:0]==4'b1101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_448_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_370 ) begin
      COMP_LOOP_COMP_LOOP_and_448_itm <= (operator_64_false_acc_cse_8_sva_mx0w0[3:0]==4'b1110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_449_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_370 ) begin
      COMP_LOOP_COMP_LOOP_and_449_itm <= (operator_64_false_acc_cse_8_sva_mx0w0[3:0]==4'b1111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_10_psp_sva <= 7'b0000000;
    end
    else if ( mux_2657_nl | (fsm_output[9]) ) begin
      COMP_LOOP_acc_10_psp_sva <= nl_COMP_LOOP_acc_10_psp_sva[6:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      operator_64_false_acc_cse_9_sva <= 10'b0000000000;
    end
    else if ( MUX_s_1_2_2(not_tmp_698, or_2651_nl, fsm_output[9]) ) begin
      operator_64_false_acc_cse_9_sva <= operator_64_false_acc_cse_9_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_nor_33_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_372 ) begin
      COMP_LOOP_COMP_LOOP_nor_33_itm <= ~((operator_64_false_acc_cse_9_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_331_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_372 ) begin
      COMP_LOOP_nor_331_itm <= ~((operator_64_false_acc_cse_9_sva_mx0w0[3:1]!=3'b000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_332_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_372 ) begin
      COMP_LOOP_nor_332_itm <= ~((operator_64_false_acc_cse_9_sva_mx0w0[3]) | (operator_64_false_acc_cse_9_sva_mx0w0[2])
          | (operator_64_false_acc_cse_9_sva_mx0w0[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_497_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_372 ) begin
      COMP_LOOP_COMP_LOOP_and_497_itm <= (operator_64_false_acc_cse_9_sva_mx0w0[3:0]==4'b0011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_334_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_372 ) begin
      COMP_LOOP_nor_334_itm <= ~((operator_64_false_acc_cse_9_sva_mx0w0[3]) | (operator_64_false_acc_cse_9_sva_mx0w0[1])
          | (operator_64_false_acc_cse_9_sva_mx0w0[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_499_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_372 ) begin
      COMP_LOOP_COMP_LOOP_and_499_itm <= (operator_64_false_acc_cse_9_sva_mx0w0[3:0]==4'b0101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_500_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_372 ) begin
      COMP_LOOP_COMP_LOOP_and_500_itm <= (operator_64_false_acc_cse_9_sva_mx0w0[3:0]==4'b0110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_501_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_372 ) begin
      COMP_LOOP_COMP_LOOP_and_501_itm <= (operator_64_false_acc_cse_9_sva_mx0w0[3:0]==4'b0111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_337_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_372 ) begin
      COMP_LOOP_nor_337_itm <= ~((operator_64_false_acc_cse_9_sva_mx0w0[2:0]!=3'b000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_503_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_372 ) begin
      COMP_LOOP_COMP_LOOP_and_503_itm <= (operator_64_false_acc_cse_9_sva_mx0w0[3:0]==4'b1001);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_504_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_372 ) begin
      COMP_LOOP_COMP_LOOP_and_504_itm <= (operator_64_false_acc_cse_9_sva_mx0w0[3:0]==4'b1010);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_505_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_372 ) begin
      COMP_LOOP_COMP_LOOP_and_505_itm <= (operator_64_false_acc_cse_9_sva_mx0w0[3:0]==4'b1011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_506_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_372 ) begin
      COMP_LOOP_COMP_LOOP_and_506_itm <= (operator_64_false_acc_cse_9_sva_mx0w0[3:0]==4'b1100);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_507_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_372 ) begin
      COMP_LOOP_COMP_LOOP_and_507_itm <= (operator_64_false_acc_cse_9_sva_mx0w0[3:0]==4'b1101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_508_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_372 ) begin
      COMP_LOOP_COMP_LOOP_and_508_itm <= (operator_64_false_acc_cse_9_sva_mx0w0[3:0]==4'b1110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_509_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_372 ) begin
      COMP_LOOP_COMP_LOOP_and_509_itm <= (operator_64_false_acc_cse_9_sva_mx0w0[3:0]==4'b1111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_cse_10_sva <= 10'b0000000000;
    end
    else if ( MUX_s_1_2_2(not_tmp_698, or_2732_nl, fsm_output[9]) ) begin
      COMP_LOOP_acc_cse_10_sva <= nl_COMP_LOOP_acc_cse_10_sva[9:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      operator_64_false_acc_cse_10_sva <= 10'b0000000000;
    end
    else if ( MUX_s_1_2_2(mux_2670_nl, (fsm_output[9]), or_2733_cse) ) begin
      operator_64_false_acc_cse_10_sva <= operator_64_false_acc_cse_10_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_nor_37_itm <= 1'b0;
    end
    else if ( ~ not_tmp_706 ) begin
      COMP_LOOP_COMP_LOOP_nor_37_itm <= ~((operator_64_false_acc_cse_10_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_371_itm <= 1'b0;
    end
    else if ( ~ not_tmp_706 ) begin
      COMP_LOOP_nor_371_itm <= ~((operator_64_false_acc_cse_10_sva_mx0w0[3:1]!=3'b000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_372_itm <= 1'b0;
    end
    else if ( ~ not_tmp_706 ) begin
      COMP_LOOP_nor_372_itm <= ~((operator_64_false_acc_cse_10_sva_mx0w0[3]) | (operator_64_false_acc_cse_10_sva_mx0w0[2])
          | (operator_64_false_acc_cse_10_sva_mx0w0[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_557_itm <= 1'b0;
    end
    else if ( ~ not_tmp_706 ) begin
      COMP_LOOP_COMP_LOOP_and_557_itm <= (operator_64_false_acc_cse_10_sva_mx0w0[3:0]==4'b0011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_374_itm <= 1'b0;
    end
    else if ( ~ not_tmp_706 ) begin
      COMP_LOOP_nor_374_itm <= ~((operator_64_false_acc_cse_10_sva_mx0w0[3]) | (operator_64_false_acc_cse_10_sva_mx0w0[1])
          | (operator_64_false_acc_cse_10_sva_mx0w0[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_559_itm <= 1'b0;
    end
    else if ( ~ not_tmp_706 ) begin
      COMP_LOOP_COMP_LOOP_and_559_itm <= (operator_64_false_acc_cse_10_sva_mx0w0[3:0]==4'b0101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_560_itm <= 1'b0;
    end
    else if ( ~ not_tmp_706 ) begin
      COMP_LOOP_COMP_LOOP_and_560_itm <= (operator_64_false_acc_cse_10_sva_mx0w0[3:0]==4'b0110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_561_itm <= 1'b0;
    end
    else if ( ~ not_tmp_706 ) begin
      COMP_LOOP_COMP_LOOP_and_561_itm <= (operator_64_false_acc_cse_10_sva_mx0w0[3:0]==4'b0111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_377_itm <= 1'b0;
    end
    else if ( ~ not_tmp_706 ) begin
      COMP_LOOP_nor_377_itm <= ~((operator_64_false_acc_cse_10_sva_mx0w0[2:0]!=3'b000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_563_itm <= 1'b0;
    end
    else if ( ~ not_tmp_706 ) begin
      COMP_LOOP_COMP_LOOP_and_563_itm <= (operator_64_false_acc_cse_10_sva_mx0w0[3:0]==4'b1001);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_564_itm <= 1'b0;
    end
    else if ( ~ not_tmp_706 ) begin
      COMP_LOOP_COMP_LOOP_and_564_itm <= (operator_64_false_acc_cse_10_sva_mx0w0[3:0]==4'b1010);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_565_itm <= 1'b0;
    end
    else if ( ~ not_tmp_706 ) begin
      COMP_LOOP_COMP_LOOP_and_565_itm <= (operator_64_false_acc_cse_10_sva_mx0w0[3:0]==4'b1011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_566_itm <= 1'b0;
    end
    else if ( ~ not_tmp_706 ) begin
      COMP_LOOP_COMP_LOOP_and_566_itm <= (operator_64_false_acc_cse_10_sva_mx0w0[3:0]==4'b1100);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_567_itm <= 1'b0;
    end
    else if ( ~ not_tmp_706 ) begin
      COMP_LOOP_COMP_LOOP_and_567_itm <= (operator_64_false_acc_cse_10_sva_mx0w0[3:0]==4'b1101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_568_itm <= 1'b0;
    end
    else if ( ~ not_tmp_706 ) begin
      COMP_LOOP_COMP_LOOP_and_568_itm <= (operator_64_false_acc_cse_10_sva_mx0w0[3:0]==4'b1110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_569_itm <= 1'b0;
    end
    else if ( ~ not_tmp_706 ) begin
      COMP_LOOP_COMP_LOOP_and_569_itm <= (operator_64_false_acc_cse_10_sva_mx0w0[3:0]==4'b1111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_11_psp_sva <= 9'b000000000;
    end
    else if ( MUX_s_1_2_2(mux_2681_nl, and_tmp_32, fsm_output[5]) ) begin
      COMP_LOOP_acc_11_psp_sva <= nl_COMP_LOOP_acc_11_psp_sva[8:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      operator_64_false_acc_cse_11_sva <= 10'b0000000000;
    end
    else if ( MUX_s_1_2_2(not_tmp_698, or_2743_nl, fsm_output[9]) ) begin
      operator_64_false_acc_cse_11_sva <= operator_64_false_acc_cse_11_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_nor_41_itm <= 1'b0;
      COMP_LOOP_nor_411_itm <= 1'b0;
      COMP_LOOP_nor_412_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_617_itm <= 1'b0;
      COMP_LOOP_nor_414_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_619_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_620_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_621_itm <= 1'b0;
      COMP_LOOP_nor_417_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_623_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_624_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_625_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_626_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_627_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_628_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_629_itm <= 1'b0;
    end
    else if ( mux_2688_itm ) begin
      COMP_LOOP_COMP_LOOP_nor_41_itm <= ~((operator_64_false_acc_cse_11_sva_mx0w0[3:0]!=4'b0000));
      COMP_LOOP_nor_411_itm <= ~((operator_64_false_acc_cse_11_sva_mx0w0[3:1]!=3'b000));
      COMP_LOOP_nor_412_itm <= ~((operator_64_false_acc_cse_11_sva_mx0w0[3]) | (operator_64_false_acc_cse_11_sva_mx0w0[2])
          | (operator_64_false_acc_cse_11_sva_mx0w0[0]));
      COMP_LOOP_COMP_LOOP_and_617_itm <= (operator_64_false_acc_cse_11_sva_mx0w0[3:0]==4'b0011);
      COMP_LOOP_nor_414_itm <= ~((operator_64_false_acc_cse_11_sva_mx0w0[3]) | (operator_64_false_acc_cse_11_sva_mx0w0[1])
          | (operator_64_false_acc_cse_11_sva_mx0w0[0]));
      COMP_LOOP_COMP_LOOP_and_619_itm <= (operator_64_false_acc_cse_11_sva_mx0w0[3:0]==4'b0101);
      COMP_LOOP_COMP_LOOP_and_620_itm <= (operator_64_false_acc_cse_11_sva_mx0w0[3:0]==4'b0110);
      COMP_LOOP_COMP_LOOP_and_621_itm <= (operator_64_false_acc_cse_11_sva_mx0w0[3:0]==4'b0111);
      COMP_LOOP_nor_417_itm <= ~((operator_64_false_acc_cse_11_sva_mx0w0[2:0]!=3'b000));
      COMP_LOOP_COMP_LOOP_and_623_itm <= (operator_64_false_acc_cse_11_sva_mx0w0[3:0]==4'b1001);
      COMP_LOOP_COMP_LOOP_and_624_itm <= (operator_64_false_acc_cse_11_sva_mx0w0[3:0]==4'b1010);
      COMP_LOOP_COMP_LOOP_and_625_itm <= (operator_64_false_acc_cse_11_sva_mx0w0[3:0]==4'b1011);
      COMP_LOOP_COMP_LOOP_and_626_itm <= (operator_64_false_acc_cse_11_sva_mx0w0[3:0]==4'b1100);
      COMP_LOOP_COMP_LOOP_and_627_itm <= (operator_64_false_acc_cse_11_sva_mx0w0[3:0]==4'b1101);
      COMP_LOOP_COMP_LOOP_and_628_itm <= (operator_64_false_acc_cse_11_sva_mx0w0[3:0]==4'b1110);
      COMP_LOOP_COMP_LOOP_and_629_itm <= (operator_64_false_acc_cse_11_sva_mx0w0[3:0]==4'b1111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_cse_12_sva <= 10'b0000000000;
    end
    else if ( MUX_s_1_2_2(not_tmp_698, or_2748_nl, fsm_output[9]) ) begin
      COMP_LOOP_acc_cse_12_sva <= nl_COMP_LOOP_acc_cse_12_sva[9:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      operator_64_false_acc_cse_12_sva <= 10'b0000000000;
    end
    else if ( MUX_s_1_2_2(mux_2692_nl, (fsm_output[9]), fsm_output[8]) ) begin
      operator_64_false_acc_cse_12_sva <= operator_64_false_acc_cse_12_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_nor_45_itm <= 1'b0;
      COMP_LOOP_nor_451_itm <= 1'b0;
      COMP_LOOP_nor_452_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_677_itm <= 1'b0;
      COMP_LOOP_nor_454_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_679_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_680_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_681_itm <= 1'b0;
      COMP_LOOP_nor_457_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_683_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_684_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_685_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_686_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_687_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_688_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_689_itm <= 1'b0;
    end
    else if ( mux_2703_itm ) begin
      COMP_LOOP_COMP_LOOP_nor_45_itm <= ~((operator_64_false_acc_cse_12_sva_mx0w0[3:0]!=4'b0000));
      COMP_LOOP_nor_451_itm <= ~((operator_64_false_acc_cse_12_sva_mx0w0[3:1]!=3'b000));
      COMP_LOOP_nor_452_itm <= ~((operator_64_false_acc_cse_12_sva_mx0w0[3]) | (operator_64_false_acc_cse_12_sva_mx0w0[2])
          | (operator_64_false_acc_cse_12_sva_mx0w0[0]));
      COMP_LOOP_COMP_LOOP_and_677_itm <= (operator_64_false_acc_cse_12_sva_mx0w0[3:0]==4'b0011);
      COMP_LOOP_nor_454_itm <= ~((operator_64_false_acc_cse_12_sva_mx0w0[3]) | (operator_64_false_acc_cse_12_sva_mx0w0[1])
          | (operator_64_false_acc_cse_12_sva_mx0w0[0]));
      COMP_LOOP_COMP_LOOP_and_679_itm <= (operator_64_false_acc_cse_12_sva_mx0w0[3:0]==4'b0101);
      COMP_LOOP_COMP_LOOP_and_680_itm <= (operator_64_false_acc_cse_12_sva_mx0w0[3:0]==4'b0110);
      COMP_LOOP_COMP_LOOP_and_681_itm <= (operator_64_false_acc_cse_12_sva_mx0w0[3:0]==4'b0111);
      COMP_LOOP_nor_457_itm <= ~((operator_64_false_acc_cse_12_sva_mx0w0[2:0]!=3'b000));
      COMP_LOOP_COMP_LOOP_and_683_itm <= (operator_64_false_acc_cse_12_sva_mx0w0[3:0]==4'b1001);
      COMP_LOOP_COMP_LOOP_and_684_itm <= (operator_64_false_acc_cse_12_sva_mx0w0[3:0]==4'b1010);
      COMP_LOOP_COMP_LOOP_and_685_itm <= (operator_64_false_acc_cse_12_sva_mx0w0[3:0]==4'b1011);
      COMP_LOOP_COMP_LOOP_and_686_itm <= (operator_64_false_acc_cse_12_sva_mx0w0[3:0]==4'b1100);
      COMP_LOOP_COMP_LOOP_and_687_itm <= (operator_64_false_acc_cse_12_sva_mx0w0[3:0]==4'b1101);
      COMP_LOOP_COMP_LOOP_and_688_itm <= (operator_64_false_acc_cse_12_sva_mx0w0[3:0]==4'b1110);
      COMP_LOOP_COMP_LOOP_and_689_itm <= (operator_64_false_acc_cse_12_sva_mx0w0[3:0]==4'b1111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_12_psp_sva <= 8'b00000000;
    end
    else if ( MUX_s_1_2_2(mux_2708_nl, (fsm_output[9]), fsm_output[8]) ) begin
      COMP_LOOP_acc_12_psp_sva <= z_out_2[7:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      operator_64_false_acc_cse_13_sva <= 10'b0000000000;
    end
    else if ( MUX_s_1_2_2(mux_2713_nl, (fsm_output[9]), fsm_output[8]) ) begin
      operator_64_false_acc_cse_13_sva <= operator_64_false_acc_cse_13_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_nor_49_itm <= 1'b0;
      COMP_LOOP_nor_491_itm <= 1'b0;
      COMP_LOOP_nor_492_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_737_itm <= 1'b0;
      COMP_LOOP_nor_494_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_739_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_740_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_741_itm <= 1'b0;
      COMP_LOOP_nor_497_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_743_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_744_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_745_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_746_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_747_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_748_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_749_itm <= 1'b0;
    end
    else if ( mux_2715_itm ) begin
      COMP_LOOP_COMP_LOOP_nor_49_itm <= ~((operator_64_false_acc_cse_13_sva_mx0w0[3:0]!=4'b0000));
      COMP_LOOP_nor_491_itm <= ~((operator_64_false_acc_cse_13_sva_mx0w0[3:1]!=3'b000));
      COMP_LOOP_nor_492_itm <= ~((operator_64_false_acc_cse_13_sva_mx0w0[3]) | (operator_64_false_acc_cse_13_sva_mx0w0[2])
          | (operator_64_false_acc_cse_13_sva_mx0w0[0]));
      COMP_LOOP_COMP_LOOP_and_737_itm <= (operator_64_false_acc_cse_13_sva_mx0w0[3:0]==4'b0011);
      COMP_LOOP_nor_494_itm <= ~((operator_64_false_acc_cse_13_sva_mx0w0[3]) | (operator_64_false_acc_cse_13_sva_mx0w0[1])
          | (operator_64_false_acc_cse_13_sva_mx0w0[0]));
      COMP_LOOP_COMP_LOOP_and_739_itm <= (operator_64_false_acc_cse_13_sva_mx0w0[3:0]==4'b0101);
      COMP_LOOP_COMP_LOOP_and_740_itm <= (operator_64_false_acc_cse_13_sva_mx0w0[3:0]==4'b0110);
      COMP_LOOP_COMP_LOOP_and_741_itm <= (operator_64_false_acc_cse_13_sva_mx0w0[3:0]==4'b0111);
      COMP_LOOP_nor_497_itm <= ~((operator_64_false_acc_cse_13_sva_mx0w0[2:0]!=3'b000));
      COMP_LOOP_COMP_LOOP_and_743_itm <= (operator_64_false_acc_cse_13_sva_mx0w0[3:0]==4'b1001);
      COMP_LOOP_COMP_LOOP_and_744_itm <= (operator_64_false_acc_cse_13_sva_mx0w0[3:0]==4'b1010);
      COMP_LOOP_COMP_LOOP_and_745_itm <= (operator_64_false_acc_cse_13_sva_mx0w0[3:0]==4'b1011);
      COMP_LOOP_COMP_LOOP_and_746_itm <= (operator_64_false_acc_cse_13_sva_mx0w0[3:0]==4'b1100);
      COMP_LOOP_COMP_LOOP_and_747_itm <= (operator_64_false_acc_cse_13_sva_mx0w0[3:0]==4'b1101);
      COMP_LOOP_COMP_LOOP_and_748_itm <= (operator_64_false_acc_cse_13_sva_mx0w0[3:0]==4'b1110);
      COMP_LOOP_COMP_LOOP_and_749_itm <= (operator_64_false_acc_cse_13_sva_mx0w0[3:0]==4'b1111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_cse_14_sva <= 10'b0000000000;
    end
    else if ( MUX_s_1_2_2(not_tmp_698, and_410_nl, fsm_output[9]) ) begin
      COMP_LOOP_acc_cse_14_sva <= nl_COMP_LOOP_acc_cse_14_sva[9:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      operator_64_false_acc_cse_14_sva <= 10'b0000000000;
    end
    else if ( MUX_s_1_2_2(mux_2722_nl, nor_tmp_130, or_111_cse) ) begin
      operator_64_false_acc_cse_14_sva <= operator_64_false_acc_cse_14_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_nor_53_itm <= 1'b0;
      COMP_LOOP_nor_531_itm <= 1'b0;
      COMP_LOOP_nor_532_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_797_itm <= 1'b0;
      COMP_LOOP_nor_534_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_799_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_800_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_801_itm <= 1'b0;
      COMP_LOOP_nor_537_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_803_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_804_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_805_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_806_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_807_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_808_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_809_itm <= 1'b0;
    end
    else if ( mux_2727_itm ) begin
      COMP_LOOP_COMP_LOOP_nor_53_itm <= ~((operator_64_false_acc_cse_14_sva_mx0w0[3:0]!=4'b0000));
      COMP_LOOP_nor_531_itm <= ~((operator_64_false_acc_cse_14_sva_mx0w0[3:1]!=3'b000));
      COMP_LOOP_nor_532_itm <= ~((operator_64_false_acc_cse_14_sva_mx0w0[3]) | (operator_64_false_acc_cse_14_sva_mx0w0[2])
          | (operator_64_false_acc_cse_14_sva_mx0w0[0]));
      COMP_LOOP_COMP_LOOP_and_797_itm <= (operator_64_false_acc_cse_14_sva_mx0w0[3:0]==4'b0011);
      COMP_LOOP_nor_534_itm <= ~((operator_64_false_acc_cse_14_sva_mx0w0[3]) | (operator_64_false_acc_cse_14_sva_mx0w0[1])
          | (operator_64_false_acc_cse_14_sva_mx0w0[0]));
      COMP_LOOP_COMP_LOOP_and_799_itm <= (operator_64_false_acc_cse_14_sva_mx0w0[3:0]==4'b0101);
      COMP_LOOP_COMP_LOOP_and_800_itm <= (operator_64_false_acc_cse_14_sva_mx0w0[3:0]==4'b0110);
      COMP_LOOP_COMP_LOOP_and_801_itm <= (operator_64_false_acc_cse_14_sva_mx0w0[3:0]==4'b0111);
      COMP_LOOP_nor_537_itm <= ~((operator_64_false_acc_cse_14_sva_mx0w0[2:0]!=3'b000));
      COMP_LOOP_COMP_LOOP_and_803_itm <= (operator_64_false_acc_cse_14_sva_mx0w0[3:0]==4'b1001);
      COMP_LOOP_COMP_LOOP_and_804_itm <= (operator_64_false_acc_cse_14_sva_mx0w0[3:0]==4'b1010);
      COMP_LOOP_COMP_LOOP_and_805_itm <= (operator_64_false_acc_cse_14_sva_mx0w0[3:0]==4'b1011);
      COMP_LOOP_COMP_LOOP_and_806_itm <= (operator_64_false_acc_cse_14_sva_mx0w0[3:0]==4'b1100);
      COMP_LOOP_COMP_LOOP_and_807_itm <= (operator_64_false_acc_cse_14_sva_mx0w0[3:0]==4'b1101);
      COMP_LOOP_COMP_LOOP_and_808_itm <= (operator_64_false_acc_cse_14_sva_mx0w0[3:0]==4'b1110);
      COMP_LOOP_COMP_LOOP_and_809_itm <= (operator_64_false_acc_cse_14_sva_mx0w0[3:0]==4'b1111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_13_psp_sva <= 9'b000000000;
    end
    else if ( ~ mux_2730_nl ) begin
      COMP_LOOP_acc_13_psp_sva <= nl_COMP_LOOP_acc_13_psp_sva[8:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      operator_64_false_acc_cse_15_sva <= 10'b0000000000;
    end
    else if ( ~ mux_2733_nl ) begin
      operator_64_false_acc_cse_15_sva <= operator_64_false_acc_cse_15_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_nor_57_itm <= 1'b0;
      COMP_LOOP_nor_571_itm <= 1'b0;
      COMP_LOOP_nor_572_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_857_itm <= 1'b0;
      COMP_LOOP_nor_574_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_859_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_860_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_861_itm <= 1'b0;
      COMP_LOOP_nor_577_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_863_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_864_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_865_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_866_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_867_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_868_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_869_itm <= 1'b0;
    end
    else if ( mux_2734_itm ) begin
      COMP_LOOP_COMP_LOOP_nor_57_itm <= ~((operator_64_false_acc_cse_15_sva_mx0w0[3:0]!=4'b0000));
      COMP_LOOP_nor_571_itm <= ~((operator_64_false_acc_cse_15_sva_mx0w0[3:1]!=3'b000));
      COMP_LOOP_nor_572_itm <= ~((operator_64_false_acc_cse_15_sva_mx0w0[3]) | (operator_64_false_acc_cse_15_sva_mx0w0[2])
          | (operator_64_false_acc_cse_15_sva_mx0w0[0]));
      COMP_LOOP_COMP_LOOP_and_857_itm <= (operator_64_false_acc_cse_15_sva_mx0w0[3:0]==4'b0011);
      COMP_LOOP_nor_574_itm <= ~((operator_64_false_acc_cse_15_sva_mx0w0[3]) | (operator_64_false_acc_cse_15_sva_mx0w0[1])
          | (operator_64_false_acc_cse_15_sva_mx0w0[0]));
      COMP_LOOP_COMP_LOOP_and_859_itm <= (operator_64_false_acc_cse_15_sva_mx0w0[3:0]==4'b0101);
      COMP_LOOP_COMP_LOOP_and_860_itm <= (operator_64_false_acc_cse_15_sva_mx0w0[3:0]==4'b0110);
      COMP_LOOP_COMP_LOOP_and_861_itm <= (operator_64_false_acc_cse_15_sva_mx0w0[3:0]==4'b0111);
      COMP_LOOP_nor_577_itm <= ~((operator_64_false_acc_cse_15_sva_mx0w0[2:0]!=3'b000));
      COMP_LOOP_COMP_LOOP_and_863_itm <= (operator_64_false_acc_cse_15_sva_mx0w0[3:0]==4'b1001);
      COMP_LOOP_COMP_LOOP_and_864_itm <= (operator_64_false_acc_cse_15_sva_mx0w0[3:0]==4'b1010);
      COMP_LOOP_COMP_LOOP_and_865_itm <= (operator_64_false_acc_cse_15_sva_mx0w0[3:0]==4'b1011);
      COMP_LOOP_COMP_LOOP_and_866_itm <= (operator_64_false_acc_cse_15_sva_mx0w0[3:0]==4'b1100);
      COMP_LOOP_COMP_LOOP_and_867_itm <= (operator_64_false_acc_cse_15_sva_mx0w0[3:0]==4'b1101);
      COMP_LOOP_COMP_LOOP_and_868_itm <= (operator_64_false_acc_cse_15_sva_mx0w0[3:0]==4'b1110);
      COMP_LOOP_COMP_LOOP_and_869_itm <= (operator_64_false_acc_cse_15_sva_mx0w0[3:0]==4'b1111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_cse_sva <= 10'b0000000000;
    end
    else if ( MUX_s_1_2_2(not_tmp_698, and_413_nl, fsm_output[9]) ) begin
      COMP_LOOP_acc_cse_sva <= nl_COMP_LOOP_acc_cse_sva[9:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      operator_64_false_acc_cse_sva <= 10'b0000000000;
    end
    else if ( MUX_s_1_2_2(not_tmp_698, and_414_nl, fsm_output[9]) ) begin
      operator_64_false_acc_cse_sva <= operator_64_false_acc_cse_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_nor_61_itm <= 1'b0;
      COMP_LOOP_nor_611_itm <= 1'b0;
      COMP_LOOP_nor_612_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_917_itm <= 1'b0;
      COMP_LOOP_nor_614_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_919_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_920_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_921_itm <= 1'b0;
      COMP_LOOP_nor_617_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_923_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_924_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_925_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_926_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_927_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_928_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_929_itm <= 1'b0;
    end
    else if ( mux_2745_itm ) begin
      COMP_LOOP_COMP_LOOP_nor_61_itm <= ~((operator_64_false_acc_cse_sva_mx0w0[3:0]!=4'b0000));
      COMP_LOOP_nor_611_itm <= ~((operator_64_false_acc_cse_sva_mx0w0[3:1]!=3'b000));
      COMP_LOOP_nor_612_itm <= ~((operator_64_false_acc_cse_sva_mx0w0[3]) | (operator_64_false_acc_cse_sva_mx0w0[2])
          | (operator_64_false_acc_cse_sva_mx0w0[0]));
      COMP_LOOP_COMP_LOOP_and_917_itm <= (operator_64_false_acc_cse_sva_mx0w0[3:0]==4'b0011);
      COMP_LOOP_nor_614_itm <= ~((operator_64_false_acc_cse_sva_mx0w0[3]) | (operator_64_false_acc_cse_sva_mx0w0[1])
          | (operator_64_false_acc_cse_sva_mx0w0[0]));
      COMP_LOOP_COMP_LOOP_and_919_itm <= (operator_64_false_acc_cse_sva_mx0w0[3:0]==4'b0101);
      COMP_LOOP_COMP_LOOP_and_920_itm <= (operator_64_false_acc_cse_sva_mx0w0[3:0]==4'b0110);
      COMP_LOOP_COMP_LOOP_and_921_itm <= (operator_64_false_acc_cse_sva_mx0w0[3:0]==4'b0111);
      COMP_LOOP_nor_617_itm <= ~((operator_64_false_acc_cse_sva_mx0w0[2:0]!=3'b000));
      COMP_LOOP_COMP_LOOP_and_923_itm <= (operator_64_false_acc_cse_sva_mx0w0[3:0]==4'b1001);
      COMP_LOOP_COMP_LOOP_and_924_itm <= (operator_64_false_acc_cse_sva_mx0w0[3:0]==4'b1010);
      COMP_LOOP_COMP_LOOP_and_925_itm <= (operator_64_false_acc_cse_sva_mx0w0[3:0]==4'b1011);
      COMP_LOOP_COMP_LOOP_and_926_itm <= (operator_64_false_acc_cse_sva_mx0w0[3:0]==4'b1100);
      COMP_LOOP_COMP_LOOP_and_927_itm <= (operator_64_false_acc_cse_sva_mx0w0[3:0]==4'b1101);
      COMP_LOOP_COMP_LOOP_and_928_itm <= (operator_64_false_acc_cse_sva_mx0w0[3:0]==4'b1110);
      COMP_LOOP_COMP_LOOP_and_929_itm <= (operator_64_false_acc_cse_sva_mx0w0[3:0]==4'b1111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      operator_64_false_slc_operator_64_false_acc_1_60_itm <= 1'b0;
    end
    else if ( and_dcpl_98 | operator_64_false_slc_operator_64_false_acc_1_60_itm_mx0c1
        | operator_64_false_slc_operator_64_false_acc_1_60_itm_mx0c2 | operator_64_false_slc_operator_64_false_acc_1_60_itm_mx0c3
        | operator_64_false_slc_operator_64_false_acc_1_60_itm_mx0c4 ) begin
      operator_64_false_slc_operator_64_false_acc_1_60_itm <= MUX1HOT_s_1_4_2(COMP_LOOP_nor_11_nl,
          (z_out_2[61]), (COMP_LOOP_slc_acc_3_12_1_slc[11]), (z_out_2[59]), {and_dcpl_98
          , COMP_LOOP_or_35_nl , operator_64_false_slc_operator_64_false_acc_1_60_itm_mx0c2
          , operator_64_false_slc_operator_64_false_acc_1_60_itm_mx0c4});
    end
  end
  always @(posedge clk) begin
    if ( tmp_1_lpi_4_dfm_mx0c0 | and_dcpl_245 | and_dcpl_249 | and_dcpl_254 | and_dcpl_258
        | and_dcpl_262 | and_dcpl_265 | and_dcpl_269 | and_dcpl_271 | and_dcpl_273
        | and_dcpl_276 | and_dcpl_278 | and_dcpl_283 | and_dcpl_285 | and_dcpl_287
        | and_dcpl_289 ) begin
      tmp_1_lpi_4_dfm <= MUX1HOT_v_64_16_2(vec_rsc_0_0_i_qa_d, vec_rsc_0_1_i_qa_d,
          vec_rsc_0_2_i_qa_d, vec_rsc_0_3_i_qa_d, vec_rsc_0_4_i_qa_d, vec_rsc_0_5_i_qa_d,
          vec_rsc_0_6_i_qa_d, vec_rsc_0_7_i_qa_d, vec_rsc_0_8_i_qa_d, vec_rsc_0_9_i_qa_d,
          vec_rsc_0_10_i_qa_d, vec_rsc_0_11_i_qa_d, vec_rsc_0_12_i_qa_d, vec_rsc_0_13_i_qa_d,
          vec_rsc_0_14_i_qa_d, vec_rsc_0_15_i_qa_d, {COMP_LOOP_or_18_nl , COMP_LOOP_or_19_nl
          , COMP_LOOP_or_20_nl , COMP_LOOP_or_21_nl , COMP_LOOP_or_22_nl , COMP_LOOP_or_23_nl
          , COMP_LOOP_or_24_nl , COMP_LOOP_or_25_nl , COMP_LOOP_or_26_nl , COMP_LOOP_or_27_nl
          , COMP_LOOP_or_28_nl , COMP_LOOP_or_29_nl , COMP_LOOP_or_30_nl , COMP_LOOP_or_31_nl
          , COMP_LOOP_or_32_nl , COMP_LOOP_or_33_nl});
    end
  end
  always @(posedge clk) begin
    if ( mux_2797_itm ) begin
      modExp_dev_exp_1_sva_8_4 <= MUX_v_5_2_2((z_out_3[8:4]), COMP_LOOP_k_9_4_sva_4_0,
          mux_2336_itm);
    end
  end
  always @(posedge clk) begin
    if ( MUX_s_1_2_2(mux_2893_nl, mux_2884_nl, fsm_output[8]) ) begin
      modExp_dev_exp_1_sva_63_9 <= MUX_v_55_2_2(55'b0000000000000000000000000000000000000000000000000000000,
          (z_out_3[63:9]), not_7089_nl);
    end
  end
  assign or_2479_nl = (fsm_output[2]) | not_tmp_572;
  assign mux_2317_nl = MUX_s_1_2_2(not_tmp_572, or_2733_cse, fsm_output[2]);
  assign mux_2318_nl = MUX_s_1_2_2(or_2479_nl, mux_2317_nl, fsm_output[1]);
  assign mux_2319_nl = MUX_s_1_2_2(mux_2318_nl, or_tmp_2391, fsm_output[5]);
  assign mux_2320_nl = MUX_s_1_2_2(mux_2319_nl, mux_tmp_2244, fsm_output[6]);
  assign mux_2314_nl = MUX_s_1_2_2(or_tmp_2402, or_tmp_2401, fsm_output[1]);
  assign nand_177_nl = ~((and_515_cse | (fsm_output[2])) & (fsm_output[8:7]==2'b11));
  assign mux_2315_nl = MUX_s_1_2_2(mux_2314_nl, nand_177_nl, fsm_output[5]);
  assign or_2477_nl = and_516_cse | not_tmp_572;
  assign mux_2313_nl = MUX_s_1_2_2(or_tmp_2324, or_2477_nl, fsm_output[5]);
  assign mux_2316_nl = MUX_s_1_2_2(mux_2315_nl, mux_2313_nl, fsm_output[6]);
  assign mux_2321_nl = MUX_s_1_2_2(mux_2320_nl, mux_2316_nl, fsm_output[4]);
  assign or_2476_nl = and_516_cse | (fsm_output[8:7]!=2'b00);
  assign mux_2310_nl = MUX_s_1_2_2((fsm_output[7]), or_2476_nl, fsm_output[5]);
  assign nand_178_nl = ~((fsm_output[2]) & (fsm_output[8]) & (fsm_output[7]));
  assign mux_2309_nl = MUX_s_1_2_2(mux_tmp_2247, nand_178_nl, fsm_output[5]);
  assign mux_2311_nl = MUX_s_1_2_2(mux_2310_nl, mux_2309_nl, fsm_output[6]);
  assign mux_2307_nl = MUX_s_1_2_2(or_tmp_2324, or_tmp_2409, fsm_output[5]);
  assign mux_2306_nl = MUX_s_1_2_2(mux_tmp_2250, or_tmp_2406, fsm_output[5]);
  assign mux_2308_nl = MUX_s_1_2_2(mux_2307_nl, mux_2306_nl, fsm_output[6]);
  assign mux_2312_nl = MUX_s_1_2_2(mux_2311_nl, mux_2308_nl, fsm_output[4]);
  assign mux_2322_nl = MUX_s_1_2_2(mux_2321_nl, mux_2312_nl, fsm_output[3]);
  assign mux_2302_nl = MUX_s_1_2_2(or_tmp_2409, mux_tmp_2250, fsm_output[5]);
  assign mux_2300_nl = MUX_s_1_2_2(or_tmp_2406, or_2733_cse, fsm_output[5]);
  assign mux_2303_nl = MUX_s_1_2_2(mux_2302_nl, mux_2300_nl, fsm_output[6]);
  assign or_2468_nl = (fsm_output[5]) | mux_tmp_2247;
  assign mux_2299_nl = MUX_s_1_2_2(or_2468_nl, or_tmp_2395, fsm_output[6]);
  assign mux_2304_nl = MUX_s_1_2_2(mux_2303_nl, mux_2299_nl, fsm_output[4]);
  assign or_2461_nl = (fsm_output[5]) | (fsm_output[2]) | (~ (fsm_output[8])) | (fsm_output[7]);
  assign mux_2296_nl = MUX_s_1_2_2(mux_tmp_2244, or_2461_nl, fsm_output[6]);
  assign mux_2292_nl = MUX_s_1_2_2(or_tmp_2393, or_tmp_2391, fsm_output[1]);
  assign or_2455_nl = (~(and_515_cse | (fsm_output[2]))) | (fsm_output[8:7]!=2'b10);
  assign mux_2293_nl = MUX_s_1_2_2(mux_2292_nl, or_2455_nl, fsm_output[5]);
  assign mux_2294_nl = MUX_s_1_2_2(or_tmp_2395, mux_2293_nl, fsm_output[6]);
  assign mux_2297_nl = MUX_s_1_2_2(mux_2296_nl, mux_2294_nl, fsm_output[4]);
  assign mux_2305_nl = MUX_s_1_2_2(mux_2304_nl, mux_2297_nl, fsm_output[3]);
  assign mux_2323_nl = MUX_s_1_2_2(mux_2322_nl, mux_2305_nl, fsm_output[9]);
  assign nor_549_nl = ~((fsm_output[2]) | (fsm_output[5]) | (fsm_output[7]) | (fsm_output[8])
      | (fsm_output[9]));
  assign and_511_nl = (fsm_output[2]) & (fsm_output[5]) & (fsm_output[7]) & (fsm_output[8])
      & (fsm_output[9]);
  assign mux_2337_nl = MUX_s_1_2_2(nor_549_nl, and_511_nl, or_2500_cse);
  assign and_512_nl = (fsm_output[5]) & (fsm_output[7]) & (fsm_output[8]) & (fsm_output[9]);
  assign mux_2338_nl = MUX_s_1_2_2(mux_2337_nl, and_512_nl, or_602_cse);
  assign and_513_nl = (fsm_output[9:7]==3'b111);
  assign mux_2339_nl = MUX_s_1_2_2(mux_2338_nl, and_513_nl, fsm_output[6]);
  assign nor_548_nl = ~((fsm_output[8:1]!=8'b00000000));
  assign operator_64_false_or_2_nl = and_dcpl_290 | COMP_LOOP_10_modExp_dev_1_while_mul_mut_mx0c5
      | (~ mux_2336_itm);
  assign nor_524_nl = ~((fsm_output[8:4]!=5'b00000));
  assign mux_2427_nl = MUX_s_1_2_2(nor_524_nl, and_tmp_24, fsm_output[9]);
  assign and_331_nl = and_dcpl_239 & and_dcpl_106;
  assign COMP_LOOP_or_2_nl = (COMP_LOOP_COMP_LOOP_nor_itm & and_dcpl_240) | (COMP_LOOP_COMP_LOOP_and_14_itm
      & and_332_m1c) | (COMP_LOOP_COMP_LOOP_and_13_itm & and_334_m1c) | (COMP_LOOP_COMP_LOOP_and_12_itm
      & and_335_m1c) | (COMP_LOOP_COMP_LOOP_and_72_itm & and_338_m1c) | (COMP_LOOP_COMP_LOOP_and_10_itm
      & and_340_m1c) | (COMP_LOOP_COMP_LOOP_and_70_itm & and_342_m1c) | (COMP_LOOP_COMP_LOOP_and_69_itm
      & and_344_m1c) | (COMP_LOOP_COMP_LOOP_and_68_itm & and_346_m1c) | (COMP_LOOP_COMP_LOOP_and_6_itm
      & and_348_m1c) | (COMP_LOOP_COMP_LOOP_and_66_itm & and_350_m1c) | (COMP_LOOP_COMP_LOOP_and_65_itm
      & and_351_m1c) | (COMP_LOOP_COMP_LOOP_and_64_itm & and_352_m1c) | (COMP_LOOP_COMP_LOOP_and_185_itm
      & and_354_m1c) | (COMP_LOOP_COMP_LOOP_and_62_itm & and_356_m1c) | (COMP_LOOP_COMP_LOOP_and_244_itm
      & and_358_m1c);
  assign COMP_LOOP_or_3_nl = (COMP_LOOP_COMP_LOOP_and_244_itm & and_dcpl_240) | (COMP_LOOP_COMP_LOOP_nor_itm
      & and_332_m1c) | (COMP_LOOP_COMP_LOOP_and_14_itm & and_334_m1c) | (COMP_LOOP_COMP_LOOP_and_13_itm
      & and_335_m1c) | (COMP_LOOP_COMP_LOOP_and_12_itm & and_338_m1c) | (COMP_LOOP_COMP_LOOP_and_72_itm
      & and_340_m1c) | (COMP_LOOP_COMP_LOOP_and_10_itm & and_342_m1c) | (COMP_LOOP_COMP_LOOP_and_70_itm
      & and_344_m1c) | (COMP_LOOP_COMP_LOOP_and_69_itm & and_346_m1c) | (COMP_LOOP_COMP_LOOP_and_68_itm
      & and_348_m1c) | (COMP_LOOP_COMP_LOOP_and_6_itm & and_350_m1c) | (COMP_LOOP_COMP_LOOP_and_66_itm
      & and_351_m1c) | (COMP_LOOP_COMP_LOOP_and_65_itm & and_352_m1c) | (COMP_LOOP_COMP_LOOP_and_64_itm
      & and_354_m1c) | (COMP_LOOP_COMP_LOOP_and_185_itm & and_356_m1c) | (COMP_LOOP_COMP_LOOP_and_62_itm
      & and_358_m1c);
  assign COMP_LOOP_or_4_nl = (COMP_LOOP_COMP_LOOP_and_62_itm & and_dcpl_240) | (COMP_LOOP_COMP_LOOP_and_244_itm
      & and_332_m1c) | (COMP_LOOP_COMP_LOOP_nor_itm & and_334_m1c) | (COMP_LOOP_COMP_LOOP_and_14_itm
      & and_335_m1c) | (COMP_LOOP_COMP_LOOP_and_13_itm & and_338_m1c) | (COMP_LOOP_COMP_LOOP_and_12_itm
      & and_340_m1c) | (COMP_LOOP_COMP_LOOP_and_72_itm & and_342_m1c) | (COMP_LOOP_COMP_LOOP_and_10_itm
      & and_344_m1c) | (COMP_LOOP_COMP_LOOP_and_70_itm & and_346_m1c) | (COMP_LOOP_COMP_LOOP_and_69_itm
      & and_348_m1c) | (COMP_LOOP_COMP_LOOP_and_68_itm & and_350_m1c) | (COMP_LOOP_COMP_LOOP_and_6_itm
      & and_351_m1c) | (COMP_LOOP_COMP_LOOP_and_66_itm & and_352_m1c) | (COMP_LOOP_COMP_LOOP_and_65_itm
      & and_354_m1c) | (COMP_LOOP_COMP_LOOP_and_64_itm & and_356_m1c) | (COMP_LOOP_COMP_LOOP_and_185_itm
      & and_358_m1c);
  assign COMP_LOOP_or_5_nl = (COMP_LOOP_COMP_LOOP_and_185_itm & and_dcpl_240) | (COMP_LOOP_COMP_LOOP_and_62_itm
      & and_332_m1c) | (COMP_LOOP_COMP_LOOP_and_244_itm & and_334_m1c) | (COMP_LOOP_COMP_LOOP_nor_itm
      & and_335_m1c) | (COMP_LOOP_COMP_LOOP_and_14_itm & and_338_m1c) | (COMP_LOOP_COMP_LOOP_and_13_itm
      & and_340_m1c) | (COMP_LOOP_COMP_LOOP_and_12_itm & and_342_m1c) | (COMP_LOOP_COMP_LOOP_and_72_itm
      & and_344_m1c) | (COMP_LOOP_COMP_LOOP_and_10_itm & and_346_m1c) | (COMP_LOOP_COMP_LOOP_and_70_itm
      & and_348_m1c) | (COMP_LOOP_COMP_LOOP_and_69_itm & and_350_m1c) | (COMP_LOOP_COMP_LOOP_and_68_itm
      & and_351_m1c) | (COMP_LOOP_COMP_LOOP_and_6_itm & and_352_m1c) | (COMP_LOOP_COMP_LOOP_and_66_itm
      & and_354_m1c) | (COMP_LOOP_COMP_LOOP_and_65_itm & and_356_m1c) | (COMP_LOOP_COMP_LOOP_and_64_itm
      & and_358_m1c);
  assign COMP_LOOP_or_6_nl = (COMP_LOOP_COMP_LOOP_and_64_itm & and_dcpl_240) | (COMP_LOOP_COMP_LOOP_and_185_itm
      & and_332_m1c) | (COMP_LOOP_COMP_LOOP_and_62_itm & and_334_m1c) | (COMP_LOOP_COMP_LOOP_and_244_itm
      & and_335_m1c) | (COMP_LOOP_COMP_LOOP_nor_itm & and_338_m1c) | (COMP_LOOP_COMP_LOOP_and_14_itm
      & and_340_m1c) | (COMP_LOOP_COMP_LOOP_and_13_itm & and_342_m1c) | (COMP_LOOP_COMP_LOOP_and_12_itm
      & and_344_m1c) | (COMP_LOOP_COMP_LOOP_and_72_itm & and_346_m1c) | (COMP_LOOP_COMP_LOOP_and_10_itm
      & and_348_m1c) | (COMP_LOOP_COMP_LOOP_and_70_itm & and_350_m1c) | (COMP_LOOP_COMP_LOOP_and_69_itm
      & and_351_m1c) | (COMP_LOOP_COMP_LOOP_and_68_itm & and_352_m1c) | (COMP_LOOP_COMP_LOOP_and_6_itm
      & and_354_m1c) | (COMP_LOOP_COMP_LOOP_and_66_itm & and_356_m1c) | (COMP_LOOP_COMP_LOOP_and_65_itm
      & and_358_m1c);
  assign COMP_LOOP_or_7_nl = (COMP_LOOP_COMP_LOOP_and_65_itm & and_dcpl_240) | (COMP_LOOP_COMP_LOOP_and_64_itm
      & and_332_m1c) | (COMP_LOOP_COMP_LOOP_and_185_itm & and_334_m1c) | (COMP_LOOP_COMP_LOOP_and_62_itm
      & and_335_m1c) | (COMP_LOOP_COMP_LOOP_and_244_itm & and_338_m1c) | (COMP_LOOP_COMP_LOOP_nor_itm
      & and_340_m1c) | (COMP_LOOP_COMP_LOOP_and_14_itm & and_342_m1c) | (COMP_LOOP_COMP_LOOP_and_13_itm
      & and_344_m1c) | (COMP_LOOP_COMP_LOOP_and_12_itm & and_346_m1c) | (COMP_LOOP_COMP_LOOP_and_72_itm
      & and_348_m1c) | (COMP_LOOP_COMP_LOOP_and_10_itm & and_350_m1c) | (COMP_LOOP_COMP_LOOP_and_70_itm
      & and_351_m1c) | (COMP_LOOP_COMP_LOOP_and_69_itm & and_352_m1c) | (COMP_LOOP_COMP_LOOP_and_68_itm
      & and_354_m1c) | (COMP_LOOP_COMP_LOOP_and_6_itm & and_356_m1c) | (COMP_LOOP_COMP_LOOP_and_66_itm
      & and_358_m1c);
  assign COMP_LOOP_or_8_nl = (COMP_LOOP_COMP_LOOP_and_66_itm & and_dcpl_240) | (COMP_LOOP_COMP_LOOP_and_65_itm
      & and_332_m1c) | (COMP_LOOP_COMP_LOOP_and_64_itm & and_334_m1c) | (COMP_LOOP_COMP_LOOP_and_185_itm
      & and_335_m1c) | (COMP_LOOP_COMP_LOOP_and_62_itm & and_338_m1c) | (COMP_LOOP_COMP_LOOP_and_244_itm
      & and_340_m1c) | (COMP_LOOP_COMP_LOOP_nor_itm & and_342_m1c) | (COMP_LOOP_COMP_LOOP_and_14_itm
      & and_344_m1c) | (COMP_LOOP_COMP_LOOP_and_13_itm & and_346_m1c) | (COMP_LOOP_COMP_LOOP_and_12_itm
      & and_348_m1c) | (COMP_LOOP_COMP_LOOP_and_72_itm & and_350_m1c) | (COMP_LOOP_COMP_LOOP_and_10_itm
      & and_351_m1c) | (COMP_LOOP_COMP_LOOP_and_70_itm & and_352_m1c) | (COMP_LOOP_COMP_LOOP_and_69_itm
      & and_354_m1c) | (COMP_LOOP_COMP_LOOP_and_68_itm & and_356_m1c) | (COMP_LOOP_COMP_LOOP_and_6_itm
      & and_358_m1c);
  assign COMP_LOOP_or_9_nl = (COMP_LOOP_COMP_LOOP_and_6_itm & and_dcpl_240) | (COMP_LOOP_COMP_LOOP_and_66_itm
      & and_332_m1c) | (COMP_LOOP_COMP_LOOP_and_65_itm & and_334_m1c) | (COMP_LOOP_COMP_LOOP_and_64_itm
      & and_335_m1c) | (COMP_LOOP_COMP_LOOP_and_185_itm & and_338_m1c) | (COMP_LOOP_COMP_LOOP_and_62_itm
      & and_340_m1c) | (COMP_LOOP_COMP_LOOP_and_244_itm & and_342_m1c) | (COMP_LOOP_COMP_LOOP_nor_itm
      & and_344_m1c) | (COMP_LOOP_COMP_LOOP_and_14_itm & and_346_m1c) | (COMP_LOOP_COMP_LOOP_and_13_itm
      & and_348_m1c) | (COMP_LOOP_COMP_LOOP_and_12_itm & and_350_m1c) | (COMP_LOOP_COMP_LOOP_and_72_itm
      & and_351_m1c) | (COMP_LOOP_COMP_LOOP_and_10_itm & and_352_m1c) | (COMP_LOOP_COMP_LOOP_and_70_itm
      & and_354_m1c) | (COMP_LOOP_COMP_LOOP_and_69_itm & and_356_m1c) | (COMP_LOOP_COMP_LOOP_and_68_itm
      & and_358_m1c);
  assign COMP_LOOP_or_10_nl = (COMP_LOOP_COMP_LOOP_and_68_itm & and_dcpl_240) | (COMP_LOOP_COMP_LOOP_and_6_itm
      & and_332_m1c) | (COMP_LOOP_COMP_LOOP_and_66_itm & and_334_m1c) | (COMP_LOOP_COMP_LOOP_and_65_itm
      & and_335_m1c) | (COMP_LOOP_COMP_LOOP_and_64_itm & and_338_m1c) | (COMP_LOOP_COMP_LOOP_and_185_itm
      & and_340_m1c) | (COMP_LOOP_COMP_LOOP_and_62_itm & and_342_m1c) | (COMP_LOOP_COMP_LOOP_and_244_itm
      & and_344_m1c) | (COMP_LOOP_COMP_LOOP_nor_itm & and_346_m1c) | (COMP_LOOP_COMP_LOOP_and_14_itm
      & and_348_m1c) | (COMP_LOOP_COMP_LOOP_and_13_itm & and_350_m1c) | (COMP_LOOP_COMP_LOOP_and_12_itm
      & and_351_m1c) | (COMP_LOOP_COMP_LOOP_and_72_itm & and_352_m1c) | (COMP_LOOP_COMP_LOOP_and_10_itm
      & and_354_m1c) | (COMP_LOOP_COMP_LOOP_and_70_itm & and_356_m1c) | (COMP_LOOP_COMP_LOOP_and_69_itm
      & and_358_m1c);
  assign COMP_LOOP_or_11_nl = (COMP_LOOP_COMP_LOOP_and_69_itm & and_dcpl_240) | (COMP_LOOP_COMP_LOOP_and_68_itm
      & and_332_m1c) | (COMP_LOOP_COMP_LOOP_and_6_itm & and_334_m1c) | (COMP_LOOP_COMP_LOOP_and_66_itm
      & and_335_m1c) | (COMP_LOOP_COMP_LOOP_and_65_itm & and_338_m1c) | (COMP_LOOP_COMP_LOOP_and_64_itm
      & and_340_m1c) | (COMP_LOOP_COMP_LOOP_and_185_itm & and_342_m1c) | (COMP_LOOP_COMP_LOOP_and_62_itm
      & and_344_m1c) | (COMP_LOOP_COMP_LOOP_and_244_itm & and_346_m1c) | (COMP_LOOP_COMP_LOOP_nor_itm
      & and_348_m1c) | (COMP_LOOP_COMP_LOOP_and_14_itm & and_350_m1c) | (COMP_LOOP_COMP_LOOP_and_13_itm
      & and_351_m1c) | (COMP_LOOP_COMP_LOOP_and_12_itm & and_352_m1c) | (COMP_LOOP_COMP_LOOP_and_72_itm
      & and_354_m1c) | (COMP_LOOP_COMP_LOOP_and_10_itm & and_356_m1c) | (COMP_LOOP_COMP_LOOP_and_70_itm
      & and_358_m1c);
  assign COMP_LOOP_or_12_nl = (COMP_LOOP_COMP_LOOP_and_70_itm & and_dcpl_240) | (COMP_LOOP_COMP_LOOP_and_69_itm
      & and_332_m1c) | (COMP_LOOP_COMP_LOOP_and_68_itm & and_334_m1c) | (COMP_LOOP_COMP_LOOP_and_6_itm
      & and_335_m1c) | (COMP_LOOP_COMP_LOOP_and_66_itm & and_338_m1c) | (COMP_LOOP_COMP_LOOP_and_65_itm
      & and_340_m1c) | (COMP_LOOP_COMP_LOOP_and_64_itm & and_342_m1c) | (COMP_LOOP_COMP_LOOP_and_185_itm
      & and_344_m1c) | (COMP_LOOP_COMP_LOOP_and_62_itm & and_346_m1c) | (COMP_LOOP_COMP_LOOP_and_244_itm
      & and_348_m1c) | (COMP_LOOP_COMP_LOOP_nor_itm & and_350_m1c) | (COMP_LOOP_COMP_LOOP_and_14_itm
      & and_351_m1c) | (COMP_LOOP_COMP_LOOP_and_13_itm & and_352_m1c) | (COMP_LOOP_COMP_LOOP_and_12_itm
      & and_354_m1c) | (COMP_LOOP_COMP_LOOP_and_72_itm & and_356_m1c) | (COMP_LOOP_COMP_LOOP_and_10_itm
      & and_358_m1c);
  assign COMP_LOOP_or_13_nl = (COMP_LOOP_COMP_LOOP_and_10_itm & and_dcpl_240) | (COMP_LOOP_COMP_LOOP_and_70_itm
      & and_332_m1c) | (COMP_LOOP_COMP_LOOP_and_69_itm & and_334_m1c) | (COMP_LOOP_COMP_LOOP_and_68_itm
      & and_335_m1c) | (COMP_LOOP_COMP_LOOP_and_6_itm & and_338_m1c) | (COMP_LOOP_COMP_LOOP_and_66_itm
      & and_340_m1c) | (COMP_LOOP_COMP_LOOP_and_65_itm & and_342_m1c) | (COMP_LOOP_COMP_LOOP_and_64_itm
      & and_344_m1c) | (COMP_LOOP_COMP_LOOP_and_185_itm & and_346_m1c) | (COMP_LOOP_COMP_LOOP_and_62_itm
      & and_348_m1c) | (COMP_LOOP_COMP_LOOP_and_244_itm & and_350_m1c) | (COMP_LOOP_COMP_LOOP_nor_itm
      & and_351_m1c) | (COMP_LOOP_COMP_LOOP_and_14_itm & and_352_m1c) | (COMP_LOOP_COMP_LOOP_and_13_itm
      & and_354_m1c) | (COMP_LOOP_COMP_LOOP_and_12_itm & and_356_m1c) | (COMP_LOOP_COMP_LOOP_and_72_itm
      & and_358_m1c);
  assign COMP_LOOP_or_14_nl = (COMP_LOOP_COMP_LOOP_and_72_itm & and_dcpl_240) | (COMP_LOOP_COMP_LOOP_and_10_itm
      & and_332_m1c) | (COMP_LOOP_COMP_LOOP_and_70_itm & and_334_m1c) | (COMP_LOOP_COMP_LOOP_and_69_itm
      & and_335_m1c) | (COMP_LOOP_COMP_LOOP_and_68_itm & and_338_m1c) | (COMP_LOOP_COMP_LOOP_and_6_itm
      & and_340_m1c) | (COMP_LOOP_COMP_LOOP_and_66_itm & and_342_m1c) | (COMP_LOOP_COMP_LOOP_and_65_itm
      & and_344_m1c) | (COMP_LOOP_COMP_LOOP_and_64_itm & and_346_m1c) | (COMP_LOOP_COMP_LOOP_and_185_itm
      & and_348_m1c) | (COMP_LOOP_COMP_LOOP_and_62_itm & and_350_m1c) | (COMP_LOOP_COMP_LOOP_and_244_itm
      & and_351_m1c) | (COMP_LOOP_COMP_LOOP_nor_itm & and_352_m1c) | (COMP_LOOP_COMP_LOOP_and_14_itm
      & and_354_m1c) | (COMP_LOOP_COMP_LOOP_and_13_itm & and_356_m1c) | (COMP_LOOP_COMP_LOOP_and_12_itm
      & and_358_m1c);
  assign COMP_LOOP_or_15_nl = (COMP_LOOP_COMP_LOOP_and_12_itm & and_dcpl_240) | (COMP_LOOP_COMP_LOOP_and_72_itm
      & and_332_m1c) | (COMP_LOOP_COMP_LOOP_and_10_itm & and_334_m1c) | (COMP_LOOP_COMP_LOOP_and_70_itm
      & and_335_m1c) | (COMP_LOOP_COMP_LOOP_and_69_itm & and_338_m1c) | (COMP_LOOP_COMP_LOOP_and_68_itm
      & and_340_m1c) | (COMP_LOOP_COMP_LOOP_and_6_itm & and_342_m1c) | (COMP_LOOP_COMP_LOOP_and_66_itm
      & and_344_m1c) | (COMP_LOOP_COMP_LOOP_and_65_itm & and_346_m1c) | (COMP_LOOP_COMP_LOOP_and_64_itm
      & and_348_m1c) | (COMP_LOOP_COMP_LOOP_and_185_itm & and_350_m1c) | (COMP_LOOP_COMP_LOOP_and_62_itm
      & and_351_m1c) | (COMP_LOOP_COMP_LOOP_and_244_itm & and_352_m1c) | (COMP_LOOP_COMP_LOOP_nor_itm
      & and_354_m1c) | (COMP_LOOP_COMP_LOOP_and_14_itm & and_356_m1c) | (COMP_LOOP_COMP_LOOP_and_13_itm
      & and_358_m1c);
  assign COMP_LOOP_or_16_nl = (COMP_LOOP_COMP_LOOP_and_13_itm & and_dcpl_240) | (COMP_LOOP_COMP_LOOP_and_12_itm
      & and_332_m1c) | (COMP_LOOP_COMP_LOOP_and_72_itm & and_334_m1c) | (COMP_LOOP_COMP_LOOP_and_10_itm
      & and_335_m1c) | (COMP_LOOP_COMP_LOOP_and_70_itm & and_338_m1c) | (COMP_LOOP_COMP_LOOP_and_69_itm
      & and_340_m1c) | (COMP_LOOP_COMP_LOOP_and_68_itm & and_342_m1c) | (COMP_LOOP_COMP_LOOP_and_6_itm
      & and_344_m1c) | (COMP_LOOP_COMP_LOOP_and_66_itm & and_346_m1c) | (COMP_LOOP_COMP_LOOP_and_65_itm
      & and_348_m1c) | (COMP_LOOP_COMP_LOOP_and_64_itm & and_350_m1c) | (COMP_LOOP_COMP_LOOP_and_185_itm
      & and_351_m1c) | (COMP_LOOP_COMP_LOOP_and_62_itm & and_352_m1c) | (COMP_LOOP_COMP_LOOP_and_244_itm
      & and_354_m1c) | (COMP_LOOP_COMP_LOOP_nor_itm & and_356_m1c) | (COMP_LOOP_COMP_LOOP_and_14_itm
      & and_358_m1c);
  assign COMP_LOOP_or_17_nl = (COMP_LOOP_COMP_LOOP_and_14_itm & and_dcpl_240) | (COMP_LOOP_COMP_LOOP_and_13_itm
      & and_332_m1c) | (COMP_LOOP_COMP_LOOP_and_12_itm & and_334_m1c) | (COMP_LOOP_COMP_LOOP_and_72_itm
      & and_335_m1c) | (COMP_LOOP_COMP_LOOP_and_10_itm & and_338_m1c) | (COMP_LOOP_COMP_LOOP_and_70_itm
      & and_340_m1c) | (COMP_LOOP_COMP_LOOP_and_69_itm & and_342_m1c) | (COMP_LOOP_COMP_LOOP_and_68_itm
      & and_344_m1c) | (COMP_LOOP_COMP_LOOP_and_6_itm & and_346_m1c) | (COMP_LOOP_COMP_LOOP_and_66_itm
      & and_348_m1c) | (COMP_LOOP_COMP_LOOP_and_65_itm & and_350_m1c) | (COMP_LOOP_COMP_LOOP_and_64_itm
      & and_351_m1c) | (COMP_LOOP_COMP_LOOP_and_185_itm & and_352_m1c) | (COMP_LOOP_COMP_LOOP_and_62_itm
      & and_354_m1c) | (COMP_LOOP_COMP_LOOP_and_244_itm & and_356_m1c) | (COMP_LOOP_COMP_LOOP_nor_itm
      & and_358_m1c);
  assign mux_2470_nl = MUX_s_1_2_2(and_dcpl_146, or_tmp_33, and_516_cse);
  assign mux_2471_nl = MUX_s_1_2_2((~ mux_2470_nl), and_711_cse, fsm_output[5]);
  assign or_2622_nl = (~ (fsm_output[2])) | (fsm_output[6]) | (fsm_output[3]);
  assign mux_2469_nl = MUX_s_1_2_2(or_2622_nl, or_307_cse, fsm_output[1]);
  assign or_2623_nl = (fsm_output[5]) | (~ mux_2469_nl);
  assign mux_2472_nl = MUX_s_1_2_2(mux_2471_nl, or_2623_nl, fsm_output[4]);
  assign mux_2465_nl = MUX_s_1_2_2(and_dcpl_146, (fsm_output[3]), fsm_output[2]);
  assign mux_2464_nl = MUX_s_1_2_2(and_dcpl_146, or_tmp_33, fsm_output[2]);
  assign mux_2466_nl = MUX_s_1_2_2(mux_2465_nl, mux_2464_nl, fsm_output[1]);
  assign mux_2467_nl = MUX_s_1_2_2((~ mux_2466_nl), nor_tmp_403, fsm_output[5]);
  assign mux_2468_nl = MUX_s_1_2_2(mux_2467_nl, or_tmp_2551, fsm_output[4]);
  assign mux_2473_nl = MUX_s_1_2_2(mux_2472_nl, mux_2468_nl, fsm_output[0]);
  assign mux_2461_nl = MUX_s_1_2_2((~ nor_tmp_399), nor_tmp_403, fsm_output[5]);
  assign mux_2462_nl = MUX_s_1_2_2((~ or_tmp_2552), mux_2461_nl, fsm_output[4]);
  assign mux_2463_nl = MUX_s_1_2_2(mux_tmp_2389, mux_2462_nl, fsm_output[0]);
  assign mux_2474_nl = MUX_s_1_2_2(mux_2473_nl, (~ mux_2463_nl), fsm_output[7]);
  assign or_2621_nl = (fsm_output[5]) | (~ or_tmp_2549);
  assign mux_2458_nl = MUX_s_1_2_2(mux_tmp_2381, or_2621_nl, fsm_output[4]);
  assign mux_2459_nl = MUX_s_1_2_2(mux_tmp_2382, mux_2458_nl, fsm_output[0]);
  assign mux_2455_nl = MUX_s_1_2_2(or_tmp_2439, (~ or_307_cse), fsm_output[5]);
  assign mux_2454_nl = MUX_s_1_2_2((~ nor_tmp_1), nor_tmp_403, fsm_output[5]);
  assign mux_2456_nl = MUX_s_1_2_2(mux_2455_nl, mux_2454_nl, fsm_output[4]);
  assign mux_2452_nl = MUX_s_1_2_2((~ nor_tmp_1), mux_tmp_2400, fsm_output[5]);
  assign mux_2453_nl = MUX_s_1_2_2((~ mux_tmp_2380), mux_2452_nl, fsm_output[4]);
  assign mux_2457_nl = MUX_s_1_2_2(mux_2456_nl, mux_2453_nl, fsm_output[0]);
  assign mux_2460_nl = MUX_s_1_2_2((~ mux_2459_nl), mux_2457_nl, fsm_output[7]);
  assign mux_2475_nl = MUX_s_1_2_2(mux_2474_nl, mux_2460_nl, fsm_output[8]);
  assign mux_2446_nl = MUX_s_1_2_2(not_tmp_617, nor_tmp_399, fsm_output[5]);
  assign mux_2447_nl = MUX_s_1_2_2(mux_2446_nl, or_tmp_2552, fsm_output[4]);
  assign mux_2444_nl = MUX_s_1_2_2(not_tmp_617, and_711_cse, fsm_output[5]);
  assign mux_2445_nl = MUX_s_1_2_2(mux_2444_nl, or_tmp_2551, fsm_output[4]);
  assign mux_2448_nl = MUX_s_1_2_2(mux_2447_nl, mux_2445_nl, fsm_output[0]);
  assign mux_2441_nl = MUX_s_1_2_2(and_dcpl_95, or_tmp_2549, fsm_output[5]);
  assign mux_2442_nl = MUX_s_1_2_2((~ mux_2441_nl), mux_tmp_2381, fsm_output[4]);
  assign mux_2443_nl = MUX_s_1_2_2(mux_2442_nl, mux_tmp_2389, fsm_output[0]);
  assign mux_2449_nl = MUX_s_1_2_2(mux_2448_nl, (~ mux_2443_nl), fsm_output[7]);
  assign mux_2434_nl = MUX_s_1_2_2(not_tmp_617, nor_tmp_1, fsm_output[5]);
  assign mux_2435_nl = MUX_s_1_2_2(mux_2434_nl, mux_tmp_2380, fsm_output[4]);
  assign mux_2436_nl = MUX_s_1_2_2(mux_2435_nl, mux_tmp_2382, fsm_output[0]);
  assign mux_2437_nl = MUX_s_1_2_2((~ mux_2436_nl), or_tmp_2548, fsm_output[7]);
  assign mux_2450_nl = MUX_s_1_2_2(mux_2449_nl, mux_2437_nl, fsm_output[8]);
  assign COMP_LOOP_COMP_LOOP_and_17_nl = (COMP_LOOP_1_operator_64_false_acc_tmp[3:0]==4'b0011);
  assign modExp_dev_while_or_nl = and_dcpl_290 | (~ mux_2336_itm);
  assign modExp_dev_while_or_1_nl = COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c3
      | COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c4 | COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c5
      | COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c6 | COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c7
      | COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c8 | COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c9
      | COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c10 |
      COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c11 | COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c12
      | COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c13;
  assign nand_486_nl = ~(and_dcpl_294 & and_dcpl_346);
  assign nor_nl = ~((fsm_output[1]) | (fsm_output[7]) | (~ (fsm_output[0])) | (~
      (fsm_output[4])) | (fsm_output[9]) | (fsm_output[8]));
  assign nor_1038_nl = ~((~ (fsm_output[1])) | (~ (fsm_output[7])) | (fsm_output[0])
      | (fsm_output[4]) | nand_490_cse);
  assign mux_2864_nl = MUX_s_1_2_2(nor_nl, nor_1038_nl, fsm_output[2]);
  assign and_421_nl = and_dcpl_109 & and_dcpl_346;
  assign and_422_nl = and_dcpl_239 & and_dcpl_256;
  assign and_423_nl = and_dcpl_244 & and_dcpl_307;
  assign and_424_nl = and_dcpl_248 & and_dcpl_263;
  assign and_425_nl = and_dcpl_253 & and_dcpl_260;
  assign and_426_nl = and_dcpl_257 & and_dcpl_313;
  assign and_427_nl = and_dcpl_261 & and_dcpl_319;
  assign and_428_nl = and_dcpl_264 & and_dcpl_317;
  assign and_429_nl = and_dcpl_268 & and_dcpl_323;
  assign and_430_nl = and_dcpl_244 & and_dcpl_321;
  assign and_431_nl = and_dcpl_239 & and_dcpl_284;
  assign and_432_nl = and_dcpl_275 & and_dcpl_279;
  assign and_433_nl = and_dcpl_248 & and_dcpl_288;
  assign and_434_nl = and_dcpl_282 & and_dcpl_331;
  assign operator_64_false_mux1h_nl = MUX1HOT_v_4_16_2((z_out_3[3:0]), (COMP_LOOP_acc_psp_sva[3:0]),
      4'b0001, 4'b0010, 4'b0011, 4'b0100, 4'b0101, 4'b0110, 4'b0111, 4'b1000, 4'b1001,
      4'b1010, 4'b1011, 4'b1100, 4'b1101, 4'b1110, {(~ mux_2336_itm) , (~ mux_2797_itm)
      , and_421_nl , and_422_nl , and_423_nl , and_424_nl , and_425_nl , and_426_nl
      , and_427_nl , and_428_nl , and_429_nl , and_430_nl , and_431_nl , and_432_nl
      , and_433_nl , and_434_nl});
  assign COMP_LOOP_nand_nl = ~(and_dcpl_268 & and_dcpl_106);
  assign operator_64_false_and_nl = MUX_v_4_2_2(4'b0000, operator_64_false_mux1h_nl,
      COMP_LOOP_nand_nl);
  assign and_435_nl = and_dcpl_257 & and_dcpl_329;
  assign operator_64_false_or_2_nl_1 = MUX_v_4_2_2(operator_64_false_and_nl, 4'b1111,
      and_435_nl);
  assign nl_operator_64_false_1_acc_nl = ({1'b1 , (~ COMP_LOOP_k_9_4_sva_4_0)}) +
      6'b000001;
  assign operator_64_false_1_acc_nl = nl_operator_64_false_1_acc_nl[5:0];
  assign mux_2587_nl = MUX_s_1_2_2(or_tmp_2548, or_tmp, fsm_output[0]);
  assign or_2696_nl = (fsm_output[7]) | mux_2587_nl;
  assign mux_2590_nl = MUX_s_1_2_2(not_tmp_664, or_2696_nl, fsm_output[8]);
  assign or_2699_nl = (fsm_output[5:4]!=2'b00);
  assign mux_2591_nl = MUX_s_1_2_2(nor_tmp_1, (fsm_output[6]), or_2699_nl);
  assign mux_2592_nl = MUX_s_1_2_2(mux_tmp_2538, (~ mux_2591_nl), fsm_output[7]);
  assign mux_2597_nl = MUX_s_1_2_2(mux_tmp_2468, (fsm_output[6]), fsm_output[5]);
  assign mux_2598_nl = MUX_s_1_2_2(mux_156_cse, mux_2597_nl, fsm_output[4]);
  assign mux_2593_nl = MUX_s_1_2_2(and_dcpl_95, and_711_cse, or_2700_cse);
  assign mux_2594_nl = MUX_s_1_2_2(mux_2593_nl, (fsm_output[6]), fsm_output[5]);
  assign mux_2596_nl = MUX_s_1_2_2(mux_156_cse, mux_2594_nl, fsm_output[4]);
  assign mux_2599_nl = MUX_s_1_2_2(mux_2598_nl, mux_2596_nl, fsm_output[0]);
  assign or_2701_nl = (fsm_output[6:1]!=6'b000000);
  assign mux_2600_nl = MUX_s_1_2_2(or_tmp, or_2701_nl, fsm_output[0]);
  assign mux_2601_nl = MUX_s_1_2_2(mux_tmp_2538, (~ mux_2600_nl), fsm_output[7]);
  assign nl_COMP_LOOP_acc_7_psp_sva  = (STAGE_VEC_LOOP_j_sva_9_0[9:1]) + conv_u2u_8_9({COMP_LOOP_k_9_4_sva_4_0
      , 3'b001});
  assign and_485_nl = (fsm_output[4]) & (fsm_output[5]) & (fsm_output[2]);
  assign mux_2611_nl = MUX_s_1_2_2((fsm_output[6]), or_165_cse, and_485_nl);
  assign mux_2612_nl = MUX_s_1_2_2(mux_tmp_2538, (~ mux_2611_nl), fsm_output[7]);
  assign or_2824_nl = (fsm_output[7:5]!=3'b000);
  assign or_2825_nl = and_515_cse | (fsm_output[7:5]!=3'b000);
  assign nand_161_nl = ~(or_2500_cse & (fsm_output[7:5]==3'b111));
  assign mux_2614_nl = MUX_s_1_2_2(or_2825_nl, nand_161_nl, fsm_output[2]);
  assign nand_162_nl = ~((fsm_output[7:5]==3'b111));
  assign mux_2615_nl = MUX_s_1_2_2(mux_2614_nl, nand_162_nl, fsm_output[3]);
  assign mux_2616_nl = MUX_s_1_2_2(or_2824_nl, mux_2615_nl, fsm_output[4]);
  assign and_482_nl = (fsm_output[5]) & (fsm_output[1]) & (fsm_output[2]);
  assign mux_2619_nl = MUX_s_1_2_2((fsm_output[6]), or_165_cse, and_482_nl);
  assign mux_2620_nl = MUX_s_1_2_2(mux_2619_nl, or_420_cse, fsm_output[4]);
  assign or_2707_nl = (fsm_output[7]) | mux_2620_nl;
  assign mux_2621_nl = MUX_s_1_2_2(not_tmp_664, or_2707_nl, fsm_output[8]);
  assign and_480_nl = (fsm_output[4]) & (fsm_output[5]) & (fsm_output[1]) & (fsm_output[2]);
  assign mux_2623_nl = MUX_s_1_2_2((fsm_output[6]), or_165_cse, and_480_nl);
  assign or_2708_nl = (fsm_output[7]) | mux_2623_nl;
  assign mux_2624_nl = MUX_s_1_2_2(not_tmp_664, or_2708_nl, fsm_output[8]);
  assign mux_2629_nl = MUX_s_1_2_2(mux_tmp_2574, and_475_cse, fsm_output[2]);
  assign mux_2630_nl = MUX_s_1_2_2(nor_510_cse, mux_2629_nl, fsm_output[4]);
  assign mux_2627_nl = MUX_s_1_2_2(nor_510_cse, mux_tmp_2574, fsm_output[2]);
  assign mux_2628_nl = MUX_s_1_2_2(mux_2627_nl, and_475_cse, fsm_output[4]);
  assign mux_2631_nl = MUX_s_1_2_2(mux_2630_nl, mux_2628_nl, and_515_cse);
  assign mux_2626_nl = MUX_s_1_2_2(mux_tmp_2574, and_475_cse, fsm_output[4]);
  assign mux_2632_nl = MUX_s_1_2_2(mux_2631_nl, mux_2626_nl, fsm_output[3]);
  assign mux_2633_nl = MUX_s_1_2_2(mux_2632_nl, (fsm_output[8]), fsm_output[7]);
  assign nl_COMP_LOOP_acc_9_psp_sva  = (STAGE_VEC_LOOP_j_sva_9_0[9:1]) + conv_u2u_8_9({COMP_LOOP_k_9_4_sva_4_0
      , 3'b011});
  assign nor_511_nl = ~((fsm_output[2]) | (fsm_output[5]) | (fsm_output[6]) | (fsm_output[8]));
  assign and_473_nl = (fsm_output[2]) & (fsm_output[5]) & (fsm_output[6]) & (fsm_output[8]);
  assign mux_2637_nl = MUX_s_1_2_2(nor_511_nl, and_473_nl, and_515_cse);
  assign mux_2638_nl = MUX_s_1_2_2(mux_2637_nl, and_475_cse, fsm_output[3]);
  assign mux_2639_nl = MUX_s_1_2_2(nor_510_cse, mux_2638_nl, fsm_output[4]);
  assign mux_2640_nl = MUX_s_1_2_2(mux_2639_nl, (fsm_output[8]), fsm_output[7]);
  assign and_393_nl = (fsm_output[7]) & or_420_cse;
  assign mux_2641_nl = MUX_s_1_2_2(not_tmp_664, and_393_nl, fsm_output[8]);
  assign nl_COMP_LOOP_acc_cse_8_sva  = STAGE_VEC_LOOP_j_sva_9_0 + conv_u2u_9_10({COMP_LOOP_k_9_4_sva_4_0
      , 4'b0111});
  assign and_397_nl = (fsm_output[7]) & or_tmp_2638;
  assign mux_2645_nl = MUX_s_1_2_2(not_tmp_664, and_397_nl, fsm_output[8]);
  assign nor_937_nl = ~(and_515_cse | (fsm_output[8:6]!=3'b000));
  assign and_754_nl = or_2500_cse & (fsm_output[8:6]==3'b111);
  assign mux_2646_nl = MUX_s_1_2_2(nor_937_nl, and_754_nl, fsm_output[3]);
  assign and_755_nl = (fsm_output[3]) & (fsm_output[6]) & (fsm_output[7]) & (fsm_output[8]);
  assign mux_2647_nl = MUX_s_1_2_2(mux_2646_nl, and_755_nl, fsm_output[2]);
  assign mux_2648_nl = MUX_s_1_2_2(nor_936_cse, mux_2647_nl, fsm_output[4]);
  assign mux_2649_nl = MUX_s_1_2_2(mux_2648_nl, and_756_cse, fsm_output[5]);
  assign nl_COMP_LOOP_acc_10_psp_sva  = (STAGE_VEC_LOOP_j_sva_9_0[9:3]) + conv_u2u_6_7({COMP_LOOP_k_9_4_sva_4_0
      , 1'b1});
  assign or_196_nl = (fsm_output[2:0]!=3'b000);
  assign mux_2655_nl = MUX_s_1_2_2(not_tmp_696, mux_tmp_302, or_196_nl);
  assign mux_2656_nl = MUX_s_1_2_2(not_tmp_696, mux_2655_nl, fsm_output[3]);
  assign mux_2653_nl = MUX_s_1_2_2(mux_tmp_302, nor_tmp_87, and_515_cse);
  assign mux_2654_nl = MUX_s_1_2_2(mux_2653_nl, nor_tmp_87, or_598_cse);
  assign mux_2657_nl = MUX_s_1_2_2(mux_2656_nl, mux_2654_nl, fsm_output[4]);
  assign or_2651_nl = (fsm_output[8:7]!=2'b00) | mux_tmp_2377;
  assign nl_COMP_LOOP_acc_cse_10_sva  = STAGE_VEC_LOOP_j_sva_9_0 + conv_u2u_9_10({COMP_LOOP_k_9_4_sva_4_0
      , 4'b1001});
  assign or_2732_nl = (fsm_output[8:7]!=2'b00) | mux_tmp_2450;
  assign mux_2666_nl = MUX_s_1_2_2(mux_tmp_2612, nor_tmp_3, fsm_output[3]);
  assign mux_2667_nl = MUX_s_1_2_2(not_tmp_703, mux_2666_nl, fsm_output[4]);
  assign mux_2668_nl = MUX_s_1_2_2(mux_2667_nl, mux_tmp_2614, and_515_cse);
  assign mux_2669_nl = MUX_s_1_2_2(mux_2668_nl, mux_tmp_2614, fsm_output[2]);
  assign mux_2670_nl = MUX_s_1_2_2(mux_2669_nl, nor_tmp_3, fsm_output[5]);
  assign nl_COMP_LOOP_acc_11_psp_sva  = (STAGE_VEC_LOOP_j_sva_9_0[9:1]) + conv_u2u_8_9({COMP_LOOP_k_9_4_sva_4_0
      , 3'b101});
  assign mux_2678_nl = MUX_s_1_2_2(mux_tmp_2626, and_tmp_11, fsm_output[3]);
  assign mux_2679_nl = MUX_s_1_2_2(mux_2678_nl, mux_tmp_2625, and_515_cse);
  assign mux_2680_nl = MUX_s_1_2_2(mux_2679_nl, mux_tmp_2625, fsm_output[2]);
  assign mux_2681_nl = MUX_s_1_2_2(mux_tmp_2626, mux_2680_nl, fsm_output[4]);
  assign or_2743_nl = (fsm_output[8]) | ((fsm_output[7]) & or_tmp);
  assign nl_COMP_LOOP_acc_cse_12_sva  = STAGE_VEC_LOOP_j_sva_9_0 + conv_u2u_9_10({COMP_LOOP_k_9_4_sva_4_0
      , 4'b1011});
  assign or_2748_nl = (fsm_output[8]) | ((fsm_output[7]) & mux_tmp_79);
  assign nor_503_nl = ~((fsm_output[5]) | (fsm_output[7]) | (fsm_output[9]));
  assign nor_504_nl = ~((fsm_output[3]) | and_515_cse | (fsm_output[5]) | (fsm_output[7])
      | (fsm_output[9]));
  assign and_409_nl = (fsm_output[3]) & or_2500_cse & (fsm_output[5]) & (fsm_output[7])
      & (fsm_output[9]);
  assign mux_2690_nl = MUX_s_1_2_2(nor_504_nl, and_409_nl, fsm_output[2]);
  assign mux_2691_nl = MUX_s_1_2_2(nor_503_nl, mux_2690_nl, fsm_output[4]);
  assign mux_2692_nl = MUX_s_1_2_2(mux_2691_nl, and_459_cse, fsm_output[6]);
  assign nor_500_nl = ~((fsm_output[6]) | (fsm_output[7]) | (fsm_output[9]));
  assign and_452_nl = or_2500_cse & (fsm_output[3:2]==2'b11);
  assign mux_2706_nl = MUX_s_1_2_2(nor_500_nl, mux_tmp_2653, and_452_nl);
  assign or_2755_nl = and_515_cse | (fsm_output[3:2]!=2'b00);
  assign mux_2705_nl = MUX_s_1_2_2(mux_tmp_2653, nor_tmp_459, or_2755_nl);
  assign mux_2707_nl = MUX_s_1_2_2(mux_2706_nl, mux_2705_nl, fsm_output[4]);
  assign mux_2708_nl = MUX_s_1_2_2(mux_2707_nl, nor_tmp_459, fsm_output[5]);
  assign nor_498_nl = ~((fsm_output[2]) | (fsm_output[5]) | (fsm_output[6]) | (fsm_output[7])
      | (fsm_output[9]));
  assign nor_499_nl = ~((fsm_output[0]) | (fsm_output[5]) | (fsm_output[6]) | (fsm_output[7])
      | (fsm_output[9]));
  assign mux_2710_nl = MUX_s_1_2_2(nor_499_nl, nor_tmp_463, fsm_output[2]);
  assign mux_2711_nl = MUX_s_1_2_2(nor_498_nl, mux_2710_nl, fsm_output[1]);
  assign mux_2712_nl = MUX_s_1_2_2(mux_2711_nl, nor_tmp_463, fsm_output[3]);
  assign mux_2713_nl = MUX_s_1_2_2(nor_497_cse, mux_2712_nl, fsm_output[4]);
  assign nl_COMP_LOOP_acc_cse_14_sva  = STAGE_VEC_LOOP_j_sva_9_0 + conv_u2u_9_10({COMP_LOOP_k_9_4_sva_4_0
      , 4'b1101});
  assign and_410_nl = (fsm_output[8]) & ((fsm_output[7]) | (fsm_output[4]) | (fsm_output[5])
      | or_tmp_2439);
  assign mux_2720_nl = MUX_s_1_2_2(mux_tmp_2666, nor_tmp_467, or_598_cse);
  assign mux_2721_nl = MUX_s_1_2_2(not_tmp_729, mux_2720_nl, fsm_output[4]);
  assign and_636_nl = (fsm_output[3:2]==2'b11);
  assign mux_2718_nl = MUX_s_1_2_2(not_tmp_729, mux_tmp_2666, and_636_nl);
  assign mux_2719_nl = MUX_s_1_2_2(mux_2718_nl, nor_tmp_467, fsm_output[4]);
  assign mux_2722_nl = MUX_s_1_2_2(mux_2721_nl, mux_2719_nl, and_515_cse);
  assign nl_COMP_LOOP_acc_13_psp_sva  = (STAGE_VEC_LOOP_j_sva_9_0[9:1]) + conv_u2u_8_9({COMP_LOOP_k_9_4_sva_4_0
      , 3'b111});
  assign or_2814_nl = (fsm_output[5]) | (fsm_output[8]) | (fsm_output[9]);
  assign or_2815_nl = (fsm_output[2]) | (fsm_output[3]) | (fsm_output[5]) | (fsm_output[8])
      | (fsm_output[9]);
  assign nand_156_nl = ~((fsm_output[2]) & (fsm_output[3]) & (fsm_output[5]) & (fsm_output[8])
      & (fsm_output[9]));
  assign mux_2728_nl = MUX_s_1_2_2(or_2815_nl, nand_156_nl, and_515_cse);
  assign mux_2729_nl = MUX_s_1_2_2(or_2814_nl, mux_2728_nl, fsm_output[4]);
  assign mux_2730_nl = MUX_s_1_2_2(mux_2729_nl, nand_490_cse, or_111_cse);
  assign or_411_nl = (fsm_output[9:8]!=2'b00);
  assign or_2777_nl = (fsm_output[2]) | and_515_cse | (fsm_output[3]) | (fsm_output[8])
      | (fsm_output[9]);
  assign mux_2731_nl = MUX_s_1_2_2(or_411_nl, or_2777_nl, fsm_output[4]);
  assign or_2812_nl = (fsm_output[6]) | mux_2731_nl;
  assign nand_154_nl = ~((fsm_output[6]) & or_602_cse & (fsm_output[9:8]==2'b11));
  assign mux_2732_nl = MUX_s_1_2_2(or_2812_nl, nand_154_nl, fsm_output[5]);
  assign mux_2733_nl = MUX_s_1_2_2(mux_2732_nl, nand_490_cse, fsm_output[7]);
  assign nl_COMP_LOOP_acc_cse_sva  = STAGE_VEC_LOOP_j_sva_9_0 + conv_u2u_9_10({COMP_LOOP_k_9_4_sva_4_0
      , 4'b1111});
  assign and_413_nl = (fsm_output[8]) & ((fsm_output[7]) | nor_tmp_427);
  assign or_2891_nl = (fsm_output[0]) | (fsm_output[4]);
  assign mux_2736_nl = MUX_s_1_2_2(mux_tmp_2449, or_420_cse, or_2891_nl);
  assign and_414_nl = (fsm_output[8:7]==2'b11) & mux_2736_nl;
  assign COMP_LOOP_nor_11_nl = ~((COMP_LOOP_1_operator_64_false_acc_tmp[3:1]!=3'b000));
  assign COMP_LOOP_or_35_nl = operator_64_false_slc_operator_64_false_acc_1_60_itm_mx0c1
      | operator_64_false_slc_operator_64_false_acc_1_60_itm_mx0c3;
  assign COMP_LOOP_or_18_nl = (COMP_LOOP_COMP_LOOP_nor_1_itm & tmp_1_lpi_4_dfm_mx0c0)
      | (COMP_LOOP_COMP_LOOP_nor_5_itm & and_dcpl_245) | (COMP_LOOP_COMP_LOOP_nor_9_itm
      & and_dcpl_249) | (COMP_LOOP_COMP_LOOP_nor_13_itm & and_dcpl_254) | (COMP_LOOP_COMP_LOOP_nor_17_itm
      & and_dcpl_258) | (COMP_LOOP_COMP_LOOP_nor_21_itm & and_dcpl_262) | (COMP_LOOP_COMP_LOOP_nor_25_itm
      & and_dcpl_265) | (COMP_LOOP_COMP_LOOP_nor_29_itm & and_dcpl_269) | (COMP_LOOP_COMP_LOOP_nor_33_itm
      & and_dcpl_271) | (COMP_LOOP_COMP_LOOP_nor_37_itm & and_dcpl_273) | (COMP_LOOP_COMP_LOOP_nor_41_itm
      & and_dcpl_276) | (COMP_LOOP_COMP_LOOP_nor_45_itm & and_dcpl_278) | (COMP_LOOP_COMP_LOOP_nor_49_itm
      & and_dcpl_283) | (COMP_LOOP_COMP_LOOP_nor_53_itm & and_dcpl_285) | (COMP_LOOP_COMP_LOOP_nor_57_itm
      & and_dcpl_287) | (COMP_LOOP_COMP_LOOP_nor_61_itm & and_dcpl_289);
  assign COMP_LOOP_or_19_nl = ((operator_64_false_acc_cse_1_sva[0]) & operator_64_false_slc_operator_64_false_acc_1_60_itm
      & tmp_1_lpi_4_dfm_mx0c0) | ((operator_64_false_acc_cse_2_sva[0]) & COMP_LOOP_nor_51_itm
      & and_dcpl_245) | ((operator_64_false_acc_cse_3_sva[0]) & COMP_LOOP_nor_91_itm
      & and_dcpl_249) | ((operator_64_false_acc_cse_4_sva[0]) & COMP_LOOP_nor_131_itm
      & and_dcpl_254) | ((operator_64_false_acc_cse_5_sva[0]) & COMP_LOOP_nor_171_itm
      & and_dcpl_258) | ((operator_64_false_acc_cse_6_sva[0]) & COMP_LOOP_nor_211_itm
      & and_dcpl_262) | ((operator_64_false_acc_cse_7_sva[0]) & COMP_LOOP_nor_251_itm
      & and_dcpl_265) | ((operator_64_false_acc_cse_8_sva[0]) & COMP_LOOP_nor_291_itm
      & and_dcpl_269) | ((operator_64_false_acc_cse_9_sva[0]) & COMP_LOOP_nor_331_itm
      & and_dcpl_271) | ((operator_64_false_acc_cse_10_sva[0]) & COMP_LOOP_nor_371_itm
      & and_dcpl_273) | ((operator_64_false_acc_cse_11_sva[0]) & COMP_LOOP_nor_411_itm
      & and_dcpl_276) | ((operator_64_false_acc_cse_12_sva[0]) & COMP_LOOP_nor_451_itm
      & and_dcpl_278) | ((operator_64_false_acc_cse_13_sva[0]) & COMP_LOOP_nor_491_itm
      & and_dcpl_283) | ((operator_64_false_acc_cse_14_sva[0]) & COMP_LOOP_nor_531_itm
      & and_dcpl_285) | ((operator_64_false_acc_cse_15_sva[0]) & COMP_LOOP_nor_571_itm
      & and_dcpl_287) | ((operator_64_false_acc_cse_sva[0]) & COMP_LOOP_nor_611_itm
      & and_dcpl_289);
  assign COMP_LOOP_or_20_nl = ((operator_64_false_acc_cse_1_sva[1]) & COMP_LOOP_nor_12_itm
      & tmp_1_lpi_4_dfm_mx0c0) | ((operator_64_false_acc_cse_2_sva[1]) & COMP_LOOP_nor_52_itm
      & and_dcpl_245) | ((operator_64_false_acc_cse_3_sva[1]) & COMP_LOOP_nor_92_itm
      & and_dcpl_249) | ((operator_64_false_acc_cse_4_sva[1]) & COMP_LOOP_nor_132_itm
      & and_dcpl_254) | ((operator_64_false_acc_cse_5_sva[1]) & COMP_LOOP_nor_172_itm
      & and_dcpl_258) | ((operator_64_false_acc_cse_6_sva[1]) & COMP_LOOP_nor_212_itm
      & and_dcpl_262) | ((operator_64_false_acc_cse_7_sva[1]) & COMP_LOOP_nor_252_itm
      & and_dcpl_265) | ((operator_64_false_acc_cse_8_sva[1]) & COMP_LOOP_nor_292_itm
      & and_dcpl_269) | ((operator_64_false_acc_cse_9_sva[1]) & COMP_LOOP_nor_332_itm
      & and_dcpl_271) | ((operator_64_false_acc_cse_10_sva[1]) & COMP_LOOP_nor_372_itm
      & and_dcpl_273) | ((operator_64_false_acc_cse_11_sva[1]) & COMP_LOOP_nor_412_itm
      & and_dcpl_276) | ((operator_64_false_acc_cse_12_sva[1]) & COMP_LOOP_nor_452_itm
      & and_dcpl_278) | ((operator_64_false_acc_cse_13_sva[1]) & COMP_LOOP_nor_492_itm
      & and_dcpl_283) | ((operator_64_false_acc_cse_14_sva[1]) & COMP_LOOP_nor_532_itm
      & and_dcpl_285) | ((operator_64_false_acc_cse_15_sva[1]) & COMP_LOOP_nor_572_itm
      & and_dcpl_287) | ((operator_64_false_acc_cse_sva[1]) & COMP_LOOP_nor_612_itm
      & and_dcpl_289);
  assign COMP_LOOP_or_21_nl = (COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm
      & tmp_1_lpi_4_dfm_mx0c0) | (COMP_LOOP_COMP_LOOP_and_77_itm & and_dcpl_245)
      | (COMP_LOOP_COMP_LOOP_and_137_itm & and_dcpl_249) | (COMP_LOOP_COMP_LOOP_and_197_itm
      & and_dcpl_254) | (COMP_LOOP_COMP_LOOP_and_257_itm & and_dcpl_258) | (COMP_LOOP_COMP_LOOP_and_317_itm
      & and_dcpl_262) | (COMP_LOOP_COMP_LOOP_and_377_itm & and_dcpl_265) | (COMP_LOOP_COMP_LOOP_and_437_itm
      & and_dcpl_269) | (COMP_LOOP_COMP_LOOP_and_497_itm & and_dcpl_271) | (COMP_LOOP_COMP_LOOP_and_557_itm
      & and_dcpl_273) | (COMP_LOOP_COMP_LOOP_and_617_itm & and_dcpl_276) | (COMP_LOOP_COMP_LOOP_and_677_itm
      & and_dcpl_278) | (COMP_LOOP_COMP_LOOP_and_737_itm & and_dcpl_283) | (COMP_LOOP_COMP_LOOP_and_797_itm
      & and_dcpl_285) | (COMP_LOOP_COMP_LOOP_and_857_itm & and_dcpl_287) | (COMP_LOOP_COMP_LOOP_and_917_itm
      & and_dcpl_289);
  assign COMP_LOOP_or_22_nl = ((operator_64_false_acc_cse_1_sva[2]) & COMP_LOOP_nor_14_itm
      & tmp_1_lpi_4_dfm_mx0c0) | ((operator_64_false_acc_cse_2_sva[2]) & COMP_LOOP_nor_54_itm
      & and_dcpl_245) | ((operator_64_false_acc_cse_3_sva[2]) & COMP_LOOP_nor_94_itm
      & and_dcpl_249) | ((operator_64_false_acc_cse_4_sva[2]) & COMP_LOOP_nor_134_itm
      & and_dcpl_254) | ((operator_64_false_acc_cse_5_sva[2]) & COMP_LOOP_nor_174_itm
      & and_dcpl_258) | ((operator_64_false_acc_cse_6_sva[2]) & COMP_LOOP_nor_214_itm
      & and_dcpl_262) | ((operator_64_false_acc_cse_7_sva[2]) & COMP_LOOP_nor_254_itm
      & and_dcpl_265) | ((operator_64_false_acc_cse_8_sva[2]) & COMP_LOOP_nor_294_itm
      & and_dcpl_269) | ((operator_64_false_acc_cse_9_sva[2]) & COMP_LOOP_nor_334_itm
      & and_dcpl_271) | ((operator_64_false_acc_cse_10_sva[2]) & COMP_LOOP_nor_374_itm
      & and_dcpl_273) | ((operator_64_false_acc_cse_11_sva[2]) & COMP_LOOP_nor_414_itm
      & and_dcpl_276) | ((operator_64_false_acc_cse_12_sva[2]) & COMP_LOOP_nor_454_itm
      & and_dcpl_278) | ((operator_64_false_acc_cse_13_sva[2]) & COMP_LOOP_nor_494_itm
      & and_dcpl_283) | ((operator_64_false_acc_cse_14_sva[2]) & COMP_LOOP_nor_534_itm
      & and_dcpl_285) | ((operator_64_false_acc_cse_15_sva[2]) & COMP_LOOP_nor_574_itm
      & and_dcpl_287) | ((operator_64_false_acc_cse_sva[2]) & COMP_LOOP_nor_614_itm
      & and_dcpl_289);
  assign COMP_LOOP_or_23_nl = (COMP_LOOP_COMP_LOOP_and_19_itm & tmp_1_lpi_4_dfm_mx0c0)
      | (COMP_LOOP_COMP_LOOP_and_79_itm & and_dcpl_245) | (COMP_LOOP_COMP_LOOP_and_139_itm
      & and_dcpl_249) | (COMP_LOOP_COMP_LOOP_and_199_itm & and_dcpl_254) | (COMP_LOOP_COMP_LOOP_and_259_itm
      & and_dcpl_258) | (COMP_LOOP_COMP_LOOP_and_319_itm & and_dcpl_262) | (COMP_LOOP_COMP_LOOP_and_379_itm
      & and_dcpl_265) | (COMP_LOOP_COMP_LOOP_and_439_itm & and_dcpl_269) | (COMP_LOOP_COMP_LOOP_and_499_itm
      & and_dcpl_271) | (COMP_LOOP_COMP_LOOP_and_559_itm & and_dcpl_273) | (COMP_LOOP_COMP_LOOP_and_619_itm
      & and_dcpl_276) | (COMP_LOOP_COMP_LOOP_and_679_itm & and_dcpl_278) | (COMP_LOOP_COMP_LOOP_and_739_itm
      & and_dcpl_283) | (COMP_LOOP_COMP_LOOP_and_799_itm & and_dcpl_285) | (COMP_LOOP_COMP_LOOP_and_859_itm
      & and_dcpl_287) | (COMP_LOOP_COMP_LOOP_and_919_itm & and_dcpl_289);
  assign COMP_LOOP_or_24_nl = (COMP_LOOP_COMP_LOOP_and_20_itm & tmp_1_lpi_4_dfm_mx0c0)
      | (COMP_LOOP_COMP_LOOP_and_80_itm & and_dcpl_245) | (COMP_LOOP_COMP_LOOP_and_140_itm
      & and_dcpl_249) | (COMP_LOOP_COMP_LOOP_and_200_itm & and_dcpl_254) | (COMP_LOOP_COMP_LOOP_and_260_itm
      & and_dcpl_258) | (COMP_LOOP_COMP_LOOP_and_320_itm & and_dcpl_262) | (COMP_LOOP_COMP_LOOP_and_380_itm
      & and_dcpl_265) | (COMP_LOOP_COMP_LOOP_and_440_itm & and_dcpl_269) | (COMP_LOOP_COMP_LOOP_and_500_itm
      & and_dcpl_271) | (COMP_LOOP_COMP_LOOP_and_560_itm & and_dcpl_273) | (COMP_LOOP_COMP_LOOP_and_620_itm
      & and_dcpl_276) | (COMP_LOOP_COMP_LOOP_and_680_itm & and_dcpl_278) | (COMP_LOOP_COMP_LOOP_and_740_itm
      & and_dcpl_283) | (COMP_LOOP_COMP_LOOP_and_800_itm & and_dcpl_285) | (COMP_LOOP_COMP_LOOP_and_860_itm
      & and_dcpl_287) | (COMP_LOOP_COMP_LOOP_and_920_itm & and_dcpl_289);
  assign COMP_LOOP_or_25_nl = (COMP_LOOP_COMP_LOOP_and_21_itm & tmp_1_lpi_4_dfm_mx0c0)
      | (COMP_LOOP_COMP_LOOP_and_81_itm & and_dcpl_245) | (COMP_LOOP_COMP_LOOP_and_141_itm
      & and_dcpl_249) | (COMP_LOOP_COMP_LOOP_and_201_itm & and_dcpl_254) | (COMP_LOOP_COMP_LOOP_and_261_itm
      & and_dcpl_258) | (COMP_LOOP_COMP_LOOP_and_321_itm & and_dcpl_262) | (COMP_LOOP_COMP_LOOP_and_381_itm
      & and_dcpl_265) | (COMP_LOOP_COMP_LOOP_and_441_itm & and_dcpl_269) | (COMP_LOOP_COMP_LOOP_and_501_itm
      & and_dcpl_271) | (COMP_LOOP_COMP_LOOP_and_561_itm & and_dcpl_273) | (COMP_LOOP_COMP_LOOP_and_621_itm
      & and_dcpl_276) | (COMP_LOOP_COMP_LOOP_and_681_itm & and_dcpl_278) | (COMP_LOOP_COMP_LOOP_and_741_itm
      & and_dcpl_283) | (COMP_LOOP_COMP_LOOP_and_801_itm & and_dcpl_285) | (COMP_LOOP_COMP_LOOP_and_861_itm
      & and_dcpl_287) | (COMP_LOOP_COMP_LOOP_and_921_itm & and_dcpl_289);
  assign COMP_LOOP_or_26_nl = ((operator_64_false_acc_cse_1_sva[3]) & COMP_LOOP_nor_17_itm
      & tmp_1_lpi_4_dfm_mx0c0) | ((operator_64_false_acc_cse_2_sva[3]) & COMP_LOOP_nor_57_itm
      & and_dcpl_245) | ((operator_64_false_acc_cse_3_sva[3]) & COMP_LOOP_nor_97_itm
      & and_dcpl_249) | ((operator_64_false_acc_cse_4_sva[3]) & COMP_LOOP_nor_137_itm
      & and_dcpl_254) | ((operator_64_false_acc_cse_5_sva[3]) & COMP_LOOP_nor_177_itm
      & and_dcpl_258) | ((operator_64_false_acc_cse_6_sva[3]) & COMP_LOOP_nor_217_itm
      & and_dcpl_262) | ((operator_64_false_acc_cse_7_sva[3]) & COMP_LOOP_nor_257_itm
      & and_dcpl_265) | ((operator_64_false_acc_cse_8_sva[3]) & COMP_LOOP_nor_297_itm
      & and_dcpl_269) | ((operator_64_false_acc_cse_9_sva[3]) & COMP_LOOP_nor_337_itm
      & and_dcpl_271) | ((operator_64_false_acc_cse_10_sva[3]) & COMP_LOOP_nor_377_itm
      & and_dcpl_273) | ((operator_64_false_acc_cse_11_sva[3]) & COMP_LOOP_nor_417_itm
      & and_dcpl_276) | ((operator_64_false_acc_cse_12_sva[3]) & COMP_LOOP_nor_457_itm
      & and_dcpl_278) | ((operator_64_false_acc_cse_13_sva[3]) & COMP_LOOP_nor_497_itm
      & and_dcpl_283) | ((operator_64_false_acc_cse_14_sva[3]) & COMP_LOOP_nor_537_itm
      & and_dcpl_285) | ((operator_64_false_acc_cse_15_sva[3]) & COMP_LOOP_nor_577_itm
      & and_dcpl_287) | ((operator_64_false_acc_cse_sva[3]) & COMP_LOOP_nor_617_itm
      & and_dcpl_289);
  assign COMP_LOOP_or_27_nl = (COMP_LOOP_COMP_LOOP_and_23_itm & tmp_1_lpi_4_dfm_mx0c0)
      | (COMP_LOOP_COMP_LOOP_and_83_itm & and_dcpl_245) | (COMP_LOOP_COMP_LOOP_and_143_itm
      & and_dcpl_249) | (COMP_LOOP_COMP_LOOP_and_203_itm & and_dcpl_254) | (COMP_LOOP_COMP_LOOP_and_263_itm
      & and_dcpl_258) | (COMP_LOOP_COMP_LOOP_and_323_itm & and_dcpl_262) | (COMP_LOOP_COMP_LOOP_and_383_itm
      & and_dcpl_265) | (COMP_LOOP_COMP_LOOP_and_443_itm & and_dcpl_269) | (COMP_LOOP_COMP_LOOP_and_503_itm
      & and_dcpl_271) | (COMP_LOOP_COMP_LOOP_and_563_itm & and_dcpl_273) | (COMP_LOOP_COMP_LOOP_and_623_itm
      & and_dcpl_276) | (COMP_LOOP_COMP_LOOP_and_683_itm & and_dcpl_278) | (COMP_LOOP_COMP_LOOP_and_743_itm
      & and_dcpl_283) | (COMP_LOOP_COMP_LOOP_and_803_itm & and_dcpl_285) | (COMP_LOOP_COMP_LOOP_and_863_itm
      & and_dcpl_287) | (COMP_LOOP_COMP_LOOP_and_923_itm & and_dcpl_289);
  assign COMP_LOOP_or_28_nl = (COMP_LOOP_COMP_LOOP_and_24_itm & tmp_1_lpi_4_dfm_mx0c0)
      | (COMP_LOOP_COMP_LOOP_and_84_itm & and_dcpl_245) | (COMP_LOOP_COMP_LOOP_and_144_itm
      & and_dcpl_249) | (COMP_LOOP_COMP_LOOP_and_204_itm & and_dcpl_254) | (COMP_LOOP_COMP_LOOP_and_264_itm
      & and_dcpl_258) | (COMP_LOOP_COMP_LOOP_and_324_itm & and_dcpl_262) | (COMP_LOOP_COMP_LOOP_and_384_itm
      & and_dcpl_265) | (COMP_LOOP_COMP_LOOP_and_444_itm & and_dcpl_269) | (COMP_LOOP_COMP_LOOP_and_504_itm
      & and_dcpl_271) | (COMP_LOOP_COMP_LOOP_and_564_itm & and_dcpl_273) | (COMP_LOOP_COMP_LOOP_and_624_itm
      & and_dcpl_276) | (COMP_LOOP_COMP_LOOP_and_684_itm & and_dcpl_278) | (COMP_LOOP_COMP_LOOP_and_744_itm
      & and_dcpl_283) | (COMP_LOOP_COMP_LOOP_and_804_itm & and_dcpl_285) | (COMP_LOOP_COMP_LOOP_and_864_itm
      & and_dcpl_287) | (COMP_LOOP_COMP_LOOP_and_924_itm & and_dcpl_289);
  assign COMP_LOOP_or_29_nl = (COMP_LOOP_COMP_LOOP_and_25_itm & tmp_1_lpi_4_dfm_mx0c0)
      | (COMP_LOOP_COMP_LOOP_and_85_itm & and_dcpl_245) | (COMP_LOOP_COMP_LOOP_and_145_itm
      & and_dcpl_249) | (COMP_LOOP_COMP_LOOP_and_205_itm & and_dcpl_254) | (COMP_LOOP_COMP_LOOP_and_265_itm
      & and_dcpl_258) | (COMP_LOOP_COMP_LOOP_and_325_itm & and_dcpl_262) | (COMP_LOOP_COMP_LOOP_and_385_itm
      & and_dcpl_265) | (COMP_LOOP_COMP_LOOP_and_445_itm & and_dcpl_269) | (COMP_LOOP_COMP_LOOP_and_505_itm
      & and_dcpl_271) | (COMP_LOOP_COMP_LOOP_and_565_itm & and_dcpl_273) | (COMP_LOOP_COMP_LOOP_and_625_itm
      & and_dcpl_276) | (COMP_LOOP_COMP_LOOP_and_685_itm & and_dcpl_278) | (COMP_LOOP_COMP_LOOP_and_745_itm
      & and_dcpl_283) | (COMP_LOOP_COMP_LOOP_and_805_itm & and_dcpl_285) | (COMP_LOOP_COMP_LOOP_and_865_itm
      & and_dcpl_287) | (COMP_LOOP_COMP_LOOP_and_925_itm & and_dcpl_289);
  assign COMP_LOOP_or_30_nl = (COMP_LOOP_COMP_LOOP_and_26_itm & tmp_1_lpi_4_dfm_mx0c0)
      | (COMP_LOOP_COMP_LOOP_and_86_itm & and_dcpl_245) | (COMP_LOOP_COMP_LOOP_and_146_itm
      & and_dcpl_249) | (COMP_LOOP_COMP_LOOP_and_206_itm & and_dcpl_254) | (COMP_LOOP_COMP_LOOP_and_266_itm
      & and_dcpl_258) | (COMP_LOOP_COMP_LOOP_and_326_itm & and_dcpl_262) | (COMP_LOOP_COMP_LOOP_and_386_itm
      & and_dcpl_265) | (COMP_LOOP_COMP_LOOP_and_446_itm & and_dcpl_269) | (COMP_LOOP_COMP_LOOP_and_506_itm
      & and_dcpl_271) | (COMP_LOOP_COMP_LOOP_and_566_itm & and_dcpl_273) | (COMP_LOOP_COMP_LOOP_and_626_itm
      & and_dcpl_276) | (COMP_LOOP_COMP_LOOP_and_686_itm & and_dcpl_278) | (COMP_LOOP_COMP_LOOP_and_746_itm
      & and_dcpl_283) | (COMP_LOOP_COMP_LOOP_and_806_itm & and_dcpl_285) | (COMP_LOOP_COMP_LOOP_and_866_itm
      & and_dcpl_287) | (COMP_LOOP_COMP_LOOP_and_926_itm & and_dcpl_289);
  assign COMP_LOOP_or_31_nl = (COMP_LOOP_COMP_LOOP_and_27_itm & tmp_1_lpi_4_dfm_mx0c0)
      | (COMP_LOOP_COMP_LOOP_and_87_itm & and_dcpl_245) | (COMP_LOOP_COMP_LOOP_and_147_itm
      & and_dcpl_249) | (COMP_LOOP_COMP_LOOP_and_207_itm & and_dcpl_254) | (COMP_LOOP_COMP_LOOP_and_267_itm
      & and_dcpl_258) | (COMP_LOOP_COMP_LOOP_and_327_itm & and_dcpl_262) | (COMP_LOOP_COMP_LOOP_and_387_itm
      & and_dcpl_265) | (COMP_LOOP_COMP_LOOP_and_447_itm & and_dcpl_269) | (COMP_LOOP_COMP_LOOP_and_507_itm
      & and_dcpl_271) | (COMP_LOOP_COMP_LOOP_and_567_itm & and_dcpl_273) | (COMP_LOOP_COMP_LOOP_and_627_itm
      & and_dcpl_276) | (COMP_LOOP_COMP_LOOP_and_687_itm & and_dcpl_278) | (COMP_LOOP_COMP_LOOP_and_747_itm
      & and_dcpl_283) | (COMP_LOOP_COMP_LOOP_and_807_itm & and_dcpl_285) | (COMP_LOOP_COMP_LOOP_and_867_itm
      & and_dcpl_287) | (COMP_LOOP_COMP_LOOP_and_927_itm & and_dcpl_289);
  assign COMP_LOOP_or_32_nl = (COMP_LOOP_COMP_LOOP_and_28_itm & tmp_1_lpi_4_dfm_mx0c0)
      | (COMP_LOOP_COMP_LOOP_and_88_itm & and_dcpl_245) | (COMP_LOOP_COMP_LOOP_and_148_itm
      & and_dcpl_249) | (COMP_LOOP_COMP_LOOP_and_208_itm & and_dcpl_254) | (COMP_LOOP_COMP_LOOP_and_268_itm
      & and_dcpl_258) | (COMP_LOOP_COMP_LOOP_and_328_itm & and_dcpl_262) | (COMP_LOOP_COMP_LOOP_and_388_itm
      & and_dcpl_265) | (COMP_LOOP_COMP_LOOP_and_448_itm & and_dcpl_269) | (COMP_LOOP_COMP_LOOP_and_508_itm
      & and_dcpl_271) | (COMP_LOOP_COMP_LOOP_and_568_itm & and_dcpl_273) | (COMP_LOOP_COMP_LOOP_and_628_itm
      & and_dcpl_276) | (COMP_LOOP_COMP_LOOP_and_688_itm & and_dcpl_278) | (COMP_LOOP_COMP_LOOP_and_748_itm
      & and_dcpl_283) | (COMP_LOOP_COMP_LOOP_and_808_itm & and_dcpl_285) | (COMP_LOOP_COMP_LOOP_and_868_itm
      & and_dcpl_287) | (COMP_LOOP_COMP_LOOP_and_928_itm & and_dcpl_289);
  assign COMP_LOOP_or_33_nl = (COMP_LOOP_COMP_LOOP_and_29_itm & tmp_1_lpi_4_dfm_mx0c0)
      | (COMP_LOOP_COMP_LOOP_and_89_itm & and_dcpl_245) | (COMP_LOOP_COMP_LOOP_and_149_itm
      & and_dcpl_249) | (COMP_LOOP_COMP_LOOP_and_209_itm & and_dcpl_254) | (COMP_LOOP_COMP_LOOP_and_269_itm
      & and_dcpl_258) | (COMP_LOOP_COMP_LOOP_and_329_itm & and_dcpl_262) | (COMP_LOOP_COMP_LOOP_and_389_itm
      & and_dcpl_265) | (COMP_LOOP_COMP_LOOP_and_449_itm & and_dcpl_269) | (COMP_LOOP_COMP_LOOP_and_509_itm
      & and_dcpl_271) | (COMP_LOOP_COMP_LOOP_and_569_itm & and_dcpl_273) | (COMP_LOOP_COMP_LOOP_and_629_itm
      & and_dcpl_276) | (COMP_LOOP_COMP_LOOP_and_689_itm & and_dcpl_278) | (COMP_LOOP_COMP_LOOP_and_749_itm
      & and_dcpl_283) | (COMP_LOOP_COMP_LOOP_and_809_itm & and_dcpl_285) | (COMP_LOOP_COMP_LOOP_and_869_itm
      & and_dcpl_287) | (COMP_LOOP_COMP_LOOP_and_929_itm & and_dcpl_289);
  assign not_7089_nl = ~ not_tmp_597;
  assign nand_nl = ~((fsm_output[7]) & (fsm_output[1]) & (fsm_output[0]) & (~ (fsm_output[9]))
      & nor_tmp_1);
  assign nor_1035_nl = ~((~ (fsm_output[0])) | (fsm_output[9]) | (~ nor_tmp_1));
  assign mux_2890_nl = MUX_s_1_2_2(nor_1035_nl, nor_tmp_1, fsm_output[1]);
  assign mux_2896_nl = MUX_s_1_2_2(mux_tmp_2815, mux_tmp_2823, nor_1040_cse);
  assign mux_2889_nl = MUX_s_1_2_2(mux_tmp_2823, mux_2896_nl, fsm_output[1]);
  assign mux_2891_nl = MUX_s_1_2_2((~ mux_2890_nl), mux_2889_nl, fsm_output[7]);
  assign mux_2892_nl = MUX_s_1_2_2(nand_nl, mux_2891_nl, fsm_output[4]);
  assign mux_2895_nl = MUX_s_1_2_2(mux_tmp_2815, mux_tmp_2823, nor_1040_cse);
  assign mux_2885_nl = MUX_s_1_2_2(mux_tmp_2813, mux_tmp_2815, or_3018_cse);
  assign mux_2887_nl = MUX_s_1_2_2(mux_2895_nl, mux_2885_nl, fsm_output[1]);
  assign or_3017_nl = (fsm_output[1]) | (~((~ (fsm_output[0])) | (fsm_output[9])))
      | (fsm_output[3]) | (fsm_output[2]) | (fsm_output[6]);
  assign mux_2888_nl = MUX_s_1_2_2(mux_2887_nl, or_3017_nl, fsm_output[7]);
  assign or_3019_nl = (fsm_output[4]) | mux_2888_nl;
  assign mux_2893_nl = MUX_s_1_2_2(mux_2892_nl, or_3019_nl, fsm_output[5]);
  assign mux_2879_nl = MUX_s_1_2_2(mux_tmp_2824, (~ mux_tmp_2812), fsm_output[9]);
  assign mux_2878_nl = MUX_s_1_2_2(mux_tmp_2823, mux_tmp_2824, fsm_output[9]);
  assign mux_2880_nl = MUX_s_1_2_2(mux_2879_nl, mux_2878_nl, fsm_output[0]);
  assign mux_2881_nl = MUX_s_1_2_2(mux_2880_nl, mux_tmp_2823, fsm_output[1]);
  assign mux_2874_nl = MUX_s_1_2_2(or_307_cse, or_165_cse, or_3018_cse);
  assign mux_2875_nl = MUX_s_1_2_2(mux_2874_nl, or_307_cse, fsm_output[1]);
  assign mux_2882_nl = MUX_s_1_2_2(mux_2881_nl, mux_2875_nl, fsm_output[7]);
  assign or_3011_nl = (fsm_output[7]) | (~((~ (fsm_output[1])) | (~ (fsm_output[0]))
      | (fsm_output[9]))) | (fsm_output[3]) | (fsm_output[2]) | (fsm_output[6]);
  assign mux_2883_nl = MUX_s_1_2_2(mux_2882_nl, or_3011_nl, fsm_output[4]);
  assign or_3008_nl = (~ (fsm_output[7])) | (fsm_output[9]) | (~ nor_tmp_1);
  assign mux_2870_nl = MUX_s_1_2_2(and_711_cse, nor_tmp_1, nor_1040_cse);
  assign mux_2871_nl = MUX_s_1_2_2(nor_tmp_1, mux_2870_nl, fsm_output[1]);
  assign or_3006_nl = (fsm_output[9]) | mux_tmp_2815;
  assign or_3005_nl = (fsm_output[9]) | mux_tmp_2813;
  assign or_3004_nl = (fsm_output[9]) | mux_tmp_2812;
  assign mux_2867_nl = MUX_s_1_2_2(or_3005_nl, or_3004_nl, fsm_output[0]);
  assign mux_2869_nl = MUX_s_1_2_2(or_3006_nl, mux_2867_nl, fsm_output[1]);
  assign mux_2872_nl = MUX_s_1_2_2((~ mux_2871_nl), mux_2869_nl, fsm_output[7]);
  assign mux_2873_nl = MUX_s_1_2_2(or_3008_nl, mux_2872_nl, fsm_output[4]);
  assign mux_2884_nl = MUX_s_1_2_2(mux_2883_nl, mux_2873_nl, fsm_output[5]);
  assign COMP_LOOP_mux_291_nl = MUX_v_64_2_2(COMP_LOOP_10_modExp_dev_1_while_mul_mut,
      modExp_dev_result_sva, and_dcpl_402);
  assign or_3024_nl = (fsm_output[1]) | (fsm_output[7]) | (fsm_output[4]) | (fsm_output[5])
      | (fsm_output[3]) | (fsm_output[8]) | (~ (fsm_output[2]));
  assign or_3025_nl = (~ (fsm_output[7])) | (fsm_output[4]) | (~ (fsm_output[5]))
      | (~ (fsm_output[3])) | (fsm_output[8]) | (fsm_output[2]);
  assign mux_2900_nl = MUX_s_1_2_2(or_3025_nl, nand_tmp_150, fsm_output[1]);
  assign mux_2899_nl = MUX_s_1_2_2(or_3024_nl, mux_2900_nl, fsm_output[6]);
  assign mux_2898_nl = MUX_s_1_2_2(or_tmp_2743, mux_2899_nl, fsm_output[9]);
  assign or_3026_nl = (~ (fsm_output[7])) | (fsm_output[4]) | mux_tmp_2749;
  assign mux_2902_nl = MUX_s_1_2_2(nand_tmp_150, or_3026_nl, fsm_output[1]);
  assign nand_491_nl = ~((fsm_output[6]) & (~ mux_2902_nl));
  assign mux_2901_nl = MUX_s_1_2_2(nand_491_nl, or_tmp_2743, fsm_output[9]);
  assign mux_2897_nl = MUX_s_1_2_2(mux_2898_nl, mux_2901_nl, fsm_output[0]);
  assign COMP_LOOP_mux1h_842_nl = MUX1HOT_v_64_3_2(COMP_LOOP_1_modulo_dev_cmp_return_rsc_z,
      r_sva, modExp_dev_result_sva, {(~ mux_2897_nl) , and_dcpl_402 , (~ mux_2835_cse)});
  assign nl_z_out = COMP_LOOP_mux_291_nl * COMP_LOOP_mux1h_842_nl;
  assign z_out = nl_z_out[63:0];
  assign COMP_LOOP_mux_292_nl = MUX_v_10_2_2(({4'b0000 , (STAGE_VEC_LOOP_j_sva_9_0[9:4])}),
      STAGE_VEC_LOOP_j_sva_9_0, and_dcpl_418);
  assign COMP_LOOP_mux_293_nl = MUX_v_10_2_2(({5'b00000 , COMP_LOOP_k_9_4_sva_4_0}),
      STAGE_MAIN_LOOP_lshift_psp_1_sva, and_dcpl_418);
  assign nl_z_out_1 = conv_u2u_10_11(COMP_LOOP_mux_292_nl) + conv_u2u_10_11(COMP_LOOP_mux_293_nl);
  assign z_out_1 = nl_z_out_1[10:0];
  assign operator_64_false_operator_64_false_or_58_nl = (~(and_dcpl_427 | and_dcpl_435
      | and_dcpl_442 | and_dcpl_449 | and_dcpl_454 | and_dcpl_458 | and_dcpl_464
      | and_dcpl_468 | and_dcpl_471 | and_dcpl_474 | and_dcpl_476 | and_dcpl_478
      | and_dcpl_481 | and_dcpl_484 | and_dcpl_487 | and_dcpl_489 | and_dcpl_496
      | and_dcpl_498)) | (~ mux_2835_cse) | and_dcpl_493 | and_dcpl_495;
  assign operator_64_false_operator_64_false_mux_58_nl = MUX_s_1_2_2((z_out_3[63]),
      (STAGE_MAIN_LOOP_div_cmp_z[63]), and_dcpl_493);
  assign operator_64_false_or_130_nl = (~(operator_64_false_operator_64_false_mux_58_nl
      | and_dcpl_478 | and_dcpl_481 | and_dcpl_484 | and_dcpl_487 | and_dcpl_489))
      | and_dcpl_427 | and_dcpl_435 | and_dcpl_442 | and_dcpl_449 | and_dcpl_454
      | and_dcpl_458 | and_dcpl_464 | and_dcpl_468 | and_dcpl_471 | and_dcpl_474
      | and_dcpl_476 | and_dcpl_496 | and_dcpl_498;
  assign operator_64_false_operator_64_false_mux_59_nl = MUX_s_1_2_2((z_out_3[62]),
      (STAGE_MAIN_LOOP_div_cmp_z[62]), and_dcpl_493);
  assign operator_64_false_or_131_nl = (~(operator_64_false_operator_64_false_mux_59_nl
      | and_dcpl_478 | and_dcpl_481 | and_dcpl_484 | and_dcpl_487 | and_dcpl_489))
      | and_dcpl_427 | and_dcpl_435 | and_dcpl_442 | and_dcpl_449 | and_dcpl_454
      | and_dcpl_458 | and_dcpl_464 | and_dcpl_468 | and_dcpl_471 | and_dcpl_474
      | and_dcpl_476 | and_dcpl_496 | and_dcpl_498;
  assign operator_64_false_operator_64_false_mux_60_nl = MUX_s_1_2_2((z_out_3[61]),
      (STAGE_MAIN_LOOP_div_cmp_z[61]), and_dcpl_493);
  assign operator_64_false_or_132_nl = (~(operator_64_false_operator_64_false_mux_60_nl
      | and_dcpl_478 | and_dcpl_487 | and_dcpl_489)) | and_dcpl_427 | and_dcpl_435
      | and_dcpl_442 | and_dcpl_449 | and_dcpl_454 | and_dcpl_458 | and_dcpl_464
      | and_dcpl_468 | and_dcpl_471 | and_dcpl_474 | and_dcpl_476 | and_dcpl_481
      | and_dcpl_484 | and_dcpl_496 | and_dcpl_498;
  assign operator_64_false_operator_64_false_mux_61_nl = MUX_s_1_2_2((z_out_3[60]),
      (STAGE_MAIN_LOOP_div_cmp_z[60]), and_dcpl_493);
  assign operator_64_false_or_133_nl = (~(operator_64_false_operator_64_false_mux_61_nl
      | and_dcpl_478 | and_dcpl_487 | and_dcpl_489)) | and_dcpl_427 | and_dcpl_435
      | and_dcpl_442 | and_dcpl_449 | and_dcpl_454 | and_dcpl_458 | and_dcpl_464
      | and_dcpl_468 | and_dcpl_471 | and_dcpl_474 | and_dcpl_476 | and_dcpl_481
      | and_dcpl_484 | and_dcpl_496 | and_dcpl_498;
  assign operator_64_false_operator_64_false_mux_62_nl = MUX_s_1_2_2((z_out_3[59]),
      (STAGE_MAIN_LOOP_div_cmp_z[59]), and_dcpl_493);
  assign operator_64_false_or_134_nl = (~(operator_64_false_operator_64_false_mux_62_nl
      | and_dcpl_478 | and_dcpl_489)) | and_dcpl_427 | and_dcpl_435 | and_dcpl_442
      | and_dcpl_449 | and_dcpl_454 | and_dcpl_458 | and_dcpl_464 | and_dcpl_468
      | and_dcpl_471 | and_dcpl_474 | and_dcpl_476 | and_dcpl_481 | and_dcpl_484
      | and_dcpl_487 | and_dcpl_496 | and_dcpl_498;
  assign operator_64_false_operator_64_false_mux_63_nl = MUX_s_1_2_2((z_out_3[58]),
      (STAGE_MAIN_LOOP_div_cmp_z[58]), and_dcpl_493);
  assign operator_64_false_or_135_nl = (~(operator_64_false_operator_64_false_mux_63_nl
      | and_dcpl_478 | and_dcpl_489)) | and_dcpl_427 | and_dcpl_435 | and_dcpl_442
      | and_dcpl_449 | and_dcpl_454 | and_dcpl_458 | and_dcpl_464 | and_dcpl_468
      | and_dcpl_471 | and_dcpl_474 | and_dcpl_476 | and_dcpl_481 | and_dcpl_484
      | and_dcpl_487 | and_dcpl_496 | and_dcpl_498;
  assign operator_64_false_operator_64_false_mux_64_nl = MUX_s_1_2_2((z_out_3[57]),
      (STAGE_MAIN_LOOP_div_cmp_z[57]), and_dcpl_493);
  assign operator_64_false_or_136_nl = (~(operator_64_false_operator_64_false_mux_64_nl
      | and_dcpl_478 | and_dcpl_489)) | and_dcpl_427 | and_dcpl_435 | and_dcpl_442
      | and_dcpl_449 | and_dcpl_454 | and_dcpl_458 | and_dcpl_464 | and_dcpl_468
      | and_dcpl_471 | and_dcpl_474 | and_dcpl_476 | and_dcpl_481 | and_dcpl_484
      | and_dcpl_487 | and_dcpl_496 | and_dcpl_498;
  assign operator_64_false_operator_64_false_mux_65_nl = MUX_s_1_2_2((z_out_3[56]),
      (STAGE_MAIN_LOOP_div_cmp_z[56]), and_dcpl_493);
  assign operator_64_false_or_137_nl = (~(operator_64_false_operator_64_false_mux_65_nl
      | and_dcpl_478 | and_dcpl_489)) | and_dcpl_427 | and_dcpl_435 | and_dcpl_442
      | and_dcpl_449 | and_dcpl_454 | and_dcpl_458 | and_dcpl_464 | and_dcpl_468
      | and_dcpl_471 | and_dcpl_474 | and_dcpl_476 | and_dcpl_481 | and_dcpl_484
      | and_dcpl_487 | and_dcpl_496 | and_dcpl_498;
  assign operator_64_false_operator_64_false_mux_66_nl = MUX_s_1_2_2((z_out_3[55]),
      (STAGE_MAIN_LOOP_div_cmp_z[55]), and_dcpl_493);
  assign operator_64_false_or_138_nl = (~(operator_64_false_operator_64_false_mux_66_nl
      | and_dcpl_478 | and_dcpl_489)) | and_dcpl_427 | and_dcpl_435 | and_dcpl_442
      | and_dcpl_449 | and_dcpl_454 | and_dcpl_458 | and_dcpl_464 | and_dcpl_468
      | and_dcpl_471 | and_dcpl_474 | and_dcpl_476 | and_dcpl_481 | and_dcpl_484
      | and_dcpl_487 | and_dcpl_496 | and_dcpl_498;
  assign operator_64_false_operator_64_false_mux_67_nl = MUX_s_1_2_2((z_out_3[54]),
      (STAGE_MAIN_LOOP_div_cmp_z[54]), and_dcpl_493);
  assign operator_64_false_or_139_nl = (~(operator_64_false_operator_64_false_mux_67_nl
      | and_dcpl_478 | and_dcpl_489)) | and_dcpl_427 | and_dcpl_435 | and_dcpl_442
      | and_dcpl_449 | and_dcpl_454 | and_dcpl_458 | and_dcpl_464 | and_dcpl_468
      | and_dcpl_471 | and_dcpl_474 | and_dcpl_476 | and_dcpl_481 | and_dcpl_484
      | and_dcpl_487 | and_dcpl_496 | and_dcpl_498;
  assign operator_64_false_operator_64_false_mux_68_nl = MUX_s_1_2_2((z_out_3[53]),
      (STAGE_MAIN_LOOP_div_cmp_z[53]), and_dcpl_493);
  assign operator_64_false_or_140_nl = (~(operator_64_false_operator_64_false_mux_68_nl
      | and_dcpl_478 | and_dcpl_489)) | and_dcpl_427 | and_dcpl_435 | and_dcpl_442
      | and_dcpl_449 | and_dcpl_454 | and_dcpl_458 | and_dcpl_464 | and_dcpl_468
      | and_dcpl_471 | and_dcpl_474 | and_dcpl_476 | and_dcpl_481 | and_dcpl_484
      | and_dcpl_487 | and_dcpl_496 | and_dcpl_498;
  assign operator_64_false_operator_64_false_mux_69_nl = MUX_s_1_2_2((z_out_3[52]),
      (STAGE_MAIN_LOOP_div_cmp_z[52]), and_dcpl_493);
  assign operator_64_false_or_141_nl = (~(operator_64_false_operator_64_false_mux_69_nl
      | and_dcpl_478 | and_dcpl_489)) | and_dcpl_427 | and_dcpl_435 | and_dcpl_442
      | and_dcpl_449 | and_dcpl_454 | and_dcpl_458 | and_dcpl_464 | and_dcpl_468
      | and_dcpl_471 | and_dcpl_474 | and_dcpl_476 | and_dcpl_481 | and_dcpl_484
      | and_dcpl_487 | and_dcpl_496 | and_dcpl_498;
  assign operator_64_false_operator_64_false_mux_70_nl = MUX_s_1_2_2((z_out_3[51]),
      (STAGE_MAIN_LOOP_div_cmp_z[51]), and_dcpl_493);
  assign operator_64_false_or_142_nl = (~(operator_64_false_operator_64_false_mux_70_nl
      | and_dcpl_478 | and_dcpl_489)) | and_dcpl_427 | and_dcpl_435 | and_dcpl_442
      | and_dcpl_449 | and_dcpl_454 | and_dcpl_458 | and_dcpl_464 | and_dcpl_468
      | and_dcpl_471 | and_dcpl_474 | and_dcpl_476 | and_dcpl_481 | and_dcpl_484
      | and_dcpl_487 | and_dcpl_496 | and_dcpl_498;
  assign operator_64_false_operator_64_false_mux_71_nl = MUX_s_1_2_2((z_out_3[50]),
      (STAGE_MAIN_LOOP_div_cmp_z[50]), and_dcpl_493);
  assign operator_64_false_or_143_nl = (~(operator_64_false_operator_64_false_mux_71_nl
      | and_dcpl_478 | and_dcpl_489)) | and_dcpl_427 | and_dcpl_435 | and_dcpl_442
      | and_dcpl_449 | and_dcpl_454 | and_dcpl_458 | and_dcpl_464 | and_dcpl_468
      | and_dcpl_471 | and_dcpl_474 | and_dcpl_476 | and_dcpl_481 | and_dcpl_484
      | and_dcpl_487 | and_dcpl_496 | and_dcpl_498;
  assign operator_64_false_operator_64_false_mux_72_nl = MUX_s_1_2_2((z_out_3[49]),
      (STAGE_MAIN_LOOP_div_cmp_z[49]), and_dcpl_493);
  assign operator_64_false_or_144_nl = (~(operator_64_false_operator_64_false_mux_72_nl
      | and_dcpl_478 | and_dcpl_489)) | and_dcpl_427 | and_dcpl_435 | and_dcpl_442
      | and_dcpl_449 | and_dcpl_454 | and_dcpl_458 | and_dcpl_464 | and_dcpl_468
      | and_dcpl_471 | and_dcpl_474 | and_dcpl_476 | and_dcpl_481 | and_dcpl_484
      | and_dcpl_487 | and_dcpl_496 | and_dcpl_498;
  assign operator_64_false_operator_64_false_mux_73_nl = MUX_s_1_2_2((z_out_3[48]),
      (STAGE_MAIN_LOOP_div_cmp_z[48]), and_dcpl_493);
  assign operator_64_false_or_145_nl = (~(operator_64_false_operator_64_false_mux_73_nl
      | and_dcpl_478 | and_dcpl_489)) | and_dcpl_427 | and_dcpl_435 | and_dcpl_442
      | and_dcpl_449 | and_dcpl_454 | and_dcpl_458 | and_dcpl_464 | and_dcpl_468
      | and_dcpl_471 | and_dcpl_474 | and_dcpl_476 | and_dcpl_481 | and_dcpl_484
      | and_dcpl_487 | and_dcpl_496 | and_dcpl_498;
  assign operator_64_false_operator_64_false_mux_74_nl = MUX_s_1_2_2((z_out_3[47]),
      (STAGE_MAIN_LOOP_div_cmp_z[47]), and_dcpl_493);
  assign operator_64_false_or_146_nl = (~(operator_64_false_operator_64_false_mux_74_nl
      | and_dcpl_478 | and_dcpl_489)) | and_dcpl_427 | and_dcpl_435 | and_dcpl_442
      | and_dcpl_449 | and_dcpl_454 | and_dcpl_458 | and_dcpl_464 | and_dcpl_468
      | and_dcpl_471 | and_dcpl_474 | and_dcpl_476 | and_dcpl_481 | and_dcpl_484
      | and_dcpl_487 | and_dcpl_496 | and_dcpl_498;
  assign operator_64_false_operator_64_false_mux_75_nl = MUX_s_1_2_2((z_out_3[46]),
      (STAGE_MAIN_LOOP_div_cmp_z[46]), and_dcpl_493);
  assign operator_64_false_or_147_nl = (~(operator_64_false_operator_64_false_mux_75_nl
      | and_dcpl_478 | and_dcpl_489)) | and_dcpl_427 | and_dcpl_435 | and_dcpl_442
      | and_dcpl_449 | and_dcpl_454 | and_dcpl_458 | and_dcpl_464 | and_dcpl_468
      | and_dcpl_471 | and_dcpl_474 | and_dcpl_476 | and_dcpl_481 | and_dcpl_484
      | and_dcpl_487 | and_dcpl_496 | and_dcpl_498;
  assign operator_64_false_operator_64_false_mux_76_nl = MUX_s_1_2_2((z_out_3[45]),
      (STAGE_MAIN_LOOP_div_cmp_z[45]), and_dcpl_493);
  assign operator_64_false_or_148_nl = (~(operator_64_false_operator_64_false_mux_76_nl
      | and_dcpl_478 | and_dcpl_489)) | and_dcpl_427 | and_dcpl_435 | and_dcpl_442
      | and_dcpl_449 | and_dcpl_454 | and_dcpl_458 | and_dcpl_464 | and_dcpl_468
      | and_dcpl_471 | and_dcpl_474 | and_dcpl_476 | and_dcpl_481 | and_dcpl_484
      | and_dcpl_487 | and_dcpl_496 | and_dcpl_498;
  assign operator_64_false_operator_64_false_mux_77_nl = MUX_s_1_2_2((z_out_3[44]),
      (STAGE_MAIN_LOOP_div_cmp_z[44]), and_dcpl_493);
  assign operator_64_false_or_149_nl = (~(operator_64_false_operator_64_false_mux_77_nl
      | and_dcpl_478 | and_dcpl_489)) | and_dcpl_427 | and_dcpl_435 | and_dcpl_442
      | and_dcpl_449 | and_dcpl_454 | and_dcpl_458 | and_dcpl_464 | and_dcpl_468
      | and_dcpl_471 | and_dcpl_474 | and_dcpl_476 | and_dcpl_481 | and_dcpl_484
      | and_dcpl_487 | and_dcpl_496 | and_dcpl_498;
  assign operator_64_false_operator_64_false_mux_78_nl = MUX_s_1_2_2((z_out_3[43]),
      (STAGE_MAIN_LOOP_div_cmp_z[43]), and_dcpl_493);
  assign operator_64_false_or_150_nl = (~(operator_64_false_operator_64_false_mux_78_nl
      | and_dcpl_478 | and_dcpl_489)) | and_dcpl_427 | and_dcpl_435 | and_dcpl_442
      | and_dcpl_449 | and_dcpl_454 | and_dcpl_458 | and_dcpl_464 | and_dcpl_468
      | and_dcpl_471 | and_dcpl_474 | and_dcpl_476 | and_dcpl_481 | and_dcpl_484
      | and_dcpl_487 | and_dcpl_496 | and_dcpl_498;
  assign operator_64_false_operator_64_false_mux_79_nl = MUX_s_1_2_2((z_out_3[42]),
      (STAGE_MAIN_LOOP_div_cmp_z[42]), and_dcpl_493);
  assign operator_64_false_or_151_nl = (~(operator_64_false_operator_64_false_mux_79_nl
      | and_dcpl_478 | and_dcpl_489)) | and_dcpl_427 | and_dcpl_435 | and_dcpl_442
      | and_dcpl_449 | and_dcpl_454 | and_dcpl_458 | and_dcpl_464 | and_dcpl_468
      | and_dcpl_471 | and_dcpl_474 | and_dcpl_476 | and_dcpl_481 | and_dcpl_484
      | and_dcpl_487 | and_dcpl_496 | and_dcpl_498;
  assign operator_64_false_operator_64_false_mux_80_nl = MUX_s_1_2_2((z_out_3[41]),
      (STAGE_MAIN_LOOP_div_cmp_z[41]), and_dcpl_493);
  assign operator_64_false_or_152_nl = (~(operator_64_false_operator_64_false_mux_80_nl
      | and_dcpl_478 | and_dcpl_489)) | and_dcpl_427 | and_dcpl_435 | and_dcpl_442
      | and_dcpl_449 | and_dcpl_454 | and_dcpl_458 | and_dcpl_464 | and_dcpl_468
      | and_dcpl_471 | and_dcpl_474 | and_dcpl_476 | and_dcpl_481 | and_dcpl_484
      | and_dcpl_487 | and_dcpl_496 | and_dcpl_498;
  assign operator_64_false_operator_64_false_mux_81_nl = MUX_s_1_2_2((z_out_3[40]),
      (STAGE_MAIN_LOOP_div_cmp_z[40]), and_dcpl_493);
  assign operator_64_false_or_153_nl = (~(operator_64_false_operator_64_false_mux_81_nl
      | and_dcpl_478 | and_dcpl_489)) | and_dcpl_427 | and_dcpl_435 | and_dcpl_442
      | and_dcpl_449 | and_dcpl_454 | and_dcpl_458 | and_dcpl_464 | and_dcpl_468
      | and_dcpl_471 | and_dcpl_474 | and_dcpl_476 | and_dcpl_481 | and_dcpl_484
      | and_dcpl_487 | and_dcpl_496 | and_dcpl_498;
  assign operator_64_false_operator_64_false_mux_82_nl = MUX_s_1_2_2((z_out_3[39]),
      (STAGE_MAIN_LOOP_div_cmp_z[39]), and_dcpl_493);
  assign operator_64_false_or_154_nl = (~(operator_64_false_operator_64_false_mux_82_nl
      | and_dcpl_478 | and_dcpl_489)) | and_dcpl_427 | and_dcpl_435 | and_dcpl_442
      | and_dcpl_449 | and_dcpl_454 | and_dcpl_458 | and_dcpl_464 | and_dcpl_468
      | and_dcpl_471 | and_dcpl_474 | and_dcpl_476 | and_dcpl_481 | and_dcpl_484
      | and_dcpl_487 | and_dcpl_496 | and_dcpl_498;
  assign operator_64_false_operator_64_false_mux_83_nl = MUX_s_1_2_2((z_out_3[38]),
      (STAGE_MAIN_LOOP_div_cmp_z[38]), and_dcpl_493);
  assign operator_64_false_or_155_nl = (~(operator_64_false_operator_64_false_mux_83_nl
      | and_dcpl_478 | and_dcpl_489)) | and_dcpl_427 | and_dcpl_435 | and_dcpl_442
      | and_dcpl_449 | and_dcpl_454 | and_dcpl_458 | and_dcpl_464 | and_dcpl_468
      | and_dcpl_471 | and_dcpl_474 | and_dcpl_476 | and_dcpl_481 | and_dcpl_484
      | and_dcpl_487 | and_dcpl_496 | and_dcpl_498;
  assign operator_64_false_operator_64_false_mux_84_nl = MUX_s_1_2_2((z_out_3[37]),
      (STAGE_MAIN_LOOP_div_cmp_z[37]), and_dcpl_493);
  assign operator_64_false_or_156_nl = (~(operator_64_false_operator_64_false_mux_84_nl
      | and_dcpl_478 | and_dcpl_489)) | and_dcpl_427 | and_dcpl_435 | and_dcpl_442
      | and_dcpl_449 | and_dcpl_454 | and_dcpl_458 | and_dcpl_464 | and_dcpl_468
      | and_dcpl_471 | and_dcpl_474 | and_dcpl_476 | and_dcpl_481 | and_dcpl_484
      | and_dcpl_487 | and_dcpl_496 | and_dcpl_498;
  assign operator_64_false_operator_64_false_mux_85_nl = MUX_s_1_2_2((z_out_3[36]),
      (STAGE_MAIN_LOOP_div_cmp_z[36]), and_dcpl_493);
  assign operator_64_false_or_157_nl = (~(operator_64_false_operator_64_false_mux_85_nl
      | and_dcpl_478 | and_dcpl_489)) | and_dcpl_427 | and_dcpl_435 | and_dcpl_442
      | and_dcpl_449 | and_dcpl_454 | and_dcpl_458 | and_dcpl_464 | and_dcpl_468
      | and_dcpl_471 | and_dcpl_474 | and_dcpl_476 | and_dcpl_481 | and_dcpl_484
      | and_dcpl_487 | and_dcpl_496 | and_dcpl_498;
  assign operator_64_false_operator_64_false_mux_86_nl = MUX_s_1_2_2((z_out_3[35]),
      (STAGE_MAIN_LOOP_div_cmp_z[35]), and_dcpl_493);
  assign operator_64_false_or_158_nl = (~(operator_64_false_operator_64_false_mux_86_nl
      | and_dcpl_478 | and_dcpl_489)) | and_dcpl_427 | and_dcpl_435 | and_dcpl_442
      | and_dcpl_449 | and_dcpl_454 | and_dcpl_458 | and_dcpl_464 | and_dcpl_468
      | and_dcpl_471 | and_dcpl_474 | and_dcpl_476 | and_dcpl_481 | and_dcpl_484
      | and_dcpl_487 | and_dcpl_496 | and_dcpl_498;
  assign operator_64_false_operator_64_false_mux_87_nl = MUX_s_1_2_2((z_out_3[34]),
      (STAGE_MAIN_LOOP_div_cmp_z[34]), and_dcpl_493);
  assign operator_64_false_or_159_nl = (~(operator_64_false_operator_64_false_mux_87_nl
      | and_dcpl_478 | and_dcpl_489)) | and_dcpl_427 | and_dcpl_435 | and_dcpl_442
      | and_dcpl_449 | and_dcpl_454 | and_dcpl_458 | and_dcpl_464 | and_dcpl_468
      | and_dcpl_471 | and_dcpl_474 | and_dcpl_476 | and_dcpl_481 | and_dcpl_484
      | and_dcpl_487 | and_dcpl_496 | and_dcpl_498;
  assign operator_64_false_operator_64_false_mux_88_nl = MUX_s_1_2_2((z_out_3[33]),
      (STAGE_MAIN_LOOP_div_cmp_z[33]), and_dcpl_493);
  assign operator_64_false_or_160_nl = (~(operator_64_false_operator_64_false_mux_88_nl
      | and_dcpl_478 | and_dcpl_489)) | and_dcpl_427 | and_dcpl_435 | and_dcpl_442
      | and_dcpl_449 | and_dcpl_454 | and_dcpl_458 | and_dcpl_464 | and_dcpl_468
      | and_dcpl_471 | and_dcpl_474 | and_dcpl_476 | and_dcpl_481 | and_dcpl_484
      | and_dcpl_487 | and_dcpl_496 | and_dcpl_498;
  assign operator_64_false_operator_64_false_mux_89_nl = MUX_s_1_2_2((z_out_3[32]),
      (STAGE_MAIN_LOOP_div_cmp_z[32]), and_dcpl_493);
  assign operator_64_false_or_161_nl = (~(operator_64_false_operator_64_false_mux_89_nl
      | and_dcpl_478 | and_dcpl_489)) | and_dcpl_427 | and_dcpl_435 | and_dcpl_442
      | and_dcpl_449 | and_dcpl_454 | and_dcpl_458 | and_dcpl_464 | and_dcpl_468
      | and_dcpl_471 | and_dcpl_474 | and_dcpl_476 | and_dcpl_481 | and_dcpl_484
      | and_dcpl_487 | and_dcpl_496 | and_dcpl_498;
  assign operator_64_false_operator_64_false_mux_90_nl = MUX_s_1_2_2((z_out_3[31]),
      (STAGE_MAIN_LOOP_div_cmp_z[31]), and_dcpl_493);
  assign operator_64_false_or_162_nl = (~(operator_64_false_operator_64_false_mux_90_nl
      | and_dcpl_478 | and_dcpl_489)) | and_dcpl_427 | and_dcpl_435 | and_dcpl_442
      | and_dcpl_449 | and_dcpl_454 | and_dcpl_458 | and_dcpl_464 | and_dcpl_468
      | and_dcpl_471 | and_dcpl_474 | and_dcpl_476 | and_dcpl_481 | and_dcpl_484
      | and_dcpl_487 | and_dcpl_496 | and_dcpl_498;
  assign operator_64_false_operator_64_false_mux_91_nl = MUX_s_1_2_2((z_out_3[30]),
      (STAGE_MAIN_LOOP_div_cmp_z[30]), and_dcpl_493);
  assign operator_64_false_or_163_nl = (~(operator_64_false_operator_64_false_mux_91_nl
      | and_dcpl_478 | and_dcpl_489)) | and_dcpl_427 | and_dcpl_435 | and_dcpl_442
      | and_dcpl_449 | and_dcpl_454 | and_dcpl_458 | and_dcpl_464 | and_dcpl_468
      | and_dcpl_471 | and_dcpl_474 | and_dcpl_476 | and_dcpl_481 | and_dcpl_484
      | and_dcpl_487 | and_dcpl_496 | and_dcpl_498;
  assign operator_64_false_operator_64_false_mux_92_nl = MUX_s_1_2_2((z_out_3[29]),
      (STAGE_MAIN_LOOP_div_cmp_z[29]), and_dcpl_493);
  assign operator_64_false_or_164_nl = (~(operator_64_false_operator_64_false_mux_92_nl
      | and_dcpl_478 | and_dcpl_489)) | and_dcpl_427 | and_dcpl_435 | and_dcpl_442
      | and_dcpl_449 | and_dcpl_454 | and_dcpl_458 | and_dcpl_464 | and_dcpl_468
      | and_dcpl_471 | and_dcpl_474 | and_dcpl_476 | and_dcpl_481 | and_dcpl_484
      | and_dcpl_487 | and_dcpl_496 | and_dcpl_498;
  assign operator_64_false_operator_64_false_mux_93_nl = MUX_s_1_2_2((z_out_3[28]),
      (STAGE_MAIN_LOOP_div_cmp_z[28]), and_dcpl_493);
  assign operator_64_false_or_165_nl = (~(operator_64_false_operator_64_false_mux_93_nl
      | and_dcpl_478 | and_dcpl_489)) | and_dcpl_427 | and_dcpl_435 | and_dcpl_442
      | and_dcpl_449 | and_dcpl_454 | and_dcpl_458 | and_dcpl_464 | and_dcpl_468
      | and_dcpl_471 | and_dcpl_474 | and_dcpl_476 | and_dcpl_481 | and_dcpl_484
      | and_dcpl_487 | and_dcpl_496 | and_dcpl_498;
  assign operator_64_false_operator_64_false_mux_94_nl = MUX_s_1_2_2((z_out_3[27]),
      (STAGE_MAIN_LOOP_div_cmp_z[27]), and_dcpl_493);
  assign operator_64_false_or_166_nl = (~(operator_64_false_operator_64_false_mux_94_nl
      | and_dcpl_478 | and_dcpl_489)) | and_dcpl_427 | and_dcpl_435 | and_dcpl_442
      | and_dcpl_449 | and_dcpl_454 | and_dcpl_458 | and_dcpl_464 | and_dcpl_468
      | and_dcpl_471 | and_dcpl_474 | and_dcpl_476 | and_dcpl_481 | and_dcpl_484
      | and_dcpl_487 | and_dcpl_496 | and_dcpl_498;
  assign operator_64_false_operator_64_false_mux_95_nl = MUX_s_1_2_2((z_out_3[26]),
      (STAGE_MAIN_LOOP_div_cmp_z[26]), and_dcpl_493);
  assign operator_64_false_or_167_nl = (~(operator_64_false_operator_64_false_mux_95_nl
      | and_dcpl_478 | and_dcpl_489)) | and_dcpl_427 | and_dcpl_435 | and_dcpl_442
      | and_dcpl_449 | and_dcpl_454 | and_dcpl_458 | and_dcpl_464 | and_dcpl_468
      | and_dcpl_471 | and_dcpl_474 | and_dcpl_476 | and_dcpl_481 | and_dcpl_484
      | and_dcpl_487 | and_dcpl_496 | and_dcpl_498;
  assign operator_64_false_operator_64_false_mux_96_nl = MUX_s_1_2_2((z_out_3[25]),
      (STAGE_MAIN_LOOP_div_cmp_z[25]), and_dcpl_493);
  assign operator_64_false_or_168_nl = (~(operator_64_false_operator_64_false_mux_96_nl
      | and_dcpl_478 | and_dcpl_489)) | and_dcpl_427 | and_dcpl_435 | and_dcpl_442
      | and_dcpl_449 | and_dcpl_454 | and_dcpl_458 | and_dcpl_464 | and_dcpl_468
      | and_dcpl_471 | and_dcpl_474 | and_dcpl_476 | and_dcpl_481 | and_dcpl_484
      | and_dcpl_487 | and_dcpl_496 | and_dcpl_498;
  assign operator_64_false_operator_64_false_mux_97_nl = MUX_s_1_2_2((z_out_3[24]),
      (STAGE_MAIN_LOOP_div_cmp_z[24]), and_dcpl_493);
  assign operator_64_false_or_169_nl = (~(operator_64_false_operator_64_false_mux_97_nl
      | and_dcpl_478 | and_dcpl_489)) | and_dcpl_427 | and_dcpl_435 | and_dcpl_442
      | and_dcpl_449 | and_dcpl_454 | and_dcpl_458 | and_dcpl_464 | and_dcpl_468
      | and_dcpl_471 | and_dcpl_474 | and_dcpl_476 | and_dcpl_481 | and_dcpl_484
      | and_dcpl_487 | and_dcpl_496 | and_dcpl_498;
  assign operator_64_false_operator_64_false_mux_98_nl = MUX_s_1_2_2((z_out_3[23]),
      (STAGE_MAIN_LOOP_div_cmp_z[23]), and_dcpl_493);
  assign operator_64_false_or_170_nl = (~(operator_64_false_operator_64_false_mux_98_nl
      | and_dcpl_478 | and_dcpl_489)) | and_dcpl_427 | and_dcpl_435 | and_dcpl_442
      | and_dcpl_449 | and_dcpl_454 | and_dcpl_458 | and_dcpl_464 | and_dcpl_468
      | and_dcpl_471 | and_dcpl_474 | and_dcpl_476 | and_dcpl_481 | and_dcpl_484
      | and_dcpl_487 | and_dcpl_496 | and_dcpl_498;
  assign operator_64_false_operator_64_false_mux_99_nl = MUX_s_1_2_2((z_out_3[22]),
      (STAGE_MAIN_LOOP_div_cmp_z[22]), and_dcpl_493);
  assign operator_64_false_or_171_nl = (~(operator_64_false_operator_64_false_mux_99_nl
      | and_dcpl_478 | and_dcpl_489)) | and_dcpl_427 | and_dcpl_435 | and_dcpl_442
      | and_dcpl_449 | and_dcpl_454 | and_dcpl_458 | and_dcpl_464 | and_dcpl_468
      | and_dcpl_471 | and_dcpl_474 | and_dcpl_476 | and_dcpl_481 | and_dcpl_484
      | and_dcpl_487 | and_dcpl_496 | and_dcpl_498;
  assign operator_64_false_operator_64_false_mux_100_nl = MUX_s_1_2_2((z_out_3[21]),
      (STAGE_MAIN_LOOP_div_cmp_z[21]), and_dcpl_493);
  assign operator_64_false_or_172_nl = (~(operator_64_false_operator_64_false_mux_100_nl
      | and_dcpl_478 | and_dcpl_489)) | and_dcpl_427 | and_dcpl_435 | and_dcpl_442
      | and_dcpl_449 | and_dcpl_454 | and_dcpl_458 | and_dcpl_464 | and_dcpl_468
      | and_dcpl_471 | and_dcpl_474 | and_dcpl_476 | and_dcpl_481 | and_dcpl_484
      | and_dcpl_487 | and_dcpl_496 | and_dcpl_498;
  assign operator_64_false_operator_64_false_mux_101_nl = MUX_s_1_2_2((z_out_3[20]),
      (STAGE_MAIN_LOOP_div_cmp_z[20]), and_dcpl_493);
  assign operator_64_false_or_173_nl = (~(operator_64_false_operator_64_false_mux_101_nl
      | and_dcpl_478 | and_dcpl_489)) | and_dcpl_427 | and_dcpl_435 | and_dcpl_442
      | and_dcpl_449 | and_dcpl_454 | and_dcpl_458 | and_dcpl_464 | and_dcpl_468
      | and_dcpl_471 | and_dcpl_474 | and_dcpl_476 | and_dcpl_481 | and_dcpl_484
      | and_dcpl_487 | and_dcpl_496 | and_dcpl_498;
  assign operator_64_false_operator_64_false_mux_102_nl = MUX_s_1_2_2((z_out_3[19]),
      (STAGE_MAIN_LOOP_div_cmp_z[19]), and_dcpl_493);
  assign operator_64_false_or_174_nl = (~(operator_64_false_operator_64_false_mux_102_nl
      | and_dcpl_478 | and_dcpl_489)) | and_dcpl_427 | and_dcpl_435 | and_dcpl_442
      | and_dcpl_449 | and_dcpl_454 | and_dcpl_458 | and_dcpl_464 | and_dcpl_468
      | and_dcpl_471 | and_dcpl_474 | and_dcpl_476 | and_dcpl_481 | and_dcpl_484
      | and_dcpl_487 | and_dcpl_496 | and_dcpl_498;
  assign operator_64_false_operator_64_false_mux_103_nl = MUX_s_1_2_2((z_out_3[18]),
      (STAGE_MAIN_LOOP_div_cmp_z[18]), and_dcpl_493);
  assign operator_64_false_or_175_nl = (~(operator_64_false_operator_64_false_mux_103_nl
      | and_dcpl_478 | and_dcpl_489)) | and_dcpl_427 | and_dcpl_435 | and_dcpl_442
      | and_dcpl_449 | and_dcpl_454 | and_dcpl_458 | and_dcpl_464 | and_dcpl_468
      | and_dcpl_471 | and_dcpl_474 | and_dcpl_476 | and_dcpl_481 | and_dcpl_484
      | and_dcpl_487 | and_dcpl_496 | and_dcpl_498;
  assign operator_64_false_operator_64_false_mux_104_nl = MUX_s_1_2_2((z_out_3[17]),
      (STAGE_MAIN_LOOP_div_cmp_z[17]), and_dcpl_493);
  assign operator_64_false_or_176_nl = (~(operator_64_false_operator_64_false_mux_104_nl
      | and_dcpl_478 | and_dcpl_489)) | and_dcpl_427 | and_dcpl_435 | and_dcpl_442
      | and_dcpl_449 | and_dcpl_454 | and_dcpl_458 | and_dcpl_464 | and_dcpl_468
      | and_dcpl_471 | and_dcpl_474 | and_dcpl_476 | and_dcpl_481 | and_dcpl_484
      | and_dcpl_487 | and_dcpl_496 | and_dcpl_498;
  assign operator_64_false_operator_64_false_mux_105_nl = MUX_s_1_2_2((z_out_3[16]),
      (STAGE_MAIN_LOOP_div_cmp_z[16]), and_dcpl_493);
  assign operator_64_false_or_177_nl = (~(operator_64_false_operator_64_false_mux_105_nl
      | and_dcpl_478 | and_dcpl_489)) | and_dcpl_427 | and_dcpl_435 | and_dcpl_442
      | and_dcpl_449 | and_dcpl_454 | and_dcpl_458 | and_dcpl_464 | and_dcpl_468
      | and_dcpl_471 | and_dcpl_474 | and_dcpl_476 | and_dcpl_481 | and_dcpl_484
      | and_dcpl_487 | and_dcpl_496 | and_dcpl_498;
  assign operator_64_false_operator_64_false_mux_106_nl = MUX_s_1_2_2((z_out_3[15]),
      (STAGE_MAIN_LOOP_div_cmp_z[15]), and_dcpl_493);
  assign operator_64_false_or_178_nl = (~(operator_64_false_operator_64_false_mux_106_nl
      | and_dcpl_478 | and_dcpl_489)) | and_dcpl_427 | and_dcpl_435 | and_dcpl_442
      | and_dcpl_449 | and_dcpl_454 | and_dcpl_458 | and_dcpl_464 | and_dcpl_468
      | and_dcpl_471 | and_dcpl_474 | and_dcpl_476 | and_dcpl_481 | and_dcpl_484
      | and_dcpl_487 | and_dcpl_496 | and_dcpl_498;
  assign operator_64_false_operator_64_false_mux_107_nl = MUX_s_1_2_2((z_out_3[14]),
      (STAGE_MAIN_LOOP_div_cmp_z[14]), and_dcpl_493);
  assign operator_64_false_or_179_nl = (~(operator_64_false_operator_64_false_mux_107_nl
      | and_dcpl_478 | and_dcpl_489)) | and_dcpl_427 | and_dcpl_435 | and_dcpl_442
      | and_dcpl_449 | and_dcpl_454 | and_dcpl_458 | and_dcpl_464 | and_dcpl_468
      | and_dcpl_471 | and_dcpl_474 | and_dcpl_476 | and_dcpl_481 | and_dcpl_484
      | and_dcpl_487 | and_dcpl_496 | and_dcpl_498;
  assign operator_64_false_operator_64_false_mux_108_nl = MUX_s_1_2_2((z_out_3[13]),
      (STAGE_MAIN_LOOP_div_cmp_z[13]), and_dcpl_493);
  assign operator_64_false_or_180_nl = (~(operator_64_false_operator_64_false_mux_108_nl
      | and_dcpl_478 | and_dcpl_489)) | and_dcpl_427 | and_dcpl_435 | and_dcpl_442
      | and_dcpl_449 | and_dcpl_454 | and_dcpl_458 | and_dcpl_464 | and_dcpl_468
      | and_dcpl_471 | and_dcpl_474 | and_dcpl_476 | and_dcpl_481 | and_dcpl_484
      | and_dcpl_487 | and_dcpl_496 | and_dcpl_498;
  assign operator_64_false_operator_64_false_mux_109_nl = MUX_s_1_2_2((z_out_3[12]),
      (STAGE_MAIN_LOOP_div_cmp_z[12]), and_dcpl_493);
  assign operator_64_false_or_181_nl = (~(operator_64_false_operator_64_false_mux_109_nl
      | and_dcpl_478 | and_dcpl_489)) | and_dcpl_427 | and_dcpl_435 | and_dcpl_442
      | and_dcpl_449 | and_dcpl_454 | and_dcpl_458 | and_dcpl_464 | and_dcpl_468
      | and_dcpl_471 | and_dcpl_474 | and_dcpl_476 | and_dcpl_481 | and_dcpl_484
      | and_dcpl_487 | and_dcpl_496 | and_dcpl_498;
  assign operator_64_false_operator_64_false_mux_110_nl = MUX_s_1_2_2((z_out_3[11]),
      (STAGE_MAIN_LOOP_div_cmp_z[11]), and_dcpl_493);
  assign operator_64_false_or_182_nl = (~(operator_64_false_operator_64_false_mux_110_nl
      | and_dcpl_478 | and_dcpl_489)) | and_dcpl_427 | and_dcpl_435 | and_dcpl_442
      | and_dcpl_449 | and_dcpl_454 | and_dcpl_458 | and_dcpl_464 | and_dcpl_468
      | and_dcpl_471 | and_dcpl_474 | and_dcpl_476 | and_dcpl_481 | and_dcpl_484
      | and_dcpl_487 | and_dcpl_496 | and_dcpl_498;
  assign operator_64_false_operator_64_false_mux_111_nl = MUX_s_1_2_2((z_out_3[10]),
      (STAGE_MAIN_LOOP_div_cmp_z[10]), and_dcpl_493);
  assign operator_64_false_or_183_nl = (~(operator_64_false_operator_64_false_mux_111_nl
      | and_dcpl_478 | and_dcpl_489)) | and_dcpl_427 | and_dcpl_435 | and_dcpl_442
      | and_dcpl_449 | and_dcpl_454 | and_dcpl_458 | and_dcpl_464 | and_dcpl_468
      | and_dcpl_471 | and_dcpl_474 | and_dcpl_476 | and_dcpl_481 | and_dcpl_484
      | and_dcpl_487 | and_dcpl_496 | and_dcpl_498;
  assign operator_64_false_operator_64_false_mux_112_nl = MUX_s_1_2_2((z_out_3[9]),
      (STAGE_MAIN_LOOP_div_cmp_z[9]), and_dcpl_493);
  assign operator_64_false_or_184_nl = (~(operator_64_false_operator_64_false_mux_112_nl
      | and_dcpl_478 | and_dcpl_489)) | and_dcpl_427 | and_dcpl_435 | and_dcpl_442
      | and_dcpl_449 | and_dcpl_454 | and_dcpl_458 | and_dcpl_464 | and_dcpl_468
      | and_dcpl_471 | and_dcpl_474 | and_dcpl_476 | and_dcpl_481 | and_dcpl_484
      | and_dcpl_487 | and_dcpl_496 | and_dcpl_498;
  assign operator_64_false_mux1h_62_nl = MUX1HOT_v_2_4_2((STAGE_MAIN_LOOP_lshift_psp_1_sva[9:8]),
      ({1'b1 , (~ (STAGE_VEC_LOOP_j_sva_9_0[9]))}), (z_out_3[8:7]), (STAGE_MAIN_LOOP_div_cmp_z[8:7]),
      {operator_64_false_or_120_itm , and_dcpl_478 , operator_64_false_or_121_cse
      , and_dcpl_493});
  assign operator_64_false_operator_64_false_nor_111_nl = ~(MUX_v_2_2_2(operator_64_false_mux1h_62_nl,
      2'b11, and_dcpl_489));
  assign operator_64_false_or_186_nl = and_dcpl_481 | and_dcpl_484 | and_dcpl_487;
  assign operator_64_false_or_185_nl = MUX_v_2_2_2(operator_64_false_operator_64_false_nor_111_nl,
      2'b11, operator_64_false_or_186_nl);
  assign operator_64_false_or_187_nl = and_dcpl_481 | and_dcpl_484;
  assign operator_64_false_mux1h_63_nl = MUX1HOT_v_7_7_2((~ (STAGE_MAIN_LOOP_lshift_psp_1_sva[7:1])),
      (STAGE_VEC_LOOP_j_sva_9_0[8:2]), (~ (STAGE_MAIN_LOOP_lshift_psp_1_sva[9:3])),
      ({2'b11 , (~ (STAGE_MAIN_LOOP_lshift_psp_1_sva[9:5]))}), (~ (z_out_3[6:0])),
      ({3'b000 , STAGE_MAIN_LOOP_acc_1_psp_sva}), (~ (STAGE_MAIN_LOOP_div_cmp_z[6:0])),
      {operator_64_false_or_120_itm , and_dcpl_478 , operator_64_false_or_187_nl
      , and_dcpl_487 , operator_64_false_or_121_cse , and_dcpl_489 , and_dcpl_493});
  assign operator_64_false_or_188_nl = (~(and_dcpl_478 | (~ mux_2835_cse) | and_dcpl_489
      | and_dcpl_493 | and_dcpl_495 | and_dcpl_496)) | and_dcpl_427 | and_dcpl_435
      | and_dcpl_442 | and_dcpl_449 | and_dcpl_454 | and_dcpl_458 | and_dcpl_464
      | and_dcpl_468 | and_dcpl_471 | and_dcpl_474 | and_dcpl_476 | and_dcpl_481
      | and_dcpl_484 | and_dcpl_487 | and_dcpl_498;
  assign operator_64_false_operator_64_false_or_59_nl = ((COMP_LOOP_slc_acc_3_12_1_slc[5])
      & (~(and_dcpl_427 | and_dcpl_435 | and_dcpl_442 | and_dcpl_449 | and_dcpl_454
      | and_dcpl_458 | and_dcpl_464 | and_dcpl_468 | and_dcpl_471 | and_dcpl_474
      | and_dcpl_476 | and_dcpl_478 | and_dcpl_481 | and_dcpl_484 | and_dcpl_487
      | (~ mux_2835_cse) | and_dcpl_493 | and_dcpl_495 | and_dcpl_496))) | and_dcpl_489;
  assign operator_64_false_operator_64_false_mux_113_nl = MUX_v_2_2_2((COMP_LOOP_k_9_4_sva_4_0[4:3]),
      (COMP_LOOP_slc_acc_3_12_1_slc[4:3]), and_dcpl_498);
  assign operator_64_false_nor_121_nl = ~(and_dcpl_478 | and_dcpl_481 | and_dcpl_484
      | and_dcpl_487 | (~ mux_2835_cse) | and_dcpl_493 | and_dcpl_495 | and_dcpl_496);
  assign operator_64_false_and_65_nl = MUX_v_2_2_2(2'b00, operator_64_false_operator_64_false_mux_113_nl,
      operator_64_false_nor_121_nl);
  assign operator_64_false_or_189_nl = MUX_v_2_2_2(operator_64_false_and_65_nl, 2'b11,
      and_dcpl_489);
  assign operator_64_false_or_191_nl = and_dcpl_427 | and_dcpl_435 | and_dcpl_442
      | and_dcpl_449 | and_dcpl_454 | and_dcpl_458 | and_dcpl_464 | and_dcpl_468
      | and_dcpl_471 | and_dcpl_474 | and_dcpl_476;
  assign operator_64_false_or_192_nl = and_dcpl_478 | and_dcpl_481 | and_dcpl_484;
  assign operator_64_false_mux1h_64_nl = MUX1HOT_v_3_4_2((COMP_LOOP_k_9_4_sva_4_0[2:0]),
      (COMP_LOOP_k_9_4_sva_4_0[4:2]), ({2'b00 , (COMP_LOOP_k_9_4_sva_4_0[4])}), (COMP_LOOP_slc_acc_3_12_1_slc[2:0]),
      {operator_64_false_or_191_nl , operator_64_false_or_192_nl , and_dcpl_487 ,
      and_dcpl_498});
  assign operator_64_false_nor_122_nl = ~((~ mux_2835_cse) | and_dcpl_493 | and_dcpl_495
      | and_dcpl_496);
  assign operator_64_false_and_66_nl = MUX_v_3_2_2(3'b000, operator_64_false_mux1h_64_nl,
      operator_64_false_nor_122_nl);
  assign operator_64_false_or_190_nl = MUX_v_3_2_2(operator_64_false_and_66_nl, 3'b111,
      and_dcpl_489);
  assign operator_64_false_operator_64_false_mux_114_nl = MUX_s_1_2_2((COMP_LOOP_k_9_4_sva_4_0[1]),
      (COMP_LOOP_k_9_4_sva_4_0[3]), and_dcpl_487);
  assign operator_64_false_or_193_nl = (operator_64_false_operator_64_false_mux_114_nl
      & (~(and_dcpl_427 | and_dcpl_435 | and_dcpl_442 | and_dcpl_449 | and_dcpl_454
      | (~ mux_2835_cse) | and_dcpl_493 | and_dcpl_495 | and_dcpl_496 | and_dcpl_498)))
      | and_dcpl_458 | and_dcpl_464 | and_dcpl_468 | and_dcpl_471 | and_dcpl_474
      | and_dcpl_476 | and_dcpl_489;
  assign operator_64_false_operator_64_false_mux_115_nl = MUX_s_1_2_2((COMP_LOOP_k_9_4_sva_4_0[0]),
      (COMP_LOOP_k_9_4_sva_4_0[2]), and_dcpl_487);
  assign operator_64_false_or_194_nl = (operator_64_false_operator_64_false_mux_115_nl
      & (~(and_dcpl_427 | and_dcpl_435 | and_dcpl_458 | and_dcpl_464 | and_dcpl_468
      | (~ mux_2835_cse) | and_dcpl_493 | and_dcpl_495 | and_dcpl_496 | and_dcpl_498)))
      | and_dcpl_442 | and_dcpl_449 | and_dcpl_454 | and_dcpl_471 | and_dcpl_474
      | and_dcpl_476 | and_dcpl_489;
  assign operator_64_false_operator_64_false_or_60_nl = ((COMP_LOOP_k_9_4_sva_4_0[1])
      & (~(and_dcpl_427 | and_dcpl_442 | and_dcpl_449 | and_dcpl_458 | and_dcpl_464
      | and_dcpl_471 | and_dcpl_474 | and_dcpl_481 | (~ mux_2835_cse) | and_dcpl_493
      | and_dcpl_495 | and_dcpl_496 | and_dcpl_498))) | and_dcpl_435 | and_dcpl_454
      | and_dcpl_468 | and_dcpl_476 | and_dcpl_478 | and_dcpl_484 | and_dcpl_489;
  assign operator_64_false_operator_64_false_or_61_nl = ((COMP_LOOP_k_9_4_sva_4_0[0])
      & (~(and_dcpl_435 | and_dcpl_442 | and_dcpl_454 | and_dcpl_458 | and_dcpl_468
      | and_dcpl_471 | and_dcpl_476 | and_dcpl_481 | and_dcpl_484 | and_dcpl_498)))
      | and_dcpl_427 | and_dcpl_449 | and_dcpl_464 | and_dcpl_474 | and_dcpl_478
      | (~ mux_2835_cse) | and_dcpl_489 | and_dcpl_493 | and_dcpl_495 | and_dcpl_496;
  assign nl_acc_1_nl = ({operator_64_false_operator_64_false_or_58_nl , operator_64_false_or_130_nl
      , operator_64_false_or_131_nl , operator_64_false_or_132_nl , operator_64_false_or_133_nl
      , operator_64_false_or_134_nl , operator_64_false_or_135_nl , operator_64_false_or_136_nl
      , operator_64_false_or_137_nl , operator_64_false_or_138_nl , operator_64_false_or_139_nl
      , operator_64_false_or_140_nl , operator_64_false_or_141_nl , operator_64_false_or_142_nl
      , operator_64_false_or_143_nl , operator_64_false_or_144_nl , operator_64_false_or_145_nl
      , operator_64_false_or_146_nl , operator_64_false_or_147_nl , operator_64_false_or_148_nl
      , operator_64_false_or_149_nl , operator_64_false_or_150_nl , operator_64_false_or_151_nl
      , operator_64_false_or_152_nl , operator_64_false_or_153_nl , operator_64_false_or_154_nl
      , operator_64_false_or_155_nl , operator_64_false_or_156_nl , operator_64_false_or_157_nl
      , operator_64_false_or_158_nl , operator_64_false_or_159_nl , operator_64_false_or_160_nl
      , operator_64_false_or_161_nl , operator_64_false_or_162_nl , operator_64_false_or_163_nl
      , operator_64_false_or_164_nl , operator_64_false_or_165_nl , operator_64_false_or_166_nl
      , operator_64_false_or_167_nl , operator_64_false_or_168_nl , operator_64_false_or_169_nl
      , operator_64_false_or_170_nl , operator_64_false_or_171_nl , operator_64_false_or_172_nl
      , operator_64_false_or_173_nl , operator_64_false_or_174_nl , operator_64_false_or_175_nl
      , operator_64_false_or_176_nl , operator_64_false_or_177_nl , operator_64_false_or_178_nl
      , operator_64_false_or_179_nl , operator_64_false_or_180_nl , operator_64_false_or_181_nl
      , operator_64_false_or_182_nl , operator_64_false_or_183_nl , operator_64_false_or_184_nl
      , operator_64_false_or_185_nl , operator_64_false_mux1h_63_nl , operator_64_false_or_188_nl})
      + conv_s2u_65_66({operator_64_false_operator_64_false_or_1_cse , operator_64_false_operator_64_false_or_1_cse
      , operator_64_false_operator_64_false_or_1_cse , operator_64_false_operator_64_false_or_1_cse
      , operator_64_false_operator_64_false_or_1_cse , operator_64_false_operator_64_false_or_1_cse
      , operator_64_false_operator_64_false_or_1_cse , operator_64_false_operator_64_false_or_1_cse
      , operator_64_false_operator_64_false_or_1_cse , operator_64_false_operator_64_false_or_1_cse
      , operator_64_false_operator_64_false_or_1_cse , operator_64_false_operator_64_false_or_1_cse
      , operator_64_false_operator_64_false_or_1_cse , operator_64_false_operator_64_false_or_1_cse
      , operator_64_false_operator_64_false_or_1_cse , operator_64_false_operator_64_false_or_1_cse
      , operator_64_false_operator_64_false_or_1_cse , operator_64_false_operator_64_false_or_1_cse
      , operator_64_false_operator_64_false_or_1_cse , operator_64_false_operator_64_false_or_1_cse
      , operator_64_false_operator_64_false_or_1_cse , operator_64_false_operator_64_false_or_1_cse
      , operator_64_false_operator_64_false_or_1_cse , operator_64_false_operator_64_false_or_1_cse
      , operator_64_false_operator_64_false_or_1_cse , operator_64_false_operator_64_false_or_1_cse
      , operator_64_false_operator_64_false_or_1_cse , operator_64_false_operator_64_false_or_1_cse
      , operator_64_false_operator_64_false_or_1_cse , operator_64_false_operator_64_false_or_1_cse
      , operator_64_false_operator_64_false_or_1_cse , operator_64_false_operator_64_false_or_1_cse
      , operator_64_false_operator_64_false_or_1_cse , operator_64_false_operator_64_false_or_1_cse
      , operator_64_false_operator_64_false_or_1_cse , operator_64_false_operator_64_false_or_1_cse
      , operator_64_false_operator_64_false_or_1_cse , operator_64_false_operator_64_false_or_1_cse
      , operator_64_false_operator_64_false_or_1_cse , operator_64_false_operator_64_false_or_1_cse
      , operator_64_false_operator_64_false_or_1_cse , operator_64_false_operator_64_false_or_1_cse
      , operator_64_false_operator_64_false_or_1_cse , operator_64_false_operator_64_false_or_1_cse
      , operator_64_false_operator_64_false_or_1_cse , operator_64_false_operator_64_false_or_1_cse
      , operator_64_false_operator_64_false_or_1_cse , operator_64_false_operator_64_false_or_1_cse
      , operator_64_false_operator_64_false_or_1_cse , operator_64_false_operator_64_false_or_1_cse
      , operator_64_false_operator_64_false_or_1_cse , operator_64_false_operator_64_false_or_1_cse
      , operator_64_false_operator_64_false_or_1_cse , operator_64_false_operator_64_false_or_1_cse
      , operator_64_false_operator_64_false_or_59_nl , operator_64_false_or_189_nl
      , operator_64_false_or_190_nl , operator_64_false_or_193_nl , operator_64_false_or_194_nl
      , operator_64_false_operator_64_false_or_60_nl , operator_64_false_operator_64_false_or_61_nl
      , 1'b1});
  assign acc_1_nl = nl_acc_1_nl[65:0];
  assign z_out_2 = readslicef_66_65_1(acc_1_nl);
  assign operator_64_false_or_7_nl = and_dcpl_511 | (~ mux_2863_itm) | and_925_cse
      | and_dcpl_525 | and_936_cse | and_940_cse | and_945_cse | and_950_cse | and_953_cse
      | and_957_cse | and_960_cse | and_964_cse | and_966_cse | and_970_cse | and_973_cse
      | and_975_cse | and_978_cse;
  assign operator_64_false_mux1h_3_nl = MUX1HOT_v_64_4_2(p_sva, tmp_10_lpi_4_dfm,
      ({modExp_dev_exp_1_sva_63_9 , modExp_dev_exp_1_sva_8_4 , (COMP_LOOP_acc_psp_sva[3:0])}),
      z_out_5, {and_dcpl_507 , operator_64_false_or_7_nl , (~ mux_2835_cse) , and_920_cse});
  assign operator_64_false_operator_64_false_nand_1_nl = ~((and_dcpl_507 | and_dcpl_511
      | (~ mux_2835_cse) | and_920_cse | and_925_cse | and_dcpl_525 | and_936_cse
      | and_940_cse | and_945_cse | and_950_cse | and_953_cse | and_957_cse | and_960_cse
      | and_964_cse | and_966_cse | and_970_cse | and_973_cse | and_975_cse | and_978_cse)
      & mux_2863_itm);
  assign operator_64_false_or_10_nl = and_925_cse | and_dcpl_525 | and_936_cse |
      and_940_cse | and_945_cse | and_950_cse | and_953_cse | and_957_cse | and_960_cse
      | and_964_cse | and_966_cse | and_970_cse | and_973_cse | and_975_cse | and_978_cse;
  assign operator_64_false_mux1h_4_nl = MUX1HOT_v_64_3_2(tmp_1_lpi_4_dfm, (~ tmp_1_lpi_4_dfm),
      z_out_5, {and_920_cse , (~ mux_2863_itm) , operator_64_false_or_10_nl});
  assign operator_64_false_or_11_nl = and_dcpl_507 | and_dcpl_511 | (~ mux_2835_cse);
  assign operator_64_false_or_9_nl = MUX_v_64_2_2(operator_64_false_mux1h_4_nl, 64'b1111111111111111111111111111111111111111111111111111111111111111,
      operator_64_false_or_11_nl);
  assign nl_acc_2_nl = ({operator_64_false_mux1h_3_nl , operator_64_false_operator_64_false_nand_1_nl})
      + ({operator_64_false_or_9_nl , 1'b1});
  assign acc_2_nl = nl_acc_2_nl[64:0];
  assign z_out_3 = readslicef_65_64_1(acc_2_nl);
  assign COMP_LOOP_COMP_LOOP_or_3_nl = (~(and_dcpl_582 | and_dcpl_599)) | and_dcpl_589
      | and_dcpl_593;
  assign not_7303_nl = ~ and_dcpl_599;
  assign COMP_LOOP_and_451_nl = MUX_v_4_2_2(4'b0000, (STAGE_VEC_LOOP_j_sva_9_0[9:6]),
      not_7303_nl);
  assign COMP_LOOP_or_41_nl = and_dcpl_589 | and_dcpl_593;
  assign COMP_LOOP_COMP_LOOP_or_4_nl = MUX_v_4_2_2(COMP_LOOP_and_451_nl, 4'b1111,
      COMP_LOOP_or_41_nl);
  assign COMP_LOOP_mux1h_843_nl = MUX1HOT_v_6_3_2((STAGE_VEC_LOOP_j_sva_9_0[5:0]),
      (~ (STAGE_MAIN_LOOP_lshift_psp_1_sva[9:4])), ({1'b0 , COMP_LOOP_k_9_4_sva_4_0}),
      {and_dcpl_582 , and_dcpl_589 , and_dcpl_599});
  assign COMP_LOOP_or_42_nl = MUX_v_6_2_2(COMP_LOOP_mux1h_843_nl, 6'b111111, and_dcpl_593);
  assign COMP_LOOP_or_43_nl = (~(and_dcpl_582 | and_dcpl_593 | and_dcpl_599)) | and_dcpl_589;
  assign COMP_LOOP_nor_626_nl = ~(and_dcpl_589 | and_dcpl_593 | and_dcpl_599);
  assign COMP_LOOP_COMP_LOOP_and_992_nl = MUX_v_3_2_2(3'b000, (COMP_LOOP_k_9_4_sva_4_0[4:2]),
      COMP_LOOP_nor_626_nl);
  assign COMP_LOOP_mux_294_nl = MUX_v_2_2_2((COMP_LOOP_k_9_4_sva_4_0[1:0]), (COMP_LOOP_k_9_4_sva_4_0[4:3]),
      and_dcpl_589);
  assign COMP_LOOP_nor_627_nl = ~(and_dcpl_593 | and_dcpl_599);
  assign COMP_LOOP_COMP_LOOP_and_993_nl = MUX_v_2_2_2(2'b00, COMP_LOOP_mux_294_nl,
      COMP_LOOP_nor_627_nl);
  assign COMP_LOOP_mux1h_844_nl = MUX1HOT_v_3_3_2(3'b010, (COMP_LOOP_k_9_4_sva_4_0[2:0]),
      (STAGE_MAIN_LOOP_acc_1_psp_sva[3:1]), {and_dcpl_582 , and_dcpl_589 , and_dcpl_593});
  assign not_7304_nl = ~ and_dcpl_599;
  assign COMP_LOOP_and_452_nl = MUX_v_3_2_2(3'b000, COMP_LOOP_mux1h_844_nl, not_7304_nl);
  assign COMP_LOOP_COMP_LOOP_or_5_nl = ((STAGE_MAIN_LOOP_acc_1_psp_sva[0]) & (~ and_dcpl_589))
      | and_dcpl_582 | and_dcpl_599;
  assign nl_acc_3_nl = conv_s2s_12_13({COMP_LOOP_COMP_LOOP_or_3_nl , COMP_LOOP_COMP_LOOP_or_4_nl
      , COMP_LOOP_or_42_nl , COMP_LOOP_or_43_nl}) + conv_u2s_10_13({COMP_LOOP_COMP_LOOP_and_992_nl
      , COMP_LOOP_COMP_LOOP_and_993_nl , COMP_LOOP_and_452_nl , COMP_LOOP_COMP_LOOP_or_5_nl
      , 1'b1});
  assign acc_3_nl = nl_acc_3_nl[12:0];
  assign COMP_LOOP_slc_acc_3_12_1_slc = readslicef_13_12_1(acc_3_nl);
  assign COMP_LOOP_mux1h_845_nl = MUX1HOT_s_1_16_2(COMP_LOOP_COMP_LOOP_nor_itm, COMP_LOOP_COMP_LOOP_nor_5_itm,
      COMP_LOOP_COMP_LOOP_nor_9_itm, COMP_LOOP_COMP_LOOP_nor_13_itm, COMP_LOOP_COMP_LOOP_nor_17_itm,
      COMP_LOOP_COMP_LOOP_nor_21_itm, COMP_LOOP_COMP_LOOP_nor_25_itm, COMP_LOOP_COMP_LOOP_nor_29_itm,
      COMP_LOOP_COMP_LOOP_nor_33_itm, COMP_LOOP_COMP_LOOP_nor_37_itm, COMP_LOOP_COMP_LOOP_nor_41_itm,
      COMP_LOOP_COMP_LOOP_nor_45_itm, COMP_LOOP_COMP_LOOP_nor_49_itm, COMP_LOOP_COMP_LOOP_nor_53_itm,
      COMP_LOOP_COMP_LOOP_nor_57_itm, COMP_LOOP_COMP_LOOP_nor_61_itm, {and_920_cse
      , and_925_cse , and_dcpl_621 , and_936_cse , and_940_cse , and_945_cse , and_950_cse
      , and_953_cse , and_957_cse , and_960_cse , and_964_cse , and_966_cse , and_970_cse
      , and_973_cse , and_975_cse , and_978_cse});
  assign COMP_LOOP_COMP_LOOP_and_994_nl = (operator_64_false_acc_cse_2_sva[0]) &
      COMP_LOOP_nor_51_itm;
  assign COMP_LOOP_COMP_LOOP_and_995_nl = (operator_64_false_acc_cse_3_sva[0]) &
      COMP_LOOP_nor_91_itm;
  assign COMP_LOOP_COMP_LOOP_and_996_nl = (operator_64_false_acc_cse_4_sva[0]) &
      COMP_LOOP_nor_131_itm;
  assign COMP_LOOP_COMP_LOOP_and_997_nl = (operator_64_false_acc_cse_5_sva[0]) &
      COMP_LOOP_nor_171_itm;
  assign COMP_LOOP_COMP_LOOP_and_998_nl = (operator_64_false_acc_cse_6_sva[0]) &
      COMP_LOOP_nor_211_itm;
  assign COMP_LOOP_COMP_LOOP_and_999_nl = (operator_64_false_acc_cse_7_sva[0]) &
      COMP_LOOP_nor_251_itm;
  assign COMP_LOOP_COMP_LOOP_and_1000_nl = (operator_64_false_acc_cse_8_sva[0]) &
      COMP_LOOP_nor_291_itm;
  assign COMP_LOOP_COMP_LOOP_and_1001_nl = (operator_64_false_acc_cse_9_sva[0]) &
      COMP_LOOP_nor_331_itm;
  assign COMP_LOOP_COMP_LOOP_and_1002_nl = (operator_64_false_acc_cse_10_sva[0])
      & COMP_LOOP_nor_371_itm;
  assign COMP_LOOP_COMP_LOOP_and_1003_nl = (operator_64_false_acc_cse_11_sva[0])
      & COMP_LOOP_nor_411_itm;
  assign COMP_LOOP_COMP_LOOP_and_1004_nl = (operator_64_false_acc_cse_12_sva[0])
      & COMP_LOOP_nor_451_itm;
  assign COMP_LOOP_COMP_LOOP_and_1005_nl = (operator_64_false_acc_cse_13_sva[0])
      & COMP_LOOP_nor_491_itm;
  assign COMP_LOOP_COMP_LOOP_and_1006_nl = (operator_64_false_acc_cse_14_sva[0])
      & COMP_LOOP_nor_531_itm;
  assign COMP_LOOP_COMP_LOOP_and_1007_nl = (operator_64_false_acc_cse_15_sva[0])
      & COMP_LOOP_nor_571_itm;
  assign COMP_LOOP_COMP_LOOP_and_1008_nl = (operator_64_false_acc_cse_sva[0]) & COMP_LOOP_nor_611_itm;
  assign COMP_LOOP_mux1h_846_nl = MUX1HOT_s_1_16_2(COMP_LOOP_COMP_LOOP_and_244_itm,
      COMP_LOOP_COMP_LOOP_and_994_nl, COMP_LOOP_COMP_LOOP_and_995_nl, COMP_LOOP_COMP_LOOP_and_996_nl,
      COMP_LOOP_COMP_LOOP_and_997_nl, COMP_LOOP_COMP_LOOP_and_998_nl, COMP_LOOP_COMP_LOOP_and_999_nl,
      COMP_LOOP_COMP_LOOP_and_1000_nl, COMP_LOOP_COMP_LOOP_and_1001_nl, COMP_LOOP_COMP_LOOP_and_1002_nl,
      COMP_LOOP_COMP_LOOP_and_1003_nl, COMP_LOOP_COMP_LOOP_and_1004_nl, COMP_LOOP_COMP_LOOP_and_1005_nl,
      COMP_LOOP_COMP_LOOP_and_1006_nl, COMP_LOOP_COMP_LOOP_and_1007_nl, COMP_LOOP_COMP_LOOP_and_1008_nl,
      {and_920_cse , and_925_cse , and_dcpl_621 , and_936_cse , and_940_cse , and_945_cse
      , and_950_cse , and_953_cse , and_957_cse , and_960_cse , and_964_cse , and_966_cse
      , and_970_cse , and_973_cse , and_975_cse , and_978_cse});
  assign COMP_LOOP_COMP_LOOP_and_1009_nl = (operator_64_false_acc_cse_2_sva[1]) &
      COMP_LOOP_nor_52_itm;
  assign COMP_LOOP_COMP_LOOP_and_1010_nl = (operator_64_false_acc_cse_3_sva[1]) &
      COMP_LOOP_nor_92_itm;
  assign COMP_LOOP_COMP_LOOP_and_1011_nl = (operator_64_false_acc_cse_4_sva[1]) &
      COMP_LOOP_nor_132_itm;
  assign COMP_LOOP_COMP_LOOP_and_1012_nl = (operator_64_false_acc_cse_5_sva[1]) &
      COMP_LOOP_nor_172_itm;
  assign COMP_LOOP_COMP_LOOP_and_1013_nl = (operator_64_false_acc_cse_6_sva[1]) &
      COMP_LOOP_nor_212_itm;
  assign COMP_LOOP_COMP_LOOP_and_1014_nl = (operator_64_false_acc_cse_7_sva[1]) &
      COMP_LOOP_nor_252_itm;
  assign COMP_LOOP_COMP_LOOP_and_1015_nl = (operator_64_false_acc_cse_8_sva[1]) &
      COMP_LOOP_nor_292_itm;
  assign COMP_LOOP_COMP_LOOP_and_1016_nl = (operator_64_false_acc_cse_9_sva[1]) &
      COMP_LOOP_nor_332_itm;
  assign COMP_LOOP_COMP_LOOP_and_1017_nl = (operator_64_false_acc_cse_10_sva[1])
      & COMP_LOOP_nor_372_itm;
  assign COMP_LOOP_COMP_LOOP_and_1018_nl = (operator_64_false_acc_cse_11_sva[1])
      & COMP_LOOP_nor_412_itm;
  assign COMP_LOOP_COMP_LOOP_and_1019_nl = (operator_64_false_acc_cse_12_sva[1])
      & COMP_LOOP_nor_452_itm;
  assign COMP_LOOP_COMP_LOOP_and_1020_nl = (operator_64_false_acc_cse_13_sva[1])
      & COMP_LOOP_nor_492_itm;
  assign COMP_LOOP_COMP_LOOP_and_1021_nl = (operator_64_false_acc_cse_14_sva[1])
      & COMP_LOOP_nor_532_itm;
  assign COMP_LOOP_COMP_LOOP_and_1022_nl = (operator_64_false_acc_cse_15_sva[1])
      & COMP_LOOP_nor_572_itm;
  assign COMP_LOOP_COMP_LOOP_and_1023_nl = (operator_64_false_acc_cse_sva[1]) & COMP_LOOP_nor_612_itm;
  assign COMP_LOOP_mux1h_847_nl = MUX1HOT_s_1_16_2(COMP_LOOP_COMP_LOOP_and_62_itm,
      COMP_LOOP_COMP_LOOP_and_1009_nl, COMP_LOOP_COMP_LOOP_and_1010_nl, COMP_LOOP_COMP_LOOP_and_1011_nl,
      COMP_LOOP_COMP_LOOP_and_1012_nl, COMP_LOOP_COMP_LOOP_and_1013_nl, COMP_LOOP_COMP_LOOP_and_1014_nl,
      COMP_LOOP_COMP_LOOP_and_1015_nl, COMP_LOOP_COMP_LOOP_and_1016_nl, COMP_LOOP_COMP_LOOP_and_1017_nl,
      COMP_LOOP_COMP_LOOP_and_1018_nl, COMP_LOOP_COMP_LOOP_and_1019_nl, COMP_LOOP_COMP_LOOP_and_1020_nl,
      COMP_LOOP_COMP_LOOP_and_1021_nl, COMP_LOOP_COMP_LOOP_and_1022_nl, COMP_LOOP_COMP_LOOP_and_1023_nl,
      {and_920_cse , and_925_cse , and_dcpl_621 , and_936_cse , and_940_cse , and_945_cse
      , and_950_cse , and_953_cse , and_957_cse , and_960_cse , and_964_cse , and_966_cse
      , and_970_cse , and_973_cse , and_975_cse , and_978_cse});
  assign COMP_LOOP_mux1h_848_nl = MUX1HOT_s_1_16_2(COMP_LOOP_COMP_LOOP_and_185_itm,
      COMP_LOOP_COMP_LOOP_and_77_itm, COMP_LOOP_COMP_LOOP_and_137_itm, COMP_LOOP_COMP_LOOP_and_197_itm,
      COMP_LOOP_COMP_LOOP_and_257_itm, COMP_LOOP_COMP_LOOP_and_317_itm, COMP_LOOP_COMP_LOOP_and_377_itm,
      COMP_LOOP_COMP_LOOP_and_437_itm, COMP_LOOP_COMP_LOOP_and_497_itm, COMP_LOOP_COMP_LOOP_and_557_itm,
      COMP_LOOP_COMP_LOOP_and_617_itm, COMP_LOOP_COMP_LOOP_and_677_itm, COMP_LOOP_COMP_LOOP_and_737_itm,
      COMP_LOOP_COMP_LOOP_and_797_itm, COMP_LOOP_COMP_LOOP_and_857_itm, COMP_LOOP_COMP_LOOP_and_917_itm,
      {and_920_cse , and_925_cse , and_dcpl_621 , and_936_cse , and_940_cse , and_945_cse
      , and_950_cse , and_953_cse , and_957_cse , and_960_cse , and_964_cse , and_966_cse
      , and_970_cse , and_973_cse , and_975_cse , and_978_cse});
  assign COMP_LOOP_COMP_LOOP_and_1024_nl = (operator_64_false_acc_cse_2_sva[2]) &
      COMP_LOOP_nor_54_itm;
  assign COMP_LOOP_COMP_LOOP_and_1025_nl = (operator_64_false_acc_cse_3_sva[2]) &
      COMP_LOOP_nor_94_itm;
  assign COMP_LOOP_COMP_LOOP_and_1026_nl = (operator_64_false_acc_cse_4_sva[2]) &
      COMP_LOOP_nor_134_itm;
  assign COMP_LOOP_COMP_LOOP_and_1027_nl = (operator_64_false_acc_cse_5_sva[2]) &
      COMP_LOOP_nor_174_itm;
  assign COMP_LOOP_COMP_LOOP_and_1028_nl = (operator_64_false_acc_cse_6_sva[2]) &
      COMP_LOOP_nor_214_itm;
  assign COMP_LOOP_COMP_LOOP_and_1029_nl = (operator_64_false_acc_cse_7_sva[2]) &
      COMP_LOOP_nor_254_itm;
  assign COMP_LOOP_COMP_LOOP_and_1030_nl = (operator_64_false_acc_cse_8_sva[2]) &
      COMP_LOOP_nor_294_itm;
  assign COMP_LOOP_COMP_LOOP_and_1031_nl = (operator_64_false_acc_cse_9_sva[2]) &
      COMP_LOOP_nor_334_itm;
  assign COMP_LOOP_COMP_LOOP_and_1032_nl = (operator_64_false_acc_cse_10_sva[2])
      & COMP_LOOP_nor_374_itm;
  assign COMP_LOOP_COMP_LOOP_and_1033_nl = (operator_64_false_acc_cse_11_sva[2])
      & COMP_LOOP_nor_414_itm;
  assign COMP_LOOP_COMP_LOOP_and_1034_nl = (operator_64_false_acc_cse_12_sva[2])
      & COMP_LOOP_nor_454_itm;
  assign COMP_LOOP_COMP_LOOP_and_1035_nl = (operator_64_false_acc_cse_13_sva[2])
      & COMP_LOOP_nor_494_itm;
  assign COMP_LOOP_COMP_LOOP_and_1036_nl = (operator_64_false_acc_cse_14_sva[2])
      & COMP_LOOP_nor_534_itm;
  assign COMP_LOOP_COMP_LOOP_and_1037_nl = (operator_64_false_acc_cse_15_sva[2])
      & COMP_LOOP_nor_574_itm;
  assign COMP_LOOP_COMP_LOOP_and_1038_nl = (operator_64_false_acc_cse_sva[2]) & COMP_LOOP_nor_614_itm;
  assign COMP_LOOP_mux1h_849_nl = MUX1HOT_s_1_16_2(COMP_LOOP_COMP_LOOP_and_64_itm,
      COMP_LOOP_COMP_LOOP_and_1024_nl, COMP_LOOP_COMP_LOOP_and_1025_nl, COMP_LOOP_COMP_LOOP_and_1026_nl,
      COMP_LOOP_COMP_LOOP_and_1027_nl, COMP_LOOP_COMP_LOOP_and_1028_nl, COMP_LOOP_COMP_LOOP_and_1029_nl,
      COMP_LOOP_COMP_LOOP_and_1030_nl, COMP_LOOP_COMP_LOOP_and_1031_nl, COMP_LOOP_COMP_LOOP_and_1032_nl,
      COMP_LOOP_COMP_LOOP_and_1033_nl, COMP_LOOP_COMP_LOOP_and_1034_nl, COMP_LOOP_COMP_LOOP_and_1035_nl,
      COMP_LOOP_COMP_LOOP_and_1036_nl, COMP_LOOP_COMP_LOOP_and_1037_nl, COMP_LOOP_COMP_LOOP_and_1038_nl,
      {and_920_cse , and_925_cse , and_dcpl_621 , and_936_cse , and_940_cse , and_945_cse
      , and_950_cse , and_953_cse , and_957_cse , and_960_cse , and_964_cse , and_966_cse
      , and_970_cse , and_973_cse , and_975_cse , and_978_cse});
  assign COMP_LOOP_mux1h_850_nl = MUX1HOT_s_1_16_2(COMP_LOOP_COMP_LOOP_and_65_itm,
      COMP_LOOP_COMP_LOOP_and_79_itm, COMP_LOOP_COMP_LOOP_and_139_itm, COMP_LOOP_COMP_LOOP_and_199_itm,
      COMP_LOOP_COMP_LOOP_and_259_itm, COMP_LOOP_COMP_LOOP_and_319_itm, COMP_LOOP_COMP_LOOP_and_379_itm,
      COMP_LOOP_COMP_LOOP_and_439_itm, COMP_LOOP_COMP_LOOP_and_499_itm, COMP_LOOP_COMP_LOOP_and_559_itm,
      COMP_LOOP_COMP_LOOP_and_619_itm, COMP_LOOP_COMP_LOOP_and_679_itm, COMP_LOOP_COMP_LOOP_and_739_itm,
      COMP_LOOP_COMP_LOOP_and_799_itm, COMP_LOOP_COMP_LOOP_and_859_itm, COMP_LOOP_COMP_LOOP_and_919_itm,
      {and_920_cse , and_925_cse , and_dcpl_621 , and_936_cse , and_940_cse , and_945_cse
      , and_950_cse , and_953_cse , and_957_cse , and_960_cse , and_964_cse , and_966_cse
      , and_970_cse , and_973_cse , and_975_cse , and_978_cse});
  assign COMP_LOOP_mux1h_851_nl = MUX1HOT_s_1_16_2(COMP_LOOP_COMP_LOOP_and_66_itm,
      COMP_LOOP_COMP_LOOP_and_80_itm, COMP_LOOP_COMP_LOOP_and_140_itm, COMP_LOOP_COMP_LOOP_and_200_itm,
      COMP_LOOP_COMP_LOOP_and_260_itm, COMP_LOOP_COMP_LOOP_and_320_itm, COMP_LOOP_COMP_LOOP_and_380_itm,
      COMP_LOOP_COMP_LOOP_and_440_itm, COMP_LOOP_COMP_LOOP_and_500_itm, COMP_LOOP_COMP_LOOP_and_560_itm,
      COMP_LOOP_COMP_LOOP_and_620_itm, COMP_LOOP_COMP_LOOP_and_680_itm, COMP_LOOP_COMP_LOOP_and_740_itm,
      COMP_LOOP_COMP_LOOP_and_800_itm, COMP_LOOP_COMP_LOOP_and_860_itm, COMP_LOOP_COMP_LOOP_and_920_itm,
      {and_920_cse , and_925_cse , and_dcpl_621 , and_936_cse , and_940_cse , and_945_cse
      , and_950_cse , and_953_cse , and_957_cse , and_960_cse , and_964_cse , and_966_cse
      , and_970_cse , and_973_cse , and_975_cse , and_978_cse});
  assign COMP_LOOP_mux1h_852_nl = MUX1HOT_s_1_16_2(COMP_LOOP_COMP_LOOP_and_6_itm,
      COMP_LOOP_COMP_LOOP_and_81_itm, COMP_LOOP_COMP_LOOP_and_141_itm, COMP_LOOP_COMP_LOOP_and_201_itm,
      COMP_LOOP_COMP_LOOP_and_261_itm, COMP_LOOP_COMP_LOOP_and_321_itm, COMP_LOOP_COMP_LOOP_and_381_itm,
      COMP_LOOP_COMP_LOOP_and_441_itm, COMP_LOOP_COMP_LOOP_and_501_itm, COMP_LOOP_COMP_LOOP_and_561_itm,
      COMP_LOOP_COMP_LOOP_and_621_itm, COMP_LOOP_COMP_LOOP_and_681_itm, COMP_LOOP_COMP_LOOP_and_741_itm,
      COMP_LOOP_COMP_LOOP_and_801_itm, COMP_LOOP_COMP_LOOP_and_861_itm, COMP_LOOP_COMP_LOOP_and_921_itm,
      {and_920_cse , and_925_cse , and_dcpl_621 , and_936_cse , and_940_cse , and_945_cse
      , and_950_cse , and_953_cse , and_957_cse , and_960_cse , and_964_cse , and_966_cse
      , and_970_cse , and_973_cse , and_975_cse , and_978_cse});
  assign COMP_LOOP_COMP_LOOP_and_1039_nl = (operator_64_false_acc_cse_2_sva[3]) &
      COMP_LOOP_nor_57_itm;
  assign COMP_LOOP_COMP_LOOP_and_1040_nl = (operator_64_false_acc_cse_3_sva[3]) &
      COMP_LOOP_nor_97_itm;
  assign COMP_LOOP_COMP_LOOP_and_1041_nl = (operator_64_false_acc_cse_4_sva[3]) &
      COMP_LOOP_nor_137_itm;
  assign COMP_LOOP_COMP_LOOP_and_1042_nl = (operator_64_false_acc_cse_5_sva[3]) &
      COMP_LOOP_nor_177_itm;
  assign COMP_LOOP_COMP_LOOP_and_1043_nl = (operator_64_false_acc_cse_6_sva[3]) &
      COMP_LOOP_nor_217_itm;
  assign COMP_LOOP_COMP_LOOP_and_1044_nl = (operator_64_false_acc_cse_7_sva[3]) &
      COMP_LOOP_nor_257_itm;
  assign COMP_LOOP_COMP_LOOP_and_1045_nl = (operator_64_false_acc_cse_8_sva[3]) &
      COMP_LOOP_nor_297_itm;
  assign COMP_LOOP_COMP_LOOP_and_1046_nl = (operator_64_false_acc_cse_9_sva[3]) &
      COMP_LOOP_nor_337_itm;
  assign COMP_LOOP_COMP_LOOP_and_1047_nl = (operator_64_false_acc_cse_10_sva[3])
      & COMP_LOOP_nor_377_itm;
  assign COMP_LOOP_COMP_LOOP_and_1048_nl = (operator_64_false_acc_cse_11_sva[3])
      & COMP_LOOP_nor_417_itm;
  assign COMP_LOOP_COMP_LOOP_and_1049_nl = (operator_64_false_acc_cse_12_sva[3])
      & COMP_LOOP_nor_457_itm;
  assign COMP_LOOP_COMP_LOOP_and_1050_nl = (operator_64_false_acc_cse_13_sva[3])
      & COMP_LOOP_nor_497_itm;
  assign COMP_LOOP_COMP_LOOP_and_1051_nl = (operator_64_false_acc_cse_14_sva[3])
      & COMP_LOOP_nor_537_itm;
  assign COMP_LOOP_COMP_LOOP_and_1052_nl = (operator_64_false_acc_cse_15_sva[3])
      & COMP_LOOP_nor_577_itm;
  assign COMP_LOOP_COMP_LOOP_and_1053_nl = (operator_64_false_acc_cse_sva[3]) & COMP_LOOP_nor_617_itm;
  assign COMP_LOOP_mux1h_853_nl = MUX1HOT_s_1_16_2(COMP_LOOP_COMP_LOOP_and_68_itm,
      COMP_LOOP_COMP_LOOP_and_1039_nl, COMP_LOOP_COMP_LOOP_and_1040_nl, COMP_LOOP_COMP_LOOP_and_1041_nl,
      COMP_LOOP_COMP_LOOP_and_1042_nl, COMP_LOOP_COMP_LOOP_and_1043_nl, COMP_LOOP_COMP_LOOP_and_1044_nl,
      COMP_LOOP_COMP_LOOP_and_1045_nl, COMP_LOOP_COMP_LOOP_and_1046_nl, COMP_LOOP_COMP_LOOP_and_1047_nl,
      COMP_LOOP_COMP_LOOP_and_1048_nl, COMP_LOOP_COMP_LOOP_and_1049_nl, COMP_LOOP_COMP_LOOP_and_1050_nl,
      COMP_LOOP_COMP_LOOP_and_1051_nl, COMP_LOOP_COMP_LOOP_and_1052_nl, COMP_LOOP_COMP_LOOP_and_1053_nl,
      {and_920_cse , and_925_cse , and_dcpl_621 , and_936_cse , and_940_cse , and_945_cse
      , and_950_cse , and_953_cse , and_957_cse , and_960_cse , and_964_cse , and_966_cse
      , and_970_cse , and_973_cse , and_975_cse , and_978_cse});
  assign COMP_LOOP_mux1h_854_nl = MUX1HOT_s_1_16_2(COMP_LOOP_COMP_LOOP_and_69_itm,
      COMP_LOOP_COMP_LOOP_and_83_itm, COMP_LOOP_COMP_LOOP_and_143_itm, COMP_LOOP_COMP_LOOP_and_203_itm,
      COMP_LOOP_COMP_LOOP_and_263_itm, COMP_LOOP_COMP_LOOP_and_323_itm, COMP_LOOP_COMP_LOOP_and_383_itm,
      COMP_LOOP_COMP_LOOP_and_443_itm, COMP_LOOP_COMP_LOOP_and_503_itm, COMP_LOOP_COMP_LOOP_and_563_itm,
      COMP_LOOP_COMP_LOOP_and_623_itm, COMP_LOOP_COMP_LOOP_and_683_itm, COMP_LOOP_COMP_LOOP_and_743_itm,
      COMP_LOOP_COMP_LOOP_and_803_itm, COMP_LOOP_COMP_LOOP_and_863_itm, COMP_LOOP_COMP_LOOP_and_923_itm,
      {and_920_cse , and_925_cse , and_dcpl_621 , and_936_cse , and_940_cse , and_945_cse
      , and_950_cse , and_953_cse , and_957_cse , and_960_cse , and_964_cse , and_966_cse
      , and_970_cse , and_973_cse , and_975_cse , and_978_cse});
  assign COMP_LOOP_mux1h_855_nl = MUX1HOT_s_1_16_2(COMP_LOOP_COMP_LOOP_and_70_itm,
      COMP_LOOP_COMP_LOOP_and_84_itm, COMP_LOOP_COMP_LOOP_and_144_itm, COMP_LOOP_COMP_LOOP_and_204_itm,
      COMP_LOOP_COMP_LOOP_and_264_itm, COMP_LOOP_COMP_LOOP_and_324_itm, COMP_LOOP_COMP_LOOP_and_384_itm,
      COMP_LOOP_COMP_LOOP_and_444_itm, COMP_LOOP_COMP_LOOP_and_504_itm, COMP_LOOP_COMP_LOOP_and_564_itm,
      COMP_LOOP_COMP_LOOP_and_624_itm, COMP_LOOP_COMP_LOOP_and_684_itm, COMP_LOOP_COMP_LOOP_and_744_itm,
      COMP_LOOP_COMP_LOOP_and_804_itm, COMP_LOOP_COMP_LOOP_and_864_itm, COMP_LOOP_COMP_LOOP_and_924_itm,
      {and_920_cse , and_925_cse , and_dcpl_621 , and_936_cse , and_940_cse , and_945_cse
      , and_950_cse , and_953_cse , and_957_cse , and_960_cse , and_964_cse , and_966_cse
      , and_970_cse , and_973_cse , and_975_cse , and_978_cse});
  assign COMP_LOOP_mux1h_856_nl = MUX1HOT_s_1_16_2(COMP_LOOP_COMP_LOOP_and_10_itm,
      COMP_LOOP_COMP_LOOP_and_85_itm, COMP_LOOP_COMP_LOOP_and_145_itm, COMP_LOOP_COMP_LOOP_and_205_itm,
      COMP_LOOP_COMP_LOOP_and_265_itm, COMP_LOOP_COMP_LOOP_and_325_itm, COMP_LOOP_COMP_LOOP_and_385_itm,
      COMP_LOOP_COMP_LOOP_and_445_itm, COMP_LOOP_COMP_LOOP_and_505_itm, COMP_LOOP_COMP_LOOP_and_565_itm,
      COMP_LOOP_COMP_LOOP_and_625_itm, COMP_LOOP_COMP_LOOP_and_685_itm, COMP_LOOP_COMP_LOOP_and_745_itm,
      COMP_LOOP_COMP_LOOP_and_805_itm, COMP_LOOP_COMP_LOOP_and_865_itm, COMP_LOOP_COMP_LOOP_and_925_itm,
      {and_920_cse , and_925_cse , and_dcpl_621 , and_936_cse , and_940_cse , and_945_cse
      , and_950_cse , and_953_cse , and_957_cse , and_960_cse , and_964_cse , and_966_cse
      , and_970_cse , and_973_cse , and_975_cse , and_978_cse});
  assign COMP_LOOP_mux1h_857_nl = MUX1HOT_s_1_16_2(COMP_LOOP_COMP_LOOP_and_72_itm,
      COMP_LOOP_COMP_LOOP_and_86_itm, COMP_LOOP_COMP_LOOP_and_146_itm, COMP_LOOP_COMP_LOOP_and_206_itm,
      COMP_LOOP_COMP_LOOP_and_266_itm, COMP_LOOP_COMP_LOOP_and_326_itm, COMP_LOOP_COMP_LOOP_and_386_itm,
      COMP_LOOP_COMP_LOOP_and_446_itm, COMP_LOOP_COMP_LOOP_and_506_itm, COMP_LOOP_COMP_LOOP_and_566_itm,
      COMP_LOOP_COMP_LOOP_and_626_itm, COMP_LOOP_COMP_LOOP_and_686_itm, COMP_LOOP_COMP_LOOP_and_746_itm,
      COMP_LOOP_COMP_LOOP_and_806_itm, COMP_LOOP_COMP_LOOP_and_866_itm, COMP_LOOP_COMP_LOOP_and_926_itm,
      {and_920_cse , and_925_cse , and_dcpl_621 , and_936_cse , and_940_cse , and_945_cse
      , and_950_cse , and_953_cse , and_957_cse , and_960_cse , and_964_cse , and_966_cse
      , and_970_cse , and_973_cse , and_975_cse , and_978_cse});
  assign COMP_LOOP_mux1h_858_nl = MUX1HOT_s_1_16_2(COMP_LOOP_COMP_LOOP_and_12_itm,
      COMP_LOOP_COMP_LOOP_and_87_itm, COMP_LOOP_COMP_LOOP_and_147_itm, COMP_LOOP_COMP_LOOP_and_207_itm,
      COMP_LOOP_COMP_LOOP_and_267_itm, COMP_LOOP_COMP_LOOP_and_327_itm, COMP_LOOP_COMP_LOOP_and_387_itm,
      COMP_LOOP_COMP_LOOP_and_447_itm, COMP_LOOP_COMP_LOOP_and_507_itm, COMP_LOOP_COMP_LOOP_and_567_itm,
      COMP_LOOP_COMP_LOOP_and_627_itm, COMP_LOOP_COMP_LOOP_and_687_itm, COMP_LOOP_COMP_LOOP_and_747_itm,
      COMP_LOOP_COMP_LOOP_and_807_itm, COMP_LOOP_COMP_LOOP_and_867_itm, COMP_LOOP_COMP_LOOP_and_927_itm,
      {and_920_cse , and_925_cse , and_dcpl_621 , and_936_cse , and_940_cse , and_945_cse
      , and_950_cse , and_953_cse , and_957_cse , and_960_cse , and_964_cse , and_966_cse
      , and_970_cse , and_973_cse , and_975_cse , and_978_cse});
  assign COMP_LOOP_mux1h_859_nl = MUX1HOT_s_1_16_2(COMP_LOOP_COMP_LOOP_and_13_itm,
      COMP_LOOP_COMP_LOOP_and_88_itm, COMP_LOOP_COMP_LOOP_and_148_itm, COMP_LOOP_COMP_LOOP_and_208_itm,
      COMP_LOOP_COMP_LOOP_and_268_itm, COMP_LOOP_COMP_LOOP_and_328_itm, COMP_LOOP_COMP_LOOP_and_388_itm,
      COMP_LOOP_COMP_LOOP_and_448_itm, COMP_LOOP_COMP_LOOP_and_508_itm, COMP_LOOP_COMP_LOOP_and_568_itm,
      COMP_LOOP_COMP_LOOP_and_628_itm, COMP_LOOP_COMP_LOOP_and_688_itm, COMP_LOOP_COMP_LOOP_and_748_itm,
      COMP_LOOP_COMP_LOOP_and_808_itm, COMP_LOOP_COMP_LOOP_and_868_itm, COMP_LOOP_COMP_LOOP_and_928_itm,
      {and_920_cse , and_925_cse , and_dcpl_621 , and_936_cse , and_940_cse , and_945_cse
      , and_950_cse , and_953_cse , and_957_cse , and_960_cse , and_964_cse , and_966_cse
      , and_970_cse , and_973_cse , and_975_cse , and_978_cse});
  assign COMP_LOOP_mux1h_860_nl = MUX1HOT_s_1_16_2(COMP_LOOP_COMP_LOOP_and_14_itm,
      COMP_LOOP_COMP_LOOP_and_89_itm, COMP_LOOP_COMP_LOOP_and_149_itm, COMP_LOOP_COMP_LOOP_and_209_itm,
      COMP_LOOP_COMP_LOOP_and_269_itm, COMP_LOOP_COMP_LOOP_and_329_itm, COMP_LOOP_COMP_LOOP_and_389_itm,
      COMP_LOOP_COMP_LOOP_and_449_itm, COMP_LOOP_COMP_LOOP_and_509_itm, COMP_LOOP_COMP_LOOP_and_569_itm,
      COMP_LOOP_COMP_LOOP_and_629_itm, COMP_LOOP_COMP_LOOP_and_689_itm, COMP_LOOP_COMP_LOOP_and_749_itm,
      COMP_LOOP_COMP_LOOP_and_809_itm, COMP_LOOP_COMP_LOOP_and_869_itm, COMP_LOOP_COMP_LOOP_and_929_itm,
      {and_920_cse , and_925_cse , and_dcpl_621 , and_936_cse , and_940_cse , and_945_cse
      , and_950_cse , and_953_cse , and_957_cse , and_960_cse , and_964_cse , and_966_cse
      , and_970_cse , and_973_cse , and_975_cse , and_978_cse});
  assign z_out_5 = MUX1HOT_v_64_16_2(vec_rsc_0_0_i_qa_d, vec_rsc_0_1_i_qa_d, vec_rsc_0_2_i_qa_d,
      vec_rsc_0_3_i_qa_d, vec_rsc_0_4_i_qa_d, vec_rsc_0_5_i_qa_d, vec_rsc_0_6_i_qa_d,
      vec_rsc_0_7_i_qa_d, vec_rsc_0_8_i_qa_d, vec_rsc_0_9_i_qa_d, vec_rsc_0_10_i_qa_d,
      vec_rsc_0_11_i_qa_d, vec_rsc_0_12_i_qa_d, vec_rsc_0_13_i_qa_d, vec_rsc_0_14_i_qa_d,
      vec_rsc_0_15_i_qa_d, {COMP_LOOP_mux1h_845_nl , COMP_LOOP_mux1h_846_nl , COMP_LOOP_mux1h_847_nl
      , COMP_LOOP_mux1h_848_nl , COMP_LOOP_mux1h_849_nl , COMP_LOOP_mux1h_850_nl
      , COMP_LOOP_mux1h_851_nl , COMP_LOOP_mux1h_852_nl , COMP_LOOP_mux1h_853_nl
      , COMP_LOOP_mux1h_854_nl , COMP_LOOP_mux1h_855_nl , COMP_LOOP_mux1h_856_nl
      , COMP_LOOP_mux1h_857_nl , COMP_LOOP_mux1h_858_nl , COMP_LOOP_mux1h_859_nl
      , COMP_LOOP_mux1h_860_nl});

  function automatic [0:0] MUX1HOT_s_1_16_2;
    input [0:0] input_15;
    input [0:0] input_14;
    input [0:0] input_13;
    input [0:0] input_12;
    input [0:0] input_11;
    input [0:0] input_10;
    input [0:0] input_9;
    input [0:0] input_8;
    input [0:0] input_7;
    input [0:0] input_6;
    input [0:0] input_5;
    input [0:0] input_4;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [15:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    result = result | ( input_4 & {1{sel[4]}});
    result = result | ( input_5 & {1{sel[5]}});
    result = result | ( input_6 & {1{sel[6]}});
    result = result | ( input_7 & {1{sel[7]}});
    result = result | ( input_8 & {1{sel[8]}});
    result = result | ( input_9 & {1{sel[9]}});
    result = result | ( input_10 & {1{sel[10]}});
    result = result | ( input_11 & {1{sel[11]}});
    result = result | ( input_12 & {1{sel[12]}});
    result = result | ( input_13 & {1{sel[13]}});
    result = result | ( input_14 & {1{sel[14]}});
    result = result | ( input_15 & {1{sel[15]}});
    MUX1HOT_s_1_16_2 = result;
  end
  endfunction


  function automatic [0:0] MUX1HOT_s_1_4_2;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [3:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    MUX1HOT_s_1_4_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_4_2;
    input [1:0] input_3;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [3:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | ( input_1 & {2{sel[1]}});
    result = result | ( input_2 & {2{sel[2]}});
    result = result | ( input_3 & {2{sel[3]}});
    MUX1HOT_v_2_4_2 = result;
  end
  endfunction


  function automatic [2:0] MUX1HOT_v_3_3_2;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [2:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | ( input_1 & {3{sel[1]}});
    result = result | ( input_2 & {3{sel[2]}});
    MUX1HOT_v_3_3_2 = result;
  end
  endfunction


  function automatic [2:0] MUX1HOT_v_3_4_2;
    input [2:0] input_3;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [3:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | ( input_1 & {3{sel[1]}});
    result = result | ( input_2 & {3{sel[2]}});
    result = result | ( input_3 & {3{sel[3]}});
    MUX1HOT_v_3_4_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_16_2;
    input [3:0] input_15;
    input [3:0] input_14;
    input [3:0] input_13;
    input [3:0] input_12;
    input [3:0] input_11;
    input [3:0] input_10;
    input [3:0] input_9;
    input [3:0] input_8;
    input [3:0] input_7;
    input [3:0] input_6;
    input [3:0] input_5;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [15:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | ( input_1 & {4{sel[1]}});
    result = result | ( input_2 & {4{sel[2]}});
    result = result | ( input_3 & {4{sel[3]}});
    result = result | ( input_4 & {4{sel[4]}});
    result = result | ( input_5 & {4{sel[5]}});
    result = result | ( input_6 & {4{sel[6]}});
    result = result | ( input_7 & {4{sel[7]}});
    result = result | ( input_8 & {4{sel[8]}});
    result = result | ( input_9 & {4{sel[9]}});
    result = result | ( input_10 & {4{sel[10]}});
    result = result | ( input_11 & {4{sel[11]}});
    result = result | ( input_12 & {4{sel[12]}});
    result = result | ( input_13 & {4{sel[13]}});
    result = result | ( input_14 & {4{sel[14]}});
    result = result | ( input_15 & {4{sel[15]}});
    MUX1HOT_v_4_16_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_16_2;
    input [63:0] input_15;
    input [63:0] input_14;
    input [63:0] input_13;
    input [63:0] input_12;
    input [63:0] input_11;
    input [63:0] input_10;
    input [63:0] input_9;
    input [63:0] input_8;
    input [63:0] input_7;
    input [63:0] input_6;
    input [63:0] input_5;
    input [63:0] input_4;
    input [63:0] input_3;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [15:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    result = result | ( input_3 & {64{sel[3]}});
    result = result | ( input_4 & {64{sel[4]}});
    result = result | ( input_5 & {64{sel[5]}});
    result = result | ( input_6 & {64{sel[6]}});
    result = result | ( input_7 & {64{sel[7]}});
    result = result | ( input_8 & {64{sel[8]}});
    result = result | ( input_9 & {64{sel[9]}});
    result = result | ( input_10 & {64{sel[10]}});
    result = result | ( input_11 & {64{sel[11]}});
    result = result | ( input_12 & {64{sel[12]}});
    result = result | ( input_13 & {64{sel[13]}});
    result = result | ( input_14 & {64{sel[14]}});
    result = result | ( input_15 & {64{sel[15]}});
    MUX1HOT_v_64_16_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_18_2;
    input [63:0] input_17;
    input [63:0] input_16;
    input [63:0] input_15;
    input [63:0] input_14;
    input [63:0] input_13;
    input [63:0] input_12;
    input [63:0] input_11;
    input [63:0] input_10;
    input [63:0] input_9;
    input [63:0] input_8;
    input [63:0] input_7;
    input [63:0] input_6;
    input [63:0] input_5;
    input [63:0] input_4;
    input [63:0] input_3;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [17:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    result = result | ( input_3 & {64{sel[3]}});
    result = result | ( input_4 & {64{sel[4]}});
    result = result | ( input_5 & {64{sel[5]}});
    result = result | ( input_6 & {64{sel[6]}});
    result = result | ( input_7 & {64{sel[7]}});
    result = result | ( input_8 & {64{sel[8]}});
    result = result | ( input_9 & {64{sel[9]}});
    result = result | ( input_10 & {64{sel[10]}});
    result = result | ( input_11 & {64{sel[11]}});
    result = result | ( input_12 & {64{sel[12]}});
    result = result | ( input_13 & {64{sel[13]}});
    result = result | ( input_14 & {64{sel[14]}});
    result = result | ( input_15 & {64{sel[15]}});
    result = result | ( input_16 & {64{sel[16]}});
    result = result | ( input_17 & {64{sel[17]}});
    MUX1HOT_v_64_18_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_3_2;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [2:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    MUX1HOT_v_64_3_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_4_2;
    input [63:0] input_3;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [3:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    result = result | ( input_3 & {64{sel[3]}});
    MUX1HOT_v_64_4_2 = result;
  end
  endfunction


  function automatic [5:0] MUX1HOT_v_6_33_2;
    input [5:0] input_32;
    input [5:0] input_31;
    input [5:0] input_30;
    input [5:0] input_29;
    input [5:0] input_28;
    input [5:0] input_27;
    input [5:0] input_26;
    input [5:0] input_25;
    input [5:0] input_24;
    input [5:0] input_23;
    input [5:0] input_22;
    input [5:0] input_21;
    input [5:0] input_20;
    input [5:0] input_19;
    input [5:0] input_18;
    input [5:0] input_17;
    input [5:0] input_16;
    input [5:0] input_15;
    input [5:0] input_14;
    input [5:0] input_13;
    input [5:0] input_12;
    input [5:0] input_11;
    input [5:0] input_10;
    input [5:0] input_9;
    input [5:0] input_8;
    input [5:0] input_7;
    input [5:0] input_6;
    input [5:0] input_5;
    input [5:0] input_4;
    input [5:0] input_3;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [32:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | ( input_1 & {6{sel[1]}});
    result = result | ( input_2 & {6{sel[2]}});
    result = result | ( input_3 & {6{sel[3]}});
    result = result | ( input_4 & {6{sel[4]}});
    result = result | ( input_5 & {6{sel[5]}});
    result = result | ( input_6 & {6{sel[6]}});
    result = result | ( input_7 & {6{sel[7]}});
    result = result | ( input_8 & {6{sel[8]}});
    result = result | ( input_9 & {6{sel[9]}});
    result = result | ( input_10 & {6{sel[10]}});
    result = result | ( input_11 & {6{sel[11]}});
    result = result | ( input_12 & {6{sel[12]}});
    result = result | ( input_13 & {6{sel[13]}});
    result = result | ( input_14 & {6{sel[14]}});
    result = result | ( input_15 & {6{sel[15]}});
    result = result | ( input_16 & {6{sel[16]}});
    result = result | ( input_17 & {6{sel[17]}});
    result = result | ( input_18 & {6{sel[18]}});
    result = result | ( input_19 & {6{sel[19]}});
    result = result | ( input_20 & {6{sel[20]}});
    result = result | ( input_21 & {6{sel[21]}});
    result = result | ( input_22 & {6{sel[22]}});
    result = result | ( input_23 & {6{sel[23]}});
    result = result | ( input_24 & {6{sel[24]}});
    result = result | ( input_25 & {6{sel[25]}});
    result = result | ( input_26 & {6{sel[26]}});
    result = result | ( input_27 & {6{sel[27]}});
    result = result | ( input_28 & {6{sel[28]}});
    result = result | ( input_29 & {6{sel[29]}});
    result = result | ( input_30 & {6{sel[30]}});
    result = result | ( input_31 & {6{sel[31]}});
    result = result | ( input_32 & {6{sel[32]}});
    MUX1HOT_v_6_33_2 = result;
  end
  endfunction


  function automatic [5:0] MUX1HOT_v_6_3_2;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [2:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | ( input_1 & {6{sel[1]}});
    result = result | ( input_2 & {6{sel[2]}});
    MUX1HOT_v_6_3_2 = result;
  end
  endfunction


  function automatic [6:0] MUX1HOT_v_7_7_2;
    input [6:0] input_6;
    input [6:0] input_5;
    input [6:0] input_4;
    input [6:0] input_3;
    input [6:0] input_2;
    input [6:0] input_1;
    input [6:0] input_0;
    input [6:0] sel;
    reg [6:0] result;
  begin
    result = input_0 & {7{sel[0]}};
    result = result | ( input_1 & {7{sel[1]}});
    result = result | ( input_2 & {7{sel[2]}});
    result = result | ( input_3 & {7{sel[3]}});
    result = result | ( input_4 & {7{sel[4]}});
    result = result | ( input_5 & {7{sel[5]}});
    result = result | ( input_6 & {7{sel[6]}});
    MUX1HOT_v_7_7_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [9:0] MUX_v_10_2_2;
    input [9:0] input_0;
    input [9:0] input_1;
    input [0:0] sel;
    reg [9:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_10_2_2 = result;
  end
  endfunction


  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input [0:0] sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input [0:0] sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [0:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [54:0] MUX_v_55_2_2;
    input [54:0] input_0;
    input [54:0] input_1;
    input [0:0] sel;
    reg [54:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_55_2_2 = result;
  end
  endfunction


  function automatic [4:0] MUX_v_5_2_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input [0:0] sel;
    reg [4:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_5_2_2 = result;
  end
  endfunction


  function automatic [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function automatic [5:0] MUX_v_6_2_2;
    input [5:0] input_0;
    input [5:0] input_1;
    input [0:0] sel;
    reg [5:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_6_2_2 = result;
  end
  endfunction


  function automatic [11:0] readslicef_13_12_1;
    input [12:0] vector;
    reg [12:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_13_12_1 = tmp[11:0];
  end
  endfunction


  function automatic [63:0] readslicef_65_64_1;
    input [64:0] vector;
    reg [64:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_65_64_1 = tmp[63:0];
  end
  endfunction


  function automatic [64:0] readslicef_66_65_1;
    input [65:0] vector;
    reg [65:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_66_65_1 = tmp[64:0];
  end
  endfunction


  function automatic [0:0] readslicef_6_1_5;
    input [5:0] vector;
    reg [5:0] tmp;
  begin
    tmp = vector >> 5;
    readslicef_6_1_5 = tmp[0:0];
  end
  endfunction


  function automatic [12:0] conv_s2s_12_13 ;
    input [11:0]  vector ;
  begin
    conv_s2s_12_13 = {vector[11], vector};
  end
  endfunction


  function automatic [65:0] conv_s2u_65_66 ;
    input [64:0]  vector ;
  begin
    conv_s2u_65_66 = {vector[64], vector};
  end
  endfunction


  function automatic [12:0] conv_u2s_10_13 ;
    input [9:0]  vector ;
  begin
    conv_u2s_10_13 = {{3{1'b0}}, vector};
  end
  endfunction


  function automatic [6:0] conv_u2u_6_7 ;
    input [5:0]  vector ;
  begin
    conv_u2u_6_7 = {1'b0, vector};
  end
  endfunction


  function automatic [7:0] conv_u2u_7_8 ;
    input [6:0]  vector ;
  begin
    conv_u2u_7_8 = {1'b0, vector};
  end
  endfunction


  function automatic [8:0] conv_u2u_8_9 ;
    input [7:0]  vector ;
  begin
    conv_u2u_8_9 = {1'b0, vector};
  end
  endfunction


  function automatic [9:0] conv_u2u_9_10 ;
    input [8:0]  vector ;
  begin
    conv_u2u_9_10 = {1'b0, vector};
  end
  endfunction


  function automatic [10:0] conv_u2u_10_11 ;
    input [9:0]  vector ;
  begin
    conv_u2u_10_11 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF
// ------------------------------------------------------------------


module inPlaceNTT_DIF (
  clk, rst, vec_rsc_0_0_adra, vec_rsc_0_0_da, vec_rsc_0_0_wea, vec_rsc_0_0_qa, vec_rsc_triosy_0_0_lz,
      vec_rsc_0_1_adra, vec_rsc_0_1_da, vec_rsc_0_1_wea, vec_rsc_0_1_qa, vec_rsc_triosy_0_1_lz,
      vec_rsc_0_2_adra, vec_rsc_0_2_da, vec_rsc_0_2_wea, vec_rsc_0_2_qa, vec_rsc_triosy_0_2_lz,
      vec_rsc_0_3_adra, vec_rsc_0_3_da, vec_rsc_0_3_wea, vec_rsc_0_3_qa, vec_rsc_triosy_0_3_lz,
      vec_rsc_0_4_adra, vec_rsc_0_4_da, vec_rsc_0_4_wea, vec_rsc_0_4_qa, vec_rsc_triosy_0_4_lz,
      vec_rsc_0_5_adra, vec_rsc_0_5_da, vec_rsc_0_5_wea, vec_rsc_0_5_qa, vec_rsc_triosy_0_5_lz,
      vec_rsc_0_6_adra, vec_rsc_0_6_da, vec_rsc_0_6_wea, vec_rsc_0_6_qa, vec_rsc_triosy_0_6_lz,
      vec_rsc_0_7_adra, vec_rsc_0_7_da, vec_rsc_0_7_wea, vec_rsc_0_7_qa, vec_rsc_triosy_0_7_lz,
      vec_rsc_0_8_adra, vec_rsc_0_8_da, vec_rsc_0_8_wea, vec_rsc_0_8_qa, vec_rsc_triosy_0_8_lz,
      vec_rsc_0_9_adra, vec_rsc_0_9_da, vec_rsc_0_9_wea, vec_rsc_0_9_qa, vec_rsc_triosy_0_9_lz,
      vec_rsc_0_10_adra, vec_rsc_0_10_da, vec_rsc_0_10_wea, vec_rsc_0_10_qa, vec_rsc_triosy_0_10_lz,
      vec_rsc_0_11_adra, vec_rsc_0_11_da, vec_rsc_0_11_wea, vec_rsc_0_11_qa, vec_rsc_triosy_0_11_lz,
      vec_rsc_0_12_adra, vec_rsc_0_12_da, vec_rsc_0_12_wea, vec_rsc_0_12_qa, vec_rsc_triosy_0_12_lz,
      vec_rsc_0_13_adra, vec_rsc_0_13_da, vec_rsc_0_13_wea, vec_rsc_0_13_qa, vec_rsc_triosy_0_13_lz,
      vec_rsc_0_14_adra, vec_rsc_0_14_da, vec_rsc_0_14_wea, vec_rsc_0_14_qa, vec_rsc_triosy_0_14_lz,
      vec_rsc_0_15_adra, vec_rsc_0_15_da, vec_rsc_0_15_wea, vec_rsc_0_15_qa, vec_rsc_triosy_0_15_lz,
      p_rsc_dat, p_rsc_triosy_lz, r_rsc_dat, r_rsc_triosy_lz
);
  input clk;
  input rst;
  output [5:0] vec_rsc_0_0_adra;
  output [63:0] vec_rsc_0_0_da;
  output vec_rsc_0_0_wea;
  input [63:0] vec_rsc_0_0_qa;
  output vec_rsc_triosy_0_0_lz;
  output [5:0] vec_rsc_0_1_adra;
  output [63:0] vec_rsc_0_1_da;
  output vec_rsc_0_1_wea;
  input [63:0] vec_rsc_0_1_qa;
  output vec_rsc_triosy_0_1_lz;
  output [5:0] vec_rsc_0_2_adra;
  output [63:0] vec_rsc_0_2_da;
  output vec_rsc_0_2_wea;
  input [63:0] vec_rsc_0_2_qa;
  output vec_rsc_triosy_0_2_lz;
  output [5:0] vec_rsc_0_3_adra;
  output [63:0] vec_rsc_0_3_da;
  output vec_rsc_0_3_wea;
  input [63:0] vec_rsc_0_3_qa;
  output vec_rsc_triosy_0_3_lz;
  output [5:0] vec_rsc_0_4_adra;
  output [63:0] vec_rsc_0_4_da;
  output vec_rsc_0_4_wea;
  input [63:0] vec_rsc_0_4_qa;
  output vec_rsc_triosy_0_4_lz;
  output [5:0] vec_rsc_0_5_adra;
  output [63:0] vec_rsc_0_5_da;
  output vec_rsc_0_5_wea;
  input [63:0] vec_rsc_0_5_qa;
  output vec_rsc_triosy_0_5_lz;
  output [5:0] vec_rsc_0_6_adra;
  output [63:0] vec_rsc_0_6_da;
  output vec_rsc_0_6_wea;
  input [63:0] vec_rsc_0_6_qa;
  output vec_rsc_triosy_0_6_lz;
  output [5:0] vec_rsc_0_7_adra;
  output [63:0] vec_rsc_0_7_da;
  output vec_rsc_0_7_wea;
  input [63:0] vec_rsc_0_7_qa;
  output vec_rsc_triosy_0_7_lz;
  output [5:0] vec_rsc_0_8_adra;
  output [63:0] vec_rsc_0_8_da;
  output vec_rsc_0_8_wea;
  input [63:0] vec_rsc_0_8_qa;
  output vec_rsc_triosy_0_8_lz;
  output [5:0] vec_rsc_0_9_adra;
  output [63:0] vec_rsc_0_9_da;
  output vec_rsc_0_9_wea;
  input [63:0] vec_rsc_0_9_qa;
  output vec_rsc_triosy_0_9_lz;
  output [5:0] vec_rsc_0_10_adra;
  output [63:0] vec_rsc_0_10_da;
  output vec_rsc_0_10_wea;
  input [63:0] vec_rsc_0_10_qa;
  output vec_rsc_triosy_0_10_lz;
  output [5:0] vec_rsc_0_11_adra;
  output [63:0] vec_rsc_0_11_da;
  output vec_rsc_0_11_wea;
  input [63:0] vec_rsc_0_11_qa;
  output vec_rsc_triosy_0_11_lz;
  output [5:0] vec_rsc_0_12_adra;
  output [63:0] vec_rsc_0_12_da;
  output vec_rsc_0_12_wea;
  input [63:0] vec_rsc_0_12_qa;
  output vec_rsc_triosy_0_12_lz;
  output [5:0] vec_rsc_0_13_adra;
  output [63:0] vec_rsc_0_13_da;
  output vec_rsc_0_13_wea;
  input [63:0] vec_rsc_0_13_qa;
  output vec_rsc_triosy_0_13_lz;
  output [5:0] vec_rsc_0_14_adra;
  output [63:0] vec_rsc_0_14_da;
  output vec_rsc_0_14_wea;
  input [63:0] vec_rsc_0_14_qa;
  output vec_rsc_triosy_0_14_lz;
  output [5:0] vec_rsc_0_15_adra;
  output [63:0] vec_rsc_0_15_da;
  output vec_rsc_0_15_wea;
  input [63:0] vec_rsc_0_15_qa;
  output vec_rsc_triosy_0_15_lz;
  input [63:0] p_rsc_dat;
  output p_rsc_triosy_lz;
  input [63:0] r_rsc_dat;
  output r_rsc_triosy_lz;


  // Interconnect Declarations
  wire [63:0] vec_rsc_0_0_i_qa_d;
  wire vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_1_i_qa_d;
  wire vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_2_i_qa_d;
  wire vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_3_i_qa_d;
  wire vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_4_i_qa_d;
  wire vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_5_i_qa_d;
  wire vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_6_i_qa_d;
  wire vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_7_i_qa_d;
  wire vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_8_i_qa_d;
  wire vec_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_9_i_qa_d;
  wire vec_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_10_i_qa_d;
  wire vec_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_11_i_qa_d;
  wire vec_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_12_i_qa_d;
  wire vec_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_13_i_qa_d;
  wire vec_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_14_i_qa_d;
  wire vec_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_15_i_qa_d;
  wire vec_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [5:0] vec_rsc_0_0_i_adra_d_iff;
  wire [63:0] vec_rsc_0_0_i_da_d_iff;
  wire vec_rsc_0_0_i_wea_d_iff;
  wire vec_rsc_0_1_i_wea_d_iff;
  wire vec_rsc_0_2_i_wea_d_iff;
  wire vec_rsc_0_3_i_wea_d_iff;
  wire vec_rsc_0_4_i_wea_d_iff;
  wire vec_rsc_0_5_i_wea_d_iff;
  wire vec_rsc_0_6_i_wea_d_iff;
  wire vec_rsc_0_7_i_wea_d_iff;
  wire vec_rsc_0_8_i_wea_d_iff;
  wire vec_rsc_0_9_i_wea_d_iff;
  wire vec_rsc_0_10_i_wea_d_iff;
  wire vec_rsc_0_11_i_wea_d_iff;
  wire vec_rsc_0_12_i_wea_d_iff;
  wire vec_rsc_0_13_i_wea_d_iff;
  wire vec_rsc_0_14_i_wea_d_iff;
  wire vec_rsc_0_15_i_wea_d_iff;


  // Interconnect Declarations for Component Instantiations 
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_8_6_64_64_64_64_1_gen vec_rsc_0_0_i
      (
      .qa(vec_rsc_0_0_qa),
      .wea(vec_rsc_0_0_wea),
      .da(vec_rsc_0_0_da),
      .adra(vec_rsc_0_0_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_0_i_qa_d),
      .wea_d(vec_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_0_i_wea_d_iff)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_9_6_64_64_64_64_1_gen vec_rsc_0_1_i
      (
      .qa(vec_rsc_0_1_qa),
      .wea(vec_rsc_0_1_wea),
      .da(vec_rsc_0_1_da),
      .adra(vec_rsc_0_1_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_1_i_qa_d),
      .wea_d(vec_rsc_0_1_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_1_i_wea_d_iff)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_10_6_64_64_64_64_1_gen vec_rsc_0_2_i
      (
      .qa(vec_rsc_0_2_qa),
      .wea(vec_rsc_0_2_wea),
      .da(vec_rsc_0_2_da),
      .adra(vec_rsc_0_2_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_2_i_qa_d),
      .wea_d(vec_rsc_0_2_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_2_i_wea_d_iff)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_11_6_64_64_64_64_1_gen vec_rsc_0_3_i
      (
      .qa(vec_rsc_0_3_qa),
      .wea(vec_rsc_0_3_wea),
      .da(vec_rsc_0_3_da),
      .adra(vec_rsc_0_3_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_3_i_qa_d),
      .wea_d(vec_rsc_0_3_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_3_i_wea_d_iff)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_12_6_64_64_64_64_1_gen vec_rsc_0_4_i
      (
      .qa(vec_rsc_0_4_qa),
      .wea(vec_rsc_0_4_wea),
      .da(vec_rsc_0_4_da),
      .adra(vec_rsc_0_4_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_4_i_qa_d),
      .wea_d(vec_rsc_0_4_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_4_i_wea_d_iff)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_13_6_64_64_64_64_1_gen vec_rsc_0_5_i
      (
      .qa(vec_rsc_0_5_qa),
      .wea(vec_rsc_0_5_wea),
      .da(vec_rsc_0_5_da),
      .adra(vec_rsc_0_5_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_5_i_qa_d),
      .wea_d(vec_rsc_0_5_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_5_i_wea_d_iff)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_14_6_64_64_64_64_1_gen vec_rsc_0_6_i
      (
      .qa(vec_rsc_0_6_qa),
      .wea(vec_rsc_0_6_wea),
      .da(vec_rsc_0_6_da),
      .adra(vec_rsc_0_6_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_6_i_qa_d),
      .wea_d(vec_rsc_0_6_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_6_i_wea_d_iff)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_15_6_64_64_64_64_1_gen vec_rsc_0_7_i
      (
      .qa(vec_rsc_0_7_qa),
      .wea(vec_rsc_0_7_wea),
      .da(vec_rsc_0_7_da),
      .adra(vec_rsc_0_7_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_7_i_qa_d),
      .wea_d(vec_rsc_0_7_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_7_i_wea_d_iff)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_16_6_64_64_64_64_1_gen vec_rsc_0_8_i
      (
      .qa(vec_rsc_0_8_qa),
      .wea(vec_rsc_0_8_wea),
      .da(vec_rsc_0_8_da),
      .adra(vec_rsc_0_8_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_8_i_qa_d),
      .wea_d(vec_rsc_0_8_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_8_i_wea_d_iff)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_17_6_64_64_64_64_1_gen vec_rsc_0_9_i
      (
      .qa(vec_rsc_0_9_qa),
      .wea(vec_rsc_0_9_wea),
      .da(vec_rsc_0_9_da),
      .adra(vec_rsc_0_9_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_9_i_qa_d),
      .wea_d(vec_rsc_0_9_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_9_i_wea_d_iff)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_18_6_64_64_64_64_1_gen vec_rsc_0_10_i
      (
      .qa(vec_rsc_0_10_qa),
      .wea(vec_rsc_0_10_wea),
      .da(vec_rsc_0_10_da),
      .adra(vec_rsc_0_10_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_10_i_qa_d),
      .wea_d(vec_rsc_0_10_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_10_i_wea_d_iff)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_19_6_64_64_64_64_1_gen vec_rsc_0_11_i
      (
      .qa(vec_rsc_0_11_qa),
      .wea(vec_rsc_0_11_wea),
      .da(vec_rsc_0_11_da),
      .adra(vec_rsc_0_11_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_11_i_qa_d),
      .wea_d(vec_rsc_0_11_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_11_i_wea_d_iff)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_20_6_64_64_64_64_1_gen vec_rsc_0_12_i
      (
      .qa(vec_rsc_0_12_qa),
      .wea(vec_rsc_0_12_wea),
      .da(vec_rsc_0_12_da),
      .adra(vec_rsc_0_12_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_12_i_qa_d),
      .wea_d(vec_rsc_0_12_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_12_i_wea_d_iff)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_21_6_64_64_64_64_1_gen vec_rsc_0_13_i
      (
      .qa(vec_rsc_0_13_qa),
      .wea(vec_rsc_0_13_wea),
      .da(vec_rsc_0_13_da),
      .adra(vec_rsc_0_13_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_13_i_qa_d),
      .wea_d(vec_rsc_0_13_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_13_i_wea_d_iff)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_22_6_64_64_64_64_1_gen vec_rsc_0_14_i
      (
      .qa(vec_rsc_0_14_qa),
      .wea(vec_rsc_0_14_wea),
      .da(vec_rsc_0_14_da),
      .adra(vec_rsc_0_14_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_14_i_qa_d),
      .wea_d(vec_rsc_0_14_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_14_i_wea_d_iff)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_23_6_64_64_64_64_1_gen vec_rsc_0_15_i
      (
      .qa(vec_rsc_0_15_qa),
      .wea(vec_rsc_0_15_wea),
      .da(vec_rsc_0_15_da),
      .adra(vec_rsc_0_15_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_15_i_qa_d),
      .wea_d(vec_rsc_0_15_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_15_i_wea_d_iff)
    );
  inPlaceNTT_DIF_core inPlaceNTT_DIF_core_inst (
      .clk(clk),
      .rst(rst),
      .vec_rsc_triosy_0_0_lz(vec_rsc_triosy_0_0_lz),
      .vec_rsc_triosy_0_1_lz(vec_rsc_triosy_0_1_lz),
      .vec_rsc_triosy_0_2_lz(vec_rsc_triosy_0_2_lz),
      .vec_rsc_triosy_0_3_lz(vec_rsc_triosy_0_3_lz),
      .vec_rsc_triosy_0_4_lz(vec_rsc_triosy_0_4_lz),
      .vec_rsc_triosy_0_5_lz(vec_rsc_triosy_0_5_lz),
      .vec_rsc_triosy_0_6_lz(vec_rsc_triosy_0_6_lz),
      .vec_rsc_triosy_0_7_lz(vec_rsc_triosy_0_7_lz),
      .vec_rsc_triosy_0_8_lz(vec_rsc_triosy_0_8_lz),
      .vec_rsc_triosy_0_9_lz(vec_rsc_triosy_0_9_lz),
      .vec_rsc_triosy_0_10_lz(vec_rsc_triosy_0_10_lz),
      .vec_rsc_triosy_0_11_lz(vec_rsc_triosy_0_11_lz),
      .vec_rsc_triosy_0_12_lz(vec_rsc_triosy_0_12_lz),
      .vec_rsc_triosy_0_13_lz(vec_rsc_triosy_0_13_lz),
      .vec_rsc_triosy_0_14_lz(vec_rsc_triosy_0_14_lz),
      .vec_rsc_triosy_0_15_lz(vec_rsc_triosy_0_15_lz),
      .p_rsc_dat(p_rsc_dat),
      .p_rsc_triosy_lz(p_rsc_triosy_lz),
      .r_rsc_dat(r_rsc_dat),
      .r_rsc_triosy_lz(r_rsc_triosy_lz),
      .vec_rsc_0_0_i_qa_d(vec_rsc_0_0_i_qa_d),
      .vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_1_i_qa_d(vec_rsc_0_1_i_qa_d),
      .vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_2_i_qa_d(vec_rsc_0_2_i_qa_d),
      .vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_3_i_qa_d(vec_rsc_0_3_i_qa_d),
      .vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_4_i_qa_d(vec_rsc_0_4_i_qa_d),
      .vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_5_i_qa_d(vec_rsc_0_5_i_qa_d),
      .vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_6_i_qa_d(vec_rsc_0_6_i_qa_d),
      .vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_7_i_qa_d(vec_rsc_0_7_i_qa_d),
      .vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_8_i_qa_d(vec_rsc_0_8_i_qa_d),
      .vec_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_9_i_qa_d(vec_rsc_0_9_i_qa_d),
      .vec_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_10_i_qa_d(vec_rsc_0_10_i_qa_d),
      .vec_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_11_i_qa_d(vec_rsc_0_11_i_qa_d),
      .vec_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_12_i_qa_d(vec_rsc_0_12_i_qa_d),
      .vec_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_13_i_qa_d(vec_rsc_0_13_i_qa_d),
      .vec_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_14_i_qa_d(vec_rsc_0_14_i_qa_d),
      .vec_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_15_i_qa_d(vec_rsc_0_15_i_qa_d),
      .vec_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_0_i_adra_d_pff(vec_rsc_0_0_i_adra_d_iff),
      .vec_rsc_0_0_i_da_d_pff(vec_rsc_0_0_i_da_d_iff),
      .vec_rsc_0_0_i_wea_d_pff(vec_rsc_0_0_i_wea_d_iff),
      .vec_rsc_0_1_i_wea_d_pff(vec_rsc_0_1_i_wea_d_iff),
      .vec_rsc_0_2_i_wea_d_pff(vec_rsc_0_2_i_wea_d_iff),
      .vec_rsc_0_3_i_wea_d_pff(vec_rsc_0_3_i_wea_d_iff),
      .vec_rsc_0_4_i_wea_d_pff(vec_rsc_0_4_i_wea_d_iff),
      .vec_rsc_0_5_i_wea_d_pff(vec_rsc_0_5_i_wea_d_iff),
      .vec_rsc_0_6_i_wea_d_pff(vec_rsc_0_6_i_wea_d_iff),
      .vec_rsc_0_7_i_wea_d_pff(vec_rsc_0_7_i_wea_d_iff),
      .vec_rsc_0_8_i_wea_d_pff(vec_rsc_0_8_i_wea_d_iff),
      .vec_rsc_0_9_i_wea_d_pff(vec_rsc_0_9_i_wea_d_iff),
      .vec_rsc_0_10_i_wea_d_pff(vec_rsc_0_10_i_wea_d_iff),
      .vec_rsc_0_11_i_wea_d_pff(vec_rsc_0_11_i_wea_d_iff),
      .vec_rsc_0_12_i_wea_d_pff(vec_rsc_0_12_i_wea_d_iff),
      .vec_rsc_0_13_i_wea_d_pff(vec_rsc_0_13_i_wea_d_iff),
      .vec_rsc_0_14_i_wea_d_pff(vec_rsc_0_14_i_wea_d_iff),
      .vec_rsc_0_15_i_wea_d_pff(vec_rsc_0_15_i_wea_d_iff)
    );
endmodule



