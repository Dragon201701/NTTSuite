
//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_io_sync_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_io_sync_v2 (ld, lz);
    parameter valid = 0;

    input  ld;
    output lz;

    wire   lz;

    assign lz = ld;

endmodule


//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_rem_beh.v 
module mgc_rem(a,b,z);
   parameter width_a = 8;
   parameter width_b = 8;
   parameter signd = 1;
   input [width_a-1:0] a;
   input [width_b-1:0] b; 
   output [width_b-1:0] z;  
   reg  [width_b-1:0] z;

   always@(a or b)
     begin
	if(signd)
	  rem_s(a,b,z);
	else
          rem_u(a,b,z);
     end


//-----------------------------------------------------------------
//     -- Vectorized Overloaded Arithmetic Operators
//-----------------------------------------------------------------
   
   function [width_a-1:0] fabs_l; 
      input [width_a-1:0] arg1;
      begin
         case(arg1[width_a-1])
            1'b1:
               fabs_l = {(width_a){1'b0}} - arg1;
            default: // was: 1'b0:
               fabs_l = arg1;
         endcase
      end
   endfunction
   
   function [width_b-1:0] fabs_r; 
      input [width_b-1:0] arg1;
      begin
         case (arg1[width_b-1])
            1'b1:
               fabs_r =  {(width_b){1'b0}} - arg1;
            default: // was: 1'b0:
               fabs_r = arg1;
         endcase
      end
   endfunction

   function [width_b:0] minus;
     input [width_b:0] in1;
     input [width_b:0] in2;
     reg [width_b+1:0] tmp;
     begin
       tmp = in1 - in2;
       minus = tmp[width_b:0];
     end
   endfunction

   
   task divmod;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      output [width_b-1:0] rmod;
      
      parameter llen = width_a;
      parameter rlen = width_b;
      reg [(llen+rlen)-1:0] lbuf;
      reg [rlen:0] diff;
	  integer i;
      begin
	 lbuf = {(llen+rlen){1'b0}};
//64'b0;
	 lbuf[llen-1:0] = l;
	 for(i=width_a-1;i>=0;i=i-1)
	   begin
              diff = minus(lbuf[(llen+rlen)-1:llen-1], {1'b0,r});
	      rdiv[i] = ~diff[rlen];
	      if(diff[rlen] == 0)
		lbuf[(llen+rlen)-1:llen-1] = diff;
	      lbuf[(llen+rlen)-1:1] = lbuf[(llen+rlen)-2:0];
	   end
	 rmod = lbuf[(llen+rlen)-1:llen];
      end
   endtask
      

   task div_u;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(l, r, rdiv, rmod);
      end
   endtask
   
   task mod_u;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_b-1:0] rmod;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(l, r, rdiv, rmod);
      end
   endtask

   task rem_u; 
      input [width_a-1:0] l;
      input [width_b-1:0] r;    
      output [width_b-1:0] rmod;
      begin
	 mod_u(l,r,rmod);
      end
   endtask // rem_u

   task div_s;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(fabs_l(l), fabs_r(r),rdiv,rmod);
	 if(l[width_a-1] != r[width_b-1])
	   rdiv = {(width_a){1'b0}} - rdiv;
      end
   endtask

   task mod_s;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_b-1:0] rmod;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      reg [width_b-1:0] rnul;
      reg [width_b:0] rmod_t;
      begin
         rnul = {width_b{1'b0}};
	 divmod(fabs_l(l), fabs_r(r), rdiv, rmod);
         if (l[width_a-1])
	   rmod = {(width_b){1'b0}} - rmod;
	 if((rmod != rnul) && (l[width_a-1] != r[width_b-1]))
            begin
               rmod_t = r + rmod;
               rmod = rmod_t[width_b-1:0];
            end
      end
   endtask // mod_s
   
   task rem_s; 
      input [width_a-1:0] l;
      input [width_b-1:0] r;    
      output [width_b-1:0] rmod;   
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(fabs_l(l),fabs_r(r),rdiv,rmod);
	 if(l[width_a-1])
	   rmod = {(width_b){1'b0}} - rmod;
      end
   endtask

  endmodule

//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_div_beh.v 
module mgc_div(a,b,z);
   parameter width_a = 8;
   parameter width_b = 8;
   parameter signd = 1;
   input [width_a-1:0] a;
   input [width_b-1:0] b; 
   output [width_a-1:0] z;  
   reg  [width_a-1:0] z;

   always@(a or b)
     begin
	if(signd)
	  div_s(a,b,z);
	else
          div_u(a,b,z);
     end


//-----------------------------------------------------------------
//     -- Vectorized Overloaded Arithmetic Operators
//-----------------------------------------------------------------
   
   function [width_a-1:0] fabs_l; 
      input [width_a-1:0] arg1;
      begin
         case(arg1[width_a-1])
            1'b1:
               fabs_l = {(width_a){1'b0}} - arg1;
            default: // was: 1'b0:
               fabs_l = arg1;
         endcase
      end
   endfunction
   
   function [width_b-1:0] fabs_r; 
      input [width_b-1:0] arg1;
      begin
         case (arg1[width_b-1])
            1'b1:
               fabs_r =  {(width_b){1'b0}} - arg1;
            default: // was: 1'b0:
               fabs_r = arg1;
         endcase
      end
   endfunction

   function [width_b:0] minus;
     input [width_b:0] in1;
     input [width_b:0] in2;
     reg [width_b+1:0] tmp;
     begin
       tmp = in1 - in2;
       minus = tmp[width_b:0];
     end
   endfunction

   
   task divmod;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      output [width_b-1:0] rmod;
      
      parameter llen = width_a;
      parameter rlen = width_b;
      reg [(llen+rlen)-1:0] lbuf;
      reg [rlen:0] diff;
	  integer i;
      begin
	 lbuf = {(llen+rlen){1'b0}};
//64'b0;
	 lbuf[llen-1:0] = l;
	 for(i=width_a-1;i>=0;i=i-1)
	   begin
              diff = minus(lbuf[(llen+rlen)-1:llen-1], {1'b0,r});
	      rdiv[i] = ~diff[rlen];
	      if(diff[rlen] == 0)
		lbuf[(llen+rlen)-1:llen-1] = diff;
	      lbuf[(llen+rlen)-1:1] = lbuf[(llen+rlen)-2:0];
	   end
	 rmod = lbuf[(llen+rlen)-1:llen];
      end
   endtask
      

   task div_u;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(l, r, rdiv, rmod);
      end
   endtask
   
   task mod_u;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_b-1:0] rmod;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(l, r, rdiv, rmod);
      end
   endtask

   task rem_u; 
      input [width_a-1:0] l;
      input [width_b-1:0] r;    
      output [width_b-1:0] rmod;
      begin
	 mod_u(l,r,rmod);
      end
   endtask // rem_u

   task div_s;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(fabs_l(l), fabs_r(r),rdiv,rmod);
	 if(l[width_a-1] != r[width_b-1])
	   rdiv = {(width_a){1'b0}} - rdiv;
      end
   endtask

   task mod_s;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_b-1:0] rmod;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      reg [width_b-1:0] rnul;
      reg [width_b:0] rmod_t;
      begin
         rnul = {width_b{1'b0}};
	 divmod(fabs_l(l), fabs_r(r), rdiv, rmod);
         if (l[width_a-1])
	   rmod = {(width_b){1'b0}} - rmod;
	 if((rmod != rnul) && (l[width_a-1] != r[width_b-1]))
            begin
               rmod_t = r + rmod;
               rmod = rmod_t[width_b-1:0];
            end
      end
   endtask // mod_s
   
   task rem_s; 
      input [width_a-1:0] l;
      input [width_b-1:0] r;    
      output [width_b-1:0] rmod;   
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(fabs_l(l),fabs_r(r),rdiv,rmod);
	 if(l[width_a-1])
	   rmod = {(width_b){1'b0}} - rmod;
      end
   endtask

  endmodule

//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_shift_l_beh_v5.v 
module mgc_shift_l_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
   if (signd_a)
   begin: SGNED
      assign z = fshl_u(a,s,a[width_a-1]);
   end
   else
   begin: UNSGNED
      assign z = fshl_u(a,s,1'b0);
   end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u

endmodule

//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5c/896140 Production Release
//  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
// 
//  Generated by:   yl7897@newnano.poly.edu
//  Generated date: Thu Jul  1 00:57:50 2021
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_19_8_64_256_256_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_19_8_64_256_256_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [7:0] adra;
  input [7:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_18_8_64_256_256_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_18_8_64_256_256_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [7:0] adra;
  input [7:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_17_8_64_256_256_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_17_8_64_256_256_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [7:0] adra;
  input [7:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_16_8_64_256_256_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_16_8_64_256_256_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [7:0] adra;
  input [7:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_15_8_64_256_256_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_15_8_64_256_256_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [7:0] adra;
  input [7:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_14_8_64_256_256_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_14_8_64_256_256_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [7:0] adra;
  input [7:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_13_8_64_256_256_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_13_8_64_256_256_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [7:0] adra;
  input [7:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_12_8_64_256_256_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_12_8_64_256_256_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [7:0] adra;
  input [7:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_11_8_64_256_256_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_11_8_64_256_256_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [7:0] adra;
  input [7:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_10_8_64_256_256_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_10_8_64_256_256_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [7:0] adra;
  input [7:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_9_8_64_256_256_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_9_8_64_256_256_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [7:0] adra;
  input [7:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_8_8_64_256_256_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_8_8_64_256_256_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [7:0] adra;
  input [7:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_7_8_64_256_256_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_7_8_64_256_256_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [7:0] adra;
  input [7:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_6_8_64_256_256_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_6_8_64_256_256_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [7:0] adra;
  input [7:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_5_8_64_256_256_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_5_8_64_256_256_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [7:0] adra;
  input [7:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_4_8_64_256_256_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_4_8_64_256_256_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [7:0] adra;
  input [7:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module inPlaceNTT_DIT_core_core_fsm (
  clk, rst, fsm_output, STAGE_LOOP_C_8_tr0, modExp_while_C_38_tr0, COMP_LOOP_C_1_tr0,
      COMP_LOOP_1_modExp_1_while_C_38_tr0, COMP_LOOP_C_62_tr0, COMP_LOOP_2_modExp_1_while_C_38_tr0,
      COMP_LOOP_C_124_tr0, COMP_LOOP_3_modExp_1_while_C_38_tr0, COMP_LOOP_C_186_tr0,
      COMP_LOOP_4_modExp_1_while_C_38_tr0, COMP_LOOP_C_248_tr0, COMP_LOOP_5_modExp_1_while_C_38_tr0,
      COMP_LOOP_C_310_tr0, COMP_LOOP_6_modExp_1_while_C_38_tr0, COMP_LOOP_C_372_tr0,
      COMP_LOOP_7_modExp_1_while_C_38_tr0, COMP_LOOP_C_434_tr0, COMP_LOOP_8_modExp_1_while_C_38_tr0,
      COMP_LOOP_C_496_tr0, COMP_LOOP_9_modExp_1_while_C_38_tr0, COMP_LOOP_C_558_tr0,
      COMP_LOOP_10_modExp_1_while_C_38_tr0, COMP_LOOP_C_620_tr0, COMP_LOOP_11_modExp_1_while_C_38_tr0,
      COMP_LOOP_C_682_tr0, COMP_LOOP_12_modExp_1_while_C_38_tr0, COMP_LOOP_C_744_tr0,
      COMP_LOOP_13_modExp_1_while_C_38_tr0, COMP_LOOP_C_806_tr0, COMP_LOOP_14_modExp_1_while_C_38_tr0,
      COMP_LOOP_C_868_tr0, COMP_LOOP_15_modExp_1_while_C_38_tr0, COMP_LOOP_C_930_tr0,
      COMP_LOOP_16_modExp_1_while_C_38_tr0, COMP_LOOP_C_992_tr0, VEC_LOOP_C_0_tr0,
      STAGE_LOOP_C_9_tr0
);
  input clk;
  input rst;
  output [10:0] fsm_output;
  reg [10:0] fsm_output;
  input STAGE_LOOP_C_8_tr0;
  input modExp_while_C_38_tr0;
  input COMP_LOOP_C_1_tr0;
  input COMP_LOOP_1_modExp_1_while_C_38_tr0;
  input COMP_LOOP_C_62_tr0;
  input COMP_LOOP_2_modExp_1_while_C_38_tr0;
  input COMP_LOOP_C_124_tr0;
  input COMP_LOOP_3_modExp_1_while_C_38_tr0;
  input COMP_LOOP_C_186_tr0;
  input COMP_LOOP_4_modExp_1_while_C_38_tr0;
  input COMP_LOOP_C_248_tr0;
  input COMP_LOOP_5_modExp_1_while_C_38_tr0;
  input COMP_LOOP_C_310_tr0;
  input COMP_LOOP_6_modExp_1_while_C_38_tr0;
  input COMP_LOOP_C_372_tr0;
  input COMP_LOOP_7_modExp_1_while_C_38_tr0;
  input COMP_LOOP_C_434_tr0;
  input COMP_LOOP_8_modExp_1_while_C_38_tr0;
  input COMP_LOOP_C_496_tr0;
  input COMP_LOOP_9_modExp_1_while_C_38_tr0;
  input COMP_LOOP_C_558_tr0;
  input COMP_LOOP_10_modExp_1_while_C_38_tr0;
  input COMP_LOOP_C_620_tr0;
  input COMP_LOOP_11_modExp_1_while_C_38_tr0;
  input COMP_LOOP_C_682_tr0;
  input COMP_LOOP_12_modExp_1_while_C_38_tr0;
  input COMP_LOOP_C_744_tr0;
  input COMP_LOOP_13_modExp_1_while_C_38_tr0;
  input COMP_LOOP_C_806_tr0;
  input COMP_LOOP_14_modExp_1_while_C_38_tr0;
  input COMP_LOOP_C_868_tr0;
  input COMP_LOOP_15_modExp_1_while_C_38_tr0;
  input COMP_LOOP_C_930_tr0;
  input COMP_LOOP_16_modExp_1_while_C_38_tr0;
  input COMP_LOOP_C_992_tr0;
  input VEC_LOOP_C_0_tr0;
  input STAGE_LOOP_C_9_tr0;


  // FSM State Type Declaration for inPlaceNTT_DIT_core_core_fsm_1
  parameter
    main_C_0 = 11'd0,
    STAGE_LOOP_C_0 = 11'd1,
    STAGE_LOOP_C_1 = 11'd2,
    STAGE_LOOP_C_2 = 11'd3,
    STAGE_LOOP_C_3 = 11'd4,
    STAGE_LOOP_C_4 = 11'd5,
    STAGE_LOOP_C_5 = 11'd6,
    STAGE_LOOP_C_6 = 11'd7,
    STAGE_LOOP_C_7 = 11'd8,
    STAGE_LOOP_C_8 = 11'd9,
    modExp_while_C_0 = 11'd10,
    modExp_while_C_1 = 11'd11,
    modExp_while_C_2 = 11'd12,
    modExp_while_C_3 = 11'd13,
    modExp_while_C_4 = 11'd14,
    modExp_while_C_5 = 11'd15,
    modExp_while_C_6 = 11'd16,
    modExp_while_C_7 = 11'd17,
    modExp_while_C_8 = 11'd18,
    modExp_while_C_9 = 11'd19,
    modExp_while_C_10 = 11'd20,
    modExp_while_C_11 = 11'd21,
    modExp_while_C_12 = 11'd22,
    modExp_while_C_13 = 11'd23,
    modExp_while_C_14 = 11'd24,
    modExp_while_C_15 = 11'd25,
    modExp_while_C_16 = 11'd26,
    modExp_while_C_17 = 11'd27,
    modExp_while_C_18 = 11'd28,
    modExp_while_C_19 = 11'd29,
    modExp_while_C_20 = 11'd30,
    modExp_while_C_21 = 11'd31,
    modExp_while_C_22 = 11'd32,
    modExp_while_C_23 = 11'd33,
    modExp_while_C_24 = 11'd34,
    modExp_while_C_25 = 11'd35,
    modExp_while_C_26 = 11'd36,
    modExp_while_C_27 = 11'd37,
    modExp_while_C_28 = 11'd38,
    modExp_while_C_29 = 11'd39,
    modExp_while_C_30 = 11'd40,
    modExp_while_C_31 = 11'd41,
    modExp_while_C_32 = 11'd42,
    modExp_while_C_33 = 11'd43,
    modExp_while_C_34 = 11'd44,
    modExp_while_C_35 = 11'd45,
    modExp_while_C_36 = 11'd46,
    modExp_while_C_37 = 11'd47,
    modExp_while_C_38 = 11'd48,
    COMP_LOOP_C_0 = 11'd49,
    COMP_LOOP_C_1 = 11'd50,
    COMP_LOOP_1_modExp_1_while_C_0 = 11'd51,
    COMP_LOOP_1_modExp_1_while_C_1 = 11'd52,
    COMP_LOOP_1_modExp_1_while_C_2 = 11'd53,
    COMP_LOOP_1_modExp_1_while_C_3 = 11'd54,
    COMP_LOOP_1_modExp_1_while_C_4 = 11'd55,
    COMP_LOOP_1_modExp_1_while_C_5 = 11'd56,
    COMP_LOOP_1_modExp_1_while_C_6 = 11'd57,
    COMP_LOOP_1_modExp_1_while_C_7 = 11'd58,
    COMP_LOOP_1_modExp_1_while_C_8 = 11'd59,
    COMP_LOOP_1_modExp_1_while_C_9 = 11'd60,
    COMP_LOOP_1_modExp_1_while_C_10 = 11'd61,
    COMP_LOOP_1_modExp_1_while_C_11 = 11'd62,
    COMP_LOOP_1_modExp_1_while_C_12 = 11'd63,
    COMP_LOOP_1_modExp_1_while_C_13 = 11'd64,
    COMP_LOOP_1_modExp_1_while_C_14 = 11'd65,
    COMP_LOOP_1_modExp_1_while_C_15 = 11'd66,
    COMP_LOOP_1_modExp_1_while_C_16 = 11'd67,
    COMP_LOOP_1_modExp_1_while_C_17 = 11'd68,
    COMP_LOOP_1_modExp_1_while_C_18 = 11'd69,
    COMP_LOOP_1_modExp_1_while_C_19 = 11'd70,
    COMP_LOOP_1_modExp_1_while_C_20 = 11'd71,
    COMP_LOOP_1_modExp_1_while_C_21 = 11'd72,
    COMP_LOOP_1_modExp_1_while_C_22 = 11'd73,
    COMP_LOOP_1_modExp_1_while_C_23 = 11'd74,
    COMP_LOOP_1_modExp_1_while_C_24 = 11'd75,
    COMP_LOOP_1_modExp_1_while_C_25 = 11'd76,
    COMP_LOOP_1_modExp_1_while_C_26 = 11'd77,
    COMP_LOOP_1_modExp_1_while_C_27 = 11'd78,
    COMP_LOOP_1_modExp_1_while_C_28 = 11'd79,
    COMP_LOOP_1_modExp_1_while_C_29 = 11'd80,
    COMP_LOOP_1_modExp_1_while_C_30 = 11'd81,
    COMP_LOOP_1_modExp_1_while_C_31 = 11'd82,
    COMP_LOOP_1_modExp_1_while_C_32 = 11'd83,
    COMP_LOOP_1_modExp_1_while_C_33 = 11'd84,
    COMP_LOOP_1_modExp_1_while_C_34 = 11'd85,
    COMP_LOOP_1_modExp_1_while_C_35 = 11'd86,
    COMP_LOOP_1_modExp_1_while_C_36 = 11'd87,
    COMP_LOOP_1_modExp_1_while_C_37 = 11'd88,
    COMP_LOOP_1_modExp_1_while_C_38 = 11'd89,
    COMP_LOOP_C_2 = 11'd90,
    COMP_LOOP_C_3 = 11'd91,
    COMP_LOOP_C_4 = 11'd92,
    COMP_LOOP_C_5 = 11'd93,
    COMP_LOOP_C_6 = 11'd94,
    COMP_LOOP_C_7 = 11'd95,
    COMP_LOOP_C_8 = 11'd96,
    COMP_LOOP_C_9 = 11'd97,
    COMP_LOOP_C_10 = 11'd98,
    COMP_LOOP_C_11 = 11'd99,
    COMP_LOOP_C_12 = 11'd100,
    COMP_LOOP_C_13 = 11'd101,
    COMP_LOOP_C_14 = 11'd102,
    COMP_LOOP_C_15 = 11'd103,
    COMP_LOOP_C_16 = 11'd104,
    COMP_LOOP_C_17 = 11'd105,
    COMP_LOOP_C_18 = 11'd106,
    COMP_LOOP_C_19 = 11'd107,
    COMP_LOOP_C_20 = 11'd108,
    COMP_LOOP_C_21 = 11'd109,
    COMP_LOOP_C_22 = 11'd110,
    COMP_LOOP_C_23 = 11'd111,
    COMP_LOOP_C_24 = 11'd112,
    COMP_LOOP_C_25 = 11'd113,
    COMP_LOOP_C_26 = 11'd114,
    COMP_LOOP_C_27 = 11'd115,
    COMP_LOOP_C_28 = 11'd116,
    COMP_LOOP_C_29 = 11'd117,
    COMP_LOOP_C_30 = 11'd118,
    COMP_LOOP_C_31 = 11'd119,
    COMP_LOOP_C_32 = 11'd120,
    COMP_LOOP_C_33 = 11'd121,
    COMP_LOOP_C_34 = 11'd122,
    COMP_LOOP_C_35 = 11'd123,
    COMP_LOOP_C_36 = 11'd124,
    COMP_LOOP_C_37 = 11'd125,
    COMP_LOOP_C_38 = 11'd126,
    COMP_LOOP_C_39 = 11'd127,
    COMP_LOOP_C_40 = 11'd128,
    COMP_LOOP_C_41 = 11'd129,
    COMP_LOOP_C_42 = 11'd130,
    COMP_LOOP_C_43 = 11'd131,
    COMP_LOOP_C_44 = 11'd132,
    COMP_LOOP_C_45 = 11'd133,
    COMP_LOOP_C_46 = 11'd134,
    COMP_LOOP_C_47 = 11'd135,
    COMP_LOOP_C_48 = 11'd136,
    COMP_LOOP_C_49 = 11'd137,
    COMP_LOOP_C_50 = 11'd138,
    COMP_LOOP_C_51 = 11'd139,
    COMP_LOOP_C_52 = 11'd140,
    COMP_LOOP_C_53 = 11'd141,
    COMP_LOOP_C_54 = 11'd142,
    COMP_LOOP_C_55 = 11'd143,
    COMP_LOOP_C_56 = 11'd144,
    COMP_LOOP_C_57 = 11'd145,
    COMP_LOOP_C_58 = 11'd146,
    COMP_LOOP_C_59 = 11'd147,
    COMP_LOOP_C_60 = 11'd148,
    COMP_LOOP_C_61 = 11'd149,
    COMP_LOOP_C_62 = 11'd150,
    COMP_LOOP_C_63 = 11'd151,
    COMP_LOOP_2_modExp_1_while_C_0 = 11'd152,
    COMP_LOOP_2_modExp_1_while_C_1 = 11'd153,
    COMP_LOOP_2_modExp_1_while_C_2 = 11'd154,
    COMP_LOOP_2_modExp_1_while_C_3 = 11'd155,
    COMP_LOOP_2_modExp_1_while_C_4 = 11'd156,
    COMP_LOOP_2_modExp_1_while_C_5 = 11'd157,
    COMP_LOOP_2_modExp_1_while_C_6 = 11'd158,
    COMP_LOOP_2_modExp_1_while_C_7 = 11'd159,
    COMP_LOOP_2_modExp_1_while_C_8 = 11'd160,
    COMP_LOOP_2_modExp_1_while_C_9 = 11'd161,
    COMP_LOOP_2_modExp_1_while_C_10 = 11'd162,
    COMP_LOOP_2_modExp_1_while_C_11 = 11'd163,
    COMP_LOOP_2_modExp_1_while_C_12 = 11'd164,
    COMP_LOOP_2_modExp_1_while_C_13 = 11'd165,
    COMP_LOOP_2_modExp_1_while_C_14 = 11'd166,
    COMP_LOOP_2_modExp_1_while_C_15 = 11'd167,
    COMP_LOOP_2_modExp_1_while_C_16 = 11'd168,
    COMP_LOOP_2_modExp_1_while_C_17 = 11'd169,
    COMP_LOOP_2_modExp_1_while_C_18 = 11'd170,
    COMP_LOOP_2_modExp_1_while_C_19 = 11'd171,
    COMP_LOOP_2_modExp_1_while_C_20 = 11'd172,
    COMP_LOOP_2_modExp_1_while_C_21 = 11'd173,
    COMP_LOOP_2_modExp_1_while_C_22 = 11'd174,
    COMP_LOOP_2_modExp_1_while_C_23 = 11'd175,
    COMP_LOOP_2_modExp_1_while_C_24 = 11'd176,
    COMP_LOOP_2_modExp_1_while_C_25 = 11'd177,
    COMP_LOOP_2_modExp_1_while_C_26 = 11'd178,
    COMP_LOOP_2_modExp_1_while_C_27 = 11'd179,
    COMP_LOOP_2_modExp_1_while_C_28 = 11'd180,
    COMP_LOOP_2_modExp_1_while_C_29 = 11'd181,
    COMP_LOOP_2_modExp_1_while_C_30 = 11'd182,
    COMP_LOOP_2_modExp_1_while_C_31 = 11'd183,
    COMP_LOOP_2_modExp_1_while_C_32 = 11'd184,
    COMP_LOOP_2_modExp_1_while_C_33 = 11'd185,
    COMP_LOOP_2_modExp_1_while_C_34 = 11'd186,
    COMP_LOOP_2_modExp_1_while_C_35 = 11'd187,
    COMP_LOOP_2_modExp_1_while_C_36 = 11'd188,
    COMP_LOOP_2_modExp_1_while_C_37 = 11'd189,
    COMP_LOOP_2_modExp_1_while_C_38 = 11'd190,
    COMP_LOOP_C_64 = 11'd191,
    COMP_LOOP_C_65 = 11'd192,
    COMP_LOOP_C_66 = 11'd193,
    COMP_LOOP_C_67 = 11'd194,
    COMP_LOOP_C_68 = 11'd195,
    COMP_LOOP_C_69 = 11'd196,
    COMP_LOOP_C_70 = 11'd197,
    COMP_LOOP_C_71 = 11'd198,
    COMP_LOOP_C_72 = 11'd199,
    COMP_LOOP_C_73 = 11'd200,
    COMP_LOOP_C_74 = 11'd201,
    COMP_LOOP_C_75 = 11'd202,
    COMP_LOOP_C_76 = 11'd203,
    COMP_LOOP_C_77 = 11'd204,
    COMP_LOOP_C_78 = 11'd205,
    COMP_LOOP_C_79 = 11'd206,
    COMP_LOOP_C_80 = 11'd207,
    COMP_LOOP_C_81 = 11'd208,
    COMP_LOOP_C_82 = 11'd209,
    COMP_LOOP_C_83 = 11'd210,
    COMP_LOOP_C_84 = 11'd211,
    COMP_LOOP_C_85 = 11'd212,
    COMP_LOOP_C_86 = 11'd213,
    COMP_LOOP_C_87 = 11'd214,
    COMP_LOOP_C_88 = 11'd215,
    COMP_LOOP_C_89 = 11'd216,
    COMP_LOOP_C_90 = 11'd217,
    COMP_LOOP_C_91 = 11'd218,
    COMP_LOOP_C_92 = 11'd219,
    COMP_LOOP_C_93 = 11'd220,
    COMP_LOOP_C_94 = 11'd221,
    COMP_LOOP_C_95 = 11'd222,
    COMP_LOOP_C_96 = 11'd223,
    COMP_LOOP_C_97 = 11'd224,
    COMP_LOOP_C_98 = 11'd225,
    COMP_LOOP_C_99 = 11'd226,
    COMP_LOOP_C_100 = 11'd227,
    COMP_LOOP_C_101 = 11'd228,
    COMP_LOOP_C_102 = 11'd229,
    COMP_LOOP_C_103 = 11'd230,
    COMP_LOOP_C_104 = 11'd231,
    COMP_LOOP_C_105 = 11'd232,
    COMP_LOOP_C_106 = 11'd233,
    COMP_LOOP_C_107 = 11'd234,
    COMP_LOOP_C_108 = 11'd235,
    COMP_LOOP_C_109 = 11'd236,
    COMP_LOOP_C_110 = 11'd237,
    COMP_LOOP_C_111 = 11'd238,
    COMP_LOOP_C_112 = 11'd239,
    COMP_LOOP_C_113 = 11'd240,
    COMP_LOOP_C_114 = 11'd241,
    COMP_LOOP_C_115 = 11'd242,
    COMP_LOOP_C_116 = 11'd243,
    COMP_LOOP_C_117 = 11'd244,
    COMP_LOOP_C_118 = 11'd245,
    COMP_LOOP_C_119 = 11'd246,
    COMP_LOOP_C_120 = 11'd247,
    COMP_LOOP_C_121 = 11'd248,
    COMP_LOOP_C_122 = 11'd249,
    COMP_LOOP_C_123 = 11'd250,
    COMP_LOOP_C_124 = 11'd251,
    COMP_LOOP_C_125 = 11'd252,
    COMP_LOOP_3_modExp_1_while_C_0 = 11'd253,
    COMP_LOOP_3_modExp_1_while_C_1 = 11'd254,
    COMP_LOOP_3_modExp_1_while_C_2 = 11'd255,
    COMP_LOOP_3_modExp_1_while_C_3 = 11'd256,
    COMP_LOOP_3_modExp_1_while_C_4 = 11'd257,
    COMP_LOOP_3_modExp_1_while_C_5 = 11'd258,
    COMP_LOOP_3_modExp_1_while_C_6 = 11'd259,
    COMP_LOOP_3_modExp_1_while_C_7 = 11'd260,
    COMP_LOOP_3_modExp_1_while_C_8 = 11'd261,
    COMP_LOOP_3_modExp_1_while_C_9 = 11'd262,
    COMP_LOOP_3_modExp_1_while_C_10 = 11'd263,
    COMP_LOOP_3_modExp_1_while_C_11 = 11'd264,
    COMP_LOOP_3_modExp_1_while_C_12 = 11'd265,
    COMP_LOOP_3_modExp_1_while_C_13 = 11'd266,
    COMP_LOOP_3_modExp_1_while_C_14 = 11'd267,
    COMP_LOOP_3_modExp_1_while_C_15 = 11'd268,
    COMP_LOOP_3_modExp_1_while_C_16 = 11'd269,
    COMP_LOOP_3_modExp_1_while_C_17 = 11'd270,
    COMP_LOOP_3_modExp_1_while_C_18 = 11'd271,
    COMP_LOOP_3_modExp_1_while_C_19 = 11'd272,
    COMP_LOOP_3_modExp_1_while_C_20 = 11'd273,
    COMP_LOOP_3_modExp_1_while_C_21 = 11'd274,
    COMP_LOOP_3_modExp_1_while_C_22 = 11'd275,
    COMP_LOOP_3_modExp_1_while_C_23 = 11'd276,
    COMP_LOOP_3_modExp_1_while_C_24 = 11'd277,
    COMP_LOOP_3_modExp_1_while_C_25 = 11'd278,
    COMP_LOOP_3_modExp_1_while_C_26 = 11'd279,
    COMP_LOOP_3_modExp_1_while_C_27 = 11'd280,
    COMP_LOOP_3_modExp_1_while_C_28 = 11'd281,
    COMP_LOOP_3_modExp_1_while_C_29 = 11'd282,
    COMP_LOOP_3_modExp_1_while_C_30 = 11'd283,
    COMP_LOOP_3_modExp_1_while_C_31 = 11'd284,
    COMP_LOOP_3_modExp_1_while_C_32 = 11'd285,
    COMP_LOOP_3_modExp_1_while_C_33 = 11'd286,
    COMP_LOOP_3_modExp_1_while_C_34 = 11'd287,
    COMP_LOOP_3_modExp_1_while_C_35 = 11'd288,
    COMP_LOOP_3_modExp_1_while_C_36 = 11'd289,
    COMP_LOOP_3_modExp_1_while_C_37 = 11'd290,
    COMP_LOOP_3_modExp_1_while_C_38 = 11'd291,
    COMP_LOOP_C_126 = 11'd292,
    COMP_LOOP_C_127 = 11'd293,
    COMP_LOOP_C_128 = 11'd294,
    COMP_LOOP_C_129 = 11'd295,
    COMP_LOOP_C_130 = 11'd296,
    COMP_LOOP_C_131 = 11'd297,
    COMP_LOOP_C_132 = 11'd298,
    COMP_LOOP_C_133 = 11'd299,
    COMP_LOOP_C_134 = 11'd300,
    COMP_LOOP_C_135 = 11'd301,
    COMP_LOOP_C_136 = 11'd302,
    COMP_LOOP_C_137 = 11'd303,
    COMP_LOOP_C_138 = 11'd304,
    COMP_LOOP_C_139 = 11'd305,
    COMP_LOOP_C_140 = 11'd306,
    COMP_LOOP_C_141 = 11'd307,
    COMP_LOOP_C_142 = 11'd308,
    COMP_LOOP_C_143 = 11'd309,
    COMP_LOOP_C_144 = 11'd310,
    COMP_LOOP_C_145 = 11'd311,
    COMP_LOOP_C_146 = 11'd312,
    COMP_LOOP_C_147 = 11'd313,
    COMP_LOOP_C_148 = 11'd314,
    COMP_LOOP_C_149 = 11'd315,
    COMP_LOOP_C_150 = 11'd316,
    COMP_LOOP_C_151 = 11'd317,
    COMP_LOOP_C_152 = 11'd318,
    COMP_LOOP_C_153 = 11'd319,
    COMP_LOOP_C_154 = 11'd320,
    COMP_LOOP_C_155 = 11'd321,
    COMP_LOOP_C_156 = 11'd322,
    COMP_LOOP_C_157 = 11'd323,
    COMP_LOOP_C_158 = 11'd324,
    COMP_LOOP_C_159 = 11'd325,
    COMP_LOOP_C_160 = 11'd326,
    COMP_LOOP_C_161 = 11'd327,
    COMP_LOOP_C_162 = 11'd328,
    COMP_LOOP_C_163 = 11'd329,
    COMP_LOOP_C_164 = 11'd330,
    COMP_LOOP_C_165 = 11'd331,
    COMP_LOOP_C_166 = 11'd332,
    COMP_LOOP_C_167 = 11'd333,
    COMP_LOOP_C_168 = 11'd334,
    COMP_LOOP_C_169 = 11'd335,
    COMP_LOOP_C_170 = 11'd336,
    COMP_LOOP_C_171 = 11'd337,
    COMP_LOOP_C_172 = 11'd338,
    COMP_LOOP_C_173 = 11'd339,
    COMP_LOOP_C_174 = 11'd340,
    COMP_LOOP_C_175 = 11'd341,
    COMP_LOOP_C_176 = 11'd342,
    COMP_LOOP_C_177 = 11'd343,
    COMP_LOOP_C_178 = 11'd344,
    COMP_LOOP_C_179 = 11'd345,
    COMP_LOOP_C_180 = 11'd346,
    COMP_LOOP_C_181 = 11'd347,
    COMP_LOOP_C_182 = 11'd348,
    COMP_LOOP_C_183 = 11'd349,
    COMP_LOOP_C_184 = 11'd350,
    COMP_LOOP_C_185 = 11'd351,
    COMP_LOOP_C_186 = 11'd352,
    COMP_LOOP_C_187 = 11'd353,
    COMP_LOOP_4_modExp_1_while_C_0 = 11'd354,
    COMP_LOOP_4_modExp_1_while_C_1 = 11'd355,
    COMP_LOOP_4_modExp_1_while_C_2 = 11'd356,
    COMP_LOOP_4_modExp_1_while_C_3 = 11'd357,
    COMP_LOOP_4_modExp_1_while_C_4 = 11'd358,
    COMP_LOOP_4_modExp_1_while_C_5 = 11'd359,
    COMP_LOOP_4_modExp_1_while_C_6 = 11'd360,
    COMP_LOOP_4_modExp_1_while_C_7 = 11'd361,
    COMP_LOOP_4_modExp_1_while_C_8 = 11'd362,
    COMP_LOOP_4_modExp_1_while_C_9 = 11'd363,
    COMP_LOOP_4_modExp_1_while_C_10 = 11'd364,
    COMP_LOOP_4_modExp_1_while_C_11 = 11'd365,
    COMP_LOOP_4_modExp_1_while_C_12 = 11'd366,
    COMP_LOOP_4_modExp_1_while_C_13 = 11'd367,
    COMP_LOOP_4_modExp_1_while_C_14 = 11'd368,
    COMP_LOOP_4_modExp_1_while_C_15 = 11'd369,
    COMP_LOOP_4_modExp_1_while_C_16 = 11'd370,
    COMP_LOOP_4_modExp_1_while_C_17 = 11'd371,
    COMP_LOOP_4_modExp_1_while_C_18 = 11'd372,
    COMP_LOOP_4_modExp_1_while_C_19 = 11'd373,
    COMP_LOOP_4_modExp_1_while_C_20 = 11'd374,
    COMP_LOOP_4_modExp_1_while_C_21 = 11'd375,
    COMP_LOOP_4_modExp_1_while_C_22 = 11'd376,
    COMP_LOOP_4_modExp_1_while_C_23 = 11'd377,
    COMP_LOOP_4_modExp_1_while_C_24 = 11'd378,
    COMP_LOOP_4_modExp_1_while_C_25 = 11'd379,
    COMP_LOOP_4_modExp_1_while_C_26 = 11'd380,
    COMP_LOOP_4_modExp_1_while_C_27 = 11'd381,
    COMP_LOOP_4_modExp_1_while_C_28 = 11'd382,
    COMP_LOOP_4_modExp_1_while_C_29 = 11'd383,
    COMP_LOOP_4_modExp_1_while_C_30 = 11'd384,
    COMP_LOOP_4_modExp_1_while_C_31 = 11'd385,
    COMP_LOOP_4_modExp_1_while_C_32 = 11'd386,
    COMP_LOOP_4_modExp_1_while_C_33 = 11'd387,
    COMP_LOOP_4_modExp_1_while_C_34 = 11'd388,
    COMP_LOOP_4_modExp_1_while_C_35 = 11'd389,
    COMP_LOOP_4_modExp_1_while_C_36 = 11'd390,
    COMP_LOOP_4_modExp_1_while_C_37 = 11'd391,
    COMP_LOOP_4_modExp_1_while_C_38 = 11'd392,
    COMP_LOOP_C_188 = 11'd393,
    COMP_LOOP_C_189 = 11'd394,
    COMP_LOOP_C_190 = 11'd395,
    COMP_LOOP_C_191 = 11'd396,
    COMP_LOOP_C_192 = 11'd397,
    COMP_LOOP_C_193 = 11'd398,
    COMP_LOOP_C_194 = 11'd399,
    COMP_LOOP_C_195 = 11'd400,
    COMP_LOOP_C_196 = 11'd401,
    COMP_LOOP_C_197 = 11'd402,
    COMP_LOOP_C_198 = 11'd403,
    COMP_LOOP_C_199 = 11'd404,
    COMP_LOOP_C_200 = 11'd405,
    COMP_LOOP_C_201 = 11'd406,
    COMP_LOOP_C_202 = 11'd407,
    COMP_LOOP_C_203 = 11'd408,
    COMP_LOOP_C_204 = 11'd409,
    COMP_LOOP_C_205 = 11'd410,
    COMP_LOOP_C_206 = 11'd411,
    COMP_LOOP_C_207 = 11'd412,
    COMP_LOOP_C_208 = 11'd413,
    COMP_LOOP_C_209 = 11'd414,
    COMP_LOOP_C_210 = 11'd415,
    COMP_LOOP_C_211 = 11'd416,
    COMP_LOOP_C_212 = 11'd417,
    COMP_LOOP_C_213 = 11'd418,
    COMP_LOOP_C_214 = 11'd419,
    COMP_LOOP_C_215 = 11'd420,
    COMP_LOOP_C_216 = 11'd421,
    COMP_LOOP_C_217 = 11'd422,
    COMP_LOOP_C_218 = 11'd423,
    COMP_LOOP_C_219 = 11'd424,
    COMP_LOOP_C_220 = 11'd425,
    COMP_LOOP_C_221 = 11'd426,
    COMP_LOOP_C_222 = 11'd427,
    COMP_LOOP_C_223 = 11'd428,
    COMP_LOOP_C_224 = 11'd429,
    COMP_LOOP_C_225 = 11'd430,
    COMP_LOOP_C_226 = 11'd431,
    COMP_LOOP_C_227 = 11'd432,
    COMP_LOOP_C_228 = 11'd433,
    COMP_LOOP_C_229 = 11'd434,
    COMP_LOOP_C_230 = 11'd435,
    COMP_LOOP_C_231 = 11'd436,
    COMP_LOOP_C_232 = 11'd437,
    COMP_LOOP_C_233 = 11'd438,
    COMP_LOOP_C_234 = 11'd439,
    COMP_LOOP_C_235 = 11'd440,
    COMP_LOOP_C_236 = 11'd441,
    COMP_LOOP_C_237 = 11'd442,
    COMP_LOOP_C_238 = 11'd443,
    COMP_LOOP_C_239 = 11'd444,
    COMP_LOOP_C_240 = 11'd445,
    COMP_LOOP_C_241 = 11'd446,
    COMP_LOOP_C_242 = 11'd447,
    COMP_LOOP_C_243 = 11'd448,
    COMP_LOOP_C_244 = 11'd449,
    COMP_LOOP_C_245 = 11'd450,
    COMP_LOOP_C_246 = 11'd451,
    COMP_LOOP_C_247 = 11'd452,
    COMP_LOOP_C_248 = 11'd453,
    COMP_LOOP_C_249 = 11'd454,
    COMP_LOOP_5_modExp_1_while_C_0 = 11'd455,
    COMP_LOOP_5_modExp_1_while_C_1 = 11'd456,
    COMP_LOOP_5_modExp_1_while_C_2 = 11'd457,
    COMP_LOOP_5_modExp_1_while_C_3 = 11'd458,
    COMP_LOOP_5_modExp_1_while_C_4 = 11'd459,
    COMP_LOOP_5_modExp_1_while_C_5 = 11'd460,
    COMP_LOOP_5_modExp_1_while_C_6 = 11'd461,
    COMP_LOOP_5_modExp_1_while_C_7 = 11'd462,
    COMP_LOOP_5_modExp_1_while_C_8 = 11'd463,
    COMP_LOOP_5_modExp_1_while_C_9 = 11'd464,
    COMP_LOOP_5_modExp_1_while_C_10 = 11'd465,
    COMP_LOOP_5_modExp_1_while_C_11 = 11'd466,
    COMP_LOOP_5_modExp_1_while_C_12 = 11'd467,
    COMP_LOOP_5_modExp_1_while_C_13 = 11'd468,
    COMP_LOOP_5_modExp_1_while_C_14 = 11'd469,
    COMP_LOOP_5_modExp_1_while_C_15 = 11'd470,
    COMP_LOOP_5_modExp_1_while_C_16 = 11'd471,
    COMP_LOOP_5_modExp_1_while_C_17 = 11'd472,
    COMP_LOOP_5_modExp_1_while_C_18 = 11'd473,
    COMP_LOOP_5_modExp_1_while_C_19 = 11'd474,
    COMP_LOOP_5_modExp_1_while_C_20 = 11'd475,
    COMP_LOOP_5_modExp_1_while_C_21 = 11'd476,
    COMP_LOOP_5_modExp_1_while_C_22 = 11'd477,
    COMP_LOOP_5_modExp_1_while_C_23 = 11'd478,
    COMP_LOOP_5_modExp_1_while_C_24 = 11'd479,
    COMP_LOOP_5_modExp_1_while_C_25 = 11'd480,
    COMP_LOOP_5_modExp_1_while_C_26 = 11'd481,
    COMP_LOOP_5_modExp_1_while_C_27 = 11'd482,
    COMP_LOOP_5_modExp_1_while_C_28 = 11'd483,
    COMP_LOOP_5_modExp_1_while_C_29 = 11'd484,
    COMP_LOOP_5_modExp_1_while_C_30 = 11'd485,
    COMP_LOOP_5_modExp_1_while_C_31 = 11'd486,
    COMP_LOOP_5_modExp_1_while_C_32 = 11'd487,
    COMP_LOOP_5_modExp_1_while_C_33 = 11'd488,
    COMP_LOOP_5_modExp_1_while_C_34 = 11'd489,
    COMP_LOOP_5_modExp_1_while_C_35 = 11'd490,
    COMP_LOOP_5_modExp_1_while_C_36 = 11'd491,
    COMP_LOOP_5_modExp_1_while_C_37 = 11'd492,
    COMP_LOOP_5_modExp_1_while_C_38 = 11'd493,
    COMP_LOOP_C_250 = 11'd494,
    COMP_LOOP_C_251 = 11'd495,
    COMP_LOOP_C_252 = 11'd496,
    COMP_LOOP_C_253 = 11'd497,
    COMP_LOOP_C_254 = 11'd498,
    COMP_LOOP_C_255 = 11'd499,
    COMP_LOOP_C_256 = 11'd500,
    COMP_LOOP_C_257 = 11'd501,
    COMP_LOOP_C_258 = 11'd502,
    COMP_LOOP_C_259 = 11'd503,
    COMP_LOOP_C_260 = 11'd504,
    COMP_LOOP_C_261 = 11'd505,
    COMP_LOOP_C_262 = 11'd506,
    COMP_LOOP_C_263 = 11'd507,
    COMP_LOOP_C_264 = 11'd508,
    COMP_LOOP_C_265 = 11'd509,
    COMP_LOOP_C_266 = 11'd510,
    COMP_LOOP_C_267 = 11'd511,
    COMP_LOOP_C_268 = 11'd512,
    COMP_LOOP_C_269 = 11'd513,
    COMP_LOOP_C_270 = 11'd514,
    COMP_LOOP_C_271 = 11'd515,
    COMP_LOOP_C_272 = 11'd516,
    COMP_LOOP_C_273 = 11'd517,
    COMP_LOOP_C_274 = 11'd518,
    COMP_LOOP_C_275 = 11'd519,
    COMP_LOOP_C_276 = 11'd520,
    COMP_LOOP_C_277 = 11'd521,
    COMP_LOOP_C_278 = 11'd522,
    COMP_LOOP_C_279 = 11'd523,
    COMP_LOOP_C_280 = 11'd524,
    COMP_LOOP_C_281 = 11'd525,
    COMP_LOOP_C_282 = 11'd526,
    COMP_LOOP_C_283 = 11'd527,
    COMP_LOOP_C_284 = 11'd528,
    COMP_LOOP_C_285 = 11'd529,
    COMP_LOOP_C_286 = 11'd530,
    COMP_LOOP_C_287 = 11'd531,
    COMP_LOOP_C_288 = 11'd532,
    COMP_LOOP_C_289 = 11'd533,
    COMP_LOOP_C_290 = 11'd534,
    COMP_LOOP_C_291 = 11'd535,
    COMP_LOOP_C_292 = 11'd536,
    COMP_LOOP_C_293 = 11'd537,
    COMP_LOOP_C_294 = 11'd538,
    COMP_LOOP_C_295 = 11'd539,
    COMP_LOOP_C_296 = 11'd540,
    COMP_LOOP_C_297 = 11'd541,
    COMP_LOOP_C_298 = 11'd542,
    COMP_LOOP_C_299 = 11'd543,
    COMP_LOOP_C_300 = 11'd544,
    COMP_LOOP_C_301 = 11'd545,
    COMP_LOOP_C_302 = 11'd546,
    COMP_LOOP_C_303 = 11'd547,
    COMP_LOOP_C_304 = 11'd548,
    COMP_LOOP_C_305 = 11'd549,
    COMP_LOOP_C_306 = 11'd550,
    COMP_LOOP_C_307 = 11'd551,
    COMP_LOOP_C_308 = 11'd552,
    COMP_LOOP_C_309 = 11'd553,
    COMP_LOOP_C_310 = 11'd554,
    COMP_LOOP_C_311 = 11'd555,
    COMP_LOOP_6_modExp_1_while_C_0 = 11'd556,
    COMP_LOOP_6_modExp_1_while_C_1 = 11'd557,
    COMP_LOOP_6_modExp_1_while_C_2 = 11'd558,
    COMP_LOOP_6_modExp_1_while_C_3 = 11'd559,
    COMP_LOOP_6_modExp_1_while_C_4 = 11'd560,
    COMP_LOOP_6_modExp_1_while_C_5 = 11'd561,
    COMP_LOOP_6_modExp_1_while_C_6 = 11'd562,
    COMP_LOOP_6_modExp_1_while_C_7 = 11'd563,
    COMP_LOOP_6_modExp_1_while_C_8 = 11'd564,
    COMP_LOOP_6_modExp_1_while_C_9 = 11'd565,
    COMP_LOOP_6_modExp_1_while_C_10 = 11'd566,
    COMP_LOOP_6_modExp_1_while_C_11 = 11'd567,
    COMP_LOOP_6_modExp_1_while_C_12 = 11'd568,
    COMP_LOOP_6_modExp_1_while_C_13 = 11'd569,
    COMP_LOOP_6_modExp_1_while_C_14 = 11'd570,
    COMP_LOOP_6_modExp_1_while_C_15 = 11'd571,
    COMP_LOOP_6_modExp_1_while_C_16 = 11'd572,
    COMP_LOOP_6_modExp_1_while_C_17 = 11'd573,
    COMP_LOOP_6_modExp_1_while_C_18 = 11'd574,
    COMP_LOOP_6_modExp_1_while_C_19 = 11'd575,
    COMP_LOOP_6_modExp_1_while_C_20 = 11'd576,
    COMP_LOOP_6_modExp_1_while_C_21 = 11'd577,
    COMP_LOOP_6_modExp_1_while_C_22 = 11'd578,
    COMP_LOOP_6_modExp_1_while_C_23 = 11'd579,
    COMP_LOOP_6_modExp_1_while_C_24 = 11'd580,
    COMP_LOOP_6_modExp_1_while_C_25 = 11'd581,
    COMP_LOOP_6_modExp_1_while_C_26 = 11'd582,
    COMP_LOOP_6_modExp_1_while_C_27 = 11'd583,
    COMP_LOOP_6_modExp_1_while_C_28 = 11'd584,
    COMP_LOOP_6_modExp_1_while_C_29 = 11'd585,
    COMP_LOOP_6_modExp_1_while_C_30 = 11'd586,
    COMP_LOOP_6_modExp_1_while_C_31 = 11'd587,
    COMP_LOOP_6_modExp_1_while_C_32 = 11'd588,
    COMP_LOOP_6_modExp_1_while_C_33 = 11'd589,
    COMP_LOOP_6_modExp_1_while_C_34 = 11'd590,
    COMP_LOOP_6_modExp_1_while_C_35 = 11'd591,
    COMP_LOOP_6_modExp_1_while_C_36 = 11'd592,
    COMP_LOOP_6_modExp_1_while_C_37 = 11'd593,
    COMP_LOOP_6_modExp_1_while_C_38 = 11'd594,
    COMP_LOOP_C_312 = 11'd595,
    COMP_LOOP_C_313 = 11'd596,
    COMP_LOOP_C_314 = 11'd597,
    COMP_LOOP_C_315 = 11'd598,
    COMP_LOOP_C_316 = 11'd599,
    COMP_LOOP_C_317 = 11'd600,
    COMP_LOOP_C_318 = 11'd601,
    COMP_LOOP_C_319 = 11'd602,
    COMP_LOOP_C_320 = 11'd603,
    COMP_LOOP_C_321 = 11'd604,
    COMP_LOOP_C_322 = 11'd605,
    COMP_LOOP_C_323 = 11'd606,
    COMP_LOOP_C_324 = 11'd607,
    COMP_LOOP_C_325 = 11'd608,
    COMP_LOOP_C_326 = 11'd609,
    COMP_LOOP_C_327 = 11'd610,
    COMP_LOOP_C_328 = 11'd611,
    COMP_LOOP_C_329 = 11'd612,
    COMP_LOOP_C_330 = 11'd613,
    COMP_LOOP_C_331 = 11'd614,
    COMP_LOOP_C_332 = 11'd615,
    COMP_LOOP_C_333 = 11'd616,
    COMP_LOOP_C_334 = 11'd617,
    COMP_LOOP_C_335 = 11'd618,
    COMP_LOOP_C_336 = 11'd619,
    COMP_LOOP_C_337 = 11'd620,
    COMP_LOOP_C_338 = 11'd621,
    COMP_LOOP_C_339 = 11'd622,
    COMP_LOOP_C_340 = 11'd623,
    COMP_LOOP_C_341 = 11'd624,
    COMP_LOOP_C_342 = 11'd625,
    COMP_LOOP_C_343 = 11'd626,
    COMP_LOOP_C_344 = 11'd627,
    COMP_LOOP_C_345 = 11'd628,
    COMP_LOOP_C_346 = 11'd629,
    COMP_LOOP_C_347 = 11'd630,
    COMP_LOOP_C_348 = 11'd631,
    COMP_LOOP_C_349 = 11'd632,
    COMP_LOOP_C_350 = 11'd633,
    COMP_LOOP_C_351 = 11'd634,
    COMP_LOOP_C_352 = 11'd635,
    COMP_LOOP_C_353 = 11'd636,
    COMP_LOOP_C_354 = 11'd637,
    COMP_LOOP_C_355 = 11'd638,
    COMP_LOOP_C_356 = 11'd639,
    COMP_LOOP_C_357 = 11'd640,
    COMP_LOOP_C_358 = 11'd641,
    COMP_LOOP_C_359 = 11'd642,
    COMP_LOOP_C_360 = 11'd643,
    COMP_LOOP_C_361 = 11'd644,
    COMP_LOOP_C_362 = 11'd645,
    COMP_LOOP_C_363 = 11'd646,
    COMP_LOOP_C_364 = 11'd647,
    COMP_LOOP_C_365 = 11'd648,
    COMP_LOOP_C_366 = 11'd649,
    COMP_LOOP_C_367 = 11'd650,
    COMP_LOOP_C_368 = 11'd651,
    COMP_LOOP_C_369 = 11'd652,
    COMP_LOOP_C_370 = 11'd653,
    COMP_LOOP_C_371 = 11'd654,
    COMP_LOOP_C_372 = 11'd655,
    COMP_LOOP_C_373 = 11'd656,
    COMP_LOOP_7_modExp_1_while_C_0 = 11'd657,
    COMP_LOOP_7_modExp_1_while_C_1 = 11'd658,
    COMP_LOOP_7_modExp_1_while_C_2 = 11'd659,
    COMP_LOOP_7_modExp_1_while_C_3 = 11'd660,
    COMP_LOOP_7_modExp_1_while_C_4 = 11'd661,
    COMP_LOOP_7_modExp_1_while_C_5 = 11'd662,
    COMP_LOOP_7_modExp_1_while_C_6 = 11'd663,
    COMP_LOOP_7_modExp_1_while_C_7 = 11'd664,
    COMP_LOOP_7_modExp_1_while_C_8 = 11'd665,
    COMP_LOOP_7_modExp_1_while_C_9 = 11'd666,
    COMP_LOOP_7_modExp_1_while_C_10 = 11'd667,
    COMP_LOOP_7_modExp_1_while_C_11 = 11'd668,
    COMP_LOOP_7_modExp_1_while_C_12 = 11'd669,
    COMP_LOOP_7_modExp_1_while_C_13 = 11'd670,
    COMP_LOOP_7_modExp_1_while_C_14 = 11'd671,
    COMP_LOOP_7_modExp_1_while_C_15 = 11'd672,
    COMP_LOOP_7_modExp_1_while_C_16 = 11'd673,
    COMP_LOOP_7_modExp_1_while_C_17 = 11'd674,
    COMP_LOOP_7_modExp_1_while_C_18 = 11'd675,
    COMP_LOOP_7_modExp_1_while_C_19 = 11'd676,
    COMP_LOOP_7_modExp_1_while_C_20 = 11'd677,
    COMP_LOOP_7_modExp_1_while_C_21 = 11'd678,
    COMP_LOOP_7_modExp_1_while_C_22 = 11'd679,
    COMP_LOOP_7_modExp_1_while_C_23 = 11'd680,
    COMP_LOOP_7_modExp_1_while_C_24 = 11'd681,
    COMP_LOOP_7_modExp_1_while_C_25 = 11'd682,
    COMP_LOOP_7_modExp_1_while_C_26 = 11'd683,
    COMP_LOOP_7_modExp_1_while_C_27 = 11'd684,
    COMP_LOOP_7_modExp_1_while_C_28 = 11'd685,
    COMP_LOOP_7_modExp_1_while_C_29 = 11'd686,
    COMP_LOOP_7_modExp_1_while_C_30 = 11'd687,
    COMP_LOOP_7_modExp_1_while_C_31 = 11'd688,
    COMP_LOOP_7_modExp_1_while_C_32 = 11'd689,
    COMP_LOOP_7_modExp_1_while_C_33 = 11'd690,
    COMP_LOOP_7_modExp_1_while_C_34 = 11'd691,
    COMP_LOOP_7_modExp_1_while_C_35 = 11'd692,
    COMP_LOOP_7_modExp_1_while_C_36 = 11'd693,
    COMP_LOOP_7_modExp_1_while_C_37 = 11'd694,
    COMP_LOOP_7_modExp_1_while_C_38 = 11'd695,
    COMP_LOOP_C_374 = 11'd696,
    COMP_LOOP_C_375 = 11'd697,
    COMP_LOOP_C_376 = 11'd698,
    COMP_LOOP_C_377 = 11'd699,
    COMP_LOOP_C_378 = 11'd700,
    COMP_LOOP_C_379 = 11'd701,
    COMP_LOOP_C_380 = 11'd702,
    COMP_LOOP_C_381 = 11'd703,
    COMP_LOOP_C_382 = 11'd704,
    COMP_LOOP_C_383 = 11'd705,
    COMP_LOOP_C_384 = 11'd706,
    COMP_LOOP_C_385 = 11'd707,
    COMP_LOOP_C_386 = 11'd708,
    COMP_LOOP_C_387 = 11'd709,
    COMP_LOOP_C_388 = 11'd710,
    COMP_LOOP_C_389 = 11'd711,
    COMP_LOOP_C_390 = 11'd712,
    COMP_LOOP_C_391 = 11'd713,
    COMP_LOOP_C_392 = 11'd714,
    COMP_LOOP_C_393 = 11'd715,
    COMP_LOOP_C_394 = 11'd716,
    COMP_LOOP_C_395 = 11'd717,
    COMP_LOOP_C_396 = 11'd718,
    COMP_LOOP_C_397 = 11'd719,
    COMP_LOOP_C_398 = 11'd720,
    COMP_LOOP_C_399 = 11'd721,
    COMP_LOOP_C_400 = 11'd722,
    COMP_LOOP_C_401 = 11'd723,
    COMP_LOOP_C_402 = 11'd724,
    COMP_LOOP_C_403 = 11'd725,
    COMP_LOOP_C_404 = 11'd726,
    COMP_LOOP_C_405 = 11'd727,
    COMP_LOOP_C_406 = 11'd728,
    COMP_LOOP_C_407 = 11'd729,
    COMP_LOOP_C_408 = 11'd730,
    COMP_LOOP_C_409 = 11'd731,
    COMP_LOOP_C_410 = 11'd732,
    COMP_LOOP_C_411 = 11'd733,
    COMP_LOOP_C_412 = 11'd734,
    COMP_LOOP_C_413 = 11'd735,
    COMP_LOOP_C_414 = 11'd736,
    COMP_LOOP_C_415 = 11'd737,
    COMP_LOOP_C_416 = 11'd738,
    COMP_LOOP_C_417 = 11'd739,
    COMP_LOOP_C_418 = 11'd740,
    COMP_LOOP_C_419 = 11'd741,
    COMP_LOOP_C_420 = 11'd742,
    COMP_LOOP_C_421 = 11'd743,
    COMP_LOOP_C_422 = 11'd744,
    COMP_LOOP_C_423 = 11'd745,
    COMP_LOOP_C_424 = 11'd746,
    COMP_LOOP_C_425 = 11'd747,
    COMP_LOOP_C_426 = 11'd748,
    COMP_LOOP_C_427 = 11'd749,
    COMP_LOOP_C_428 = 11'd750,
    COMP_LOOP_C_429 = 11'd751,
    COMP_LOOP_C_430 = 11'd752,
    COMP_LOOP_C_431 = 11'd753,
    COMP_LOOP_C_432 = 11'd754,
    COMP_LOOP_C_433 = 11'd755,
    COMP_LOOP_C_434 = 11'd756,
    COMP_LOOP_C_435 = 11'd757,
    COMP_LOOP_8_modExp_1_while_C_0 = 11'd758,
    COMP_LOOP_8_modExp_1_while_C_1 = 11'd759,
    COMP_LOOP_8_modExp_1_while_C_2 = 11'd760,
    COMP_LOOP_8_modExp_1_while_C_3 = 11'd761,
    COMP_LOOP_8_modExp_1_while_C_4 = 11'd762,
    COMP_LOOP_8_modExp_1_while_C_5 = 11'd763,
    COMP_LOOP_8_modExp_1_while_C_6 = 11'd764,
    COMP_LOOP_8_modExp_1_while_C_7 = 11'd765,
    COMP_LOOP_8_modExp_1_while_C_8 = 11'd766,
    COMP_LOOP_8_modExp_1_while_C_9 = 11'd767,
    COMP_LOOP_8_modExp_1_while_C_10 = 11'd768,
    COMP_LOOP_8_modExp_1_while_C_11 = 11'd769,
    COMP_LOOP_8_modExp_1_while_C_12 = 11'd770,
    COMP_LOOP_8_modExp_1_while_C_13 = 11'd771,
    COMP_LOOP_8_modExp_1_while_C_14 = 11'd772,
    COMP_LOOP_8_modExp_1_while_C_15 = 11'd773,
    COMP_LOOP_8_modExp_1_while_C_16 = 11'd774,
    COMP_LOOP_8_modExp_1_while_C_17 = 11'd775,
    COMP_LOOP_8_modExp_1_while_C_18 = 11'd776,
    COMP_LOOP_8_modExp_1_while_C_19 = 11'd777,
    COMP_LOOP_8_modExp_1_while_C_20 = 11'd778,
    COMP_LOOP_8_modExp_1_while_C_21 = 11'd779,
    COMP_LOOP_8_modExp_1_while_C_22 = 11'd780,
    COMP_LOOP_8_modExp_1_while_C_23 = 11'd781,
    COMP_LOOP_8_modExp_1_while_C_24 = 11'd782,
    COMP_LOOP_8_modExp_1_while_C_25 = 11'd783,
    COMP_LOOP_8_modExp_1_while_C_26 = 11'd784,
    COMP_LOOP_8_modExp_1_while_C_27 = 11'd785,
    COMP_LOOP_8_modExp_1_while_C_28 = 11'd786,
    COMP_LOOP_8_modExp_1_while_C_29 = 11'd787,
    COMP_LOOP_8_modExp_1_while_C_30 = 11'd788,
    COMP_LOOP_8_modExp_1_while_C_31 = 11'd789,
    COMP_LOOP_8_modExp_1_while_C_32 = 11'd790,
    COMP_LOOP_8_modExp_1_while_C_33 = 11'd791,
    COMP_LOOP_8_modExp_1_while_C_34 = 11'd792,
    COMP_LOOP_8_modExp_1_while_C_35 = 11'd793,
    COMP_LOOP_8_modExp_1_while_C_36 = 11'd794,
    COMP_LOOP_8_modExp_1_while_C_37 = 11'd795,
    COMP_LOOP_8_modExp_1_while_C_38 = 11'd796,
    COMP_LOOP_C_436 = 11'd797,
    COMP_LOOP_C_437 = 11'd798,
    COMP_LOOP_C_438 = 11'd799,
    COMP_LOOP_C_439 = 11'd800,
    COMP_LOOP_C_440 = 11'd801,
    COMP_LOOP_C_441 = 11'd802,
    COMP_LOOP_C_442 = 11'd803,
    COMP_LOOP_C_443 = 11'd804,
    COMP_LOOP_C_444 = 11'd805,
    COMP_LOOP_C_445 = 11'd806,
    COMP_LOOP_C_446 = 11'd807,
    COMP_LOOP_C_447 = 11'd808,
    COMP_LOOP_C_448 = 11'd809,
    COMP_LOOP_C_449 = 11'd810,
    COMP_LOOP_C_450 = 11'd811,
    COMP_LOOP_C_451 = 11'd812,
    COMP_LOOP_C_452 = 11'd813,
    COMP_LOOP_C_453 = 11'd814,
    COMP_LOOP_C_454 = 11'd815,
    COMP_LOOP_C_455 = 11'd816,
    COMP_LOOP_C_456 = 11'd817,
    COMP_LOOP_C_457 = 11'd818,
    COMP_LOOP_C_458 = 11'd819,
    COMP_LOOP_C_459 = 11'd820,
    COMP_LOOP_C_460 = 11'd821,
    COMP_LOOP_C_461 = 11'd822,
    COMP_LOOP_C_462 = 11'd823,
    COMP_LOOP_C_463 = 11'd824,
    COMP_LOOP_C_464 = 11'd825,
    COMP_LOOP_C_465 = 11'd826,
    COMP_LOOP_C_466 = 11'd827,
    COMP_LOOP_C_467 = 11'd828,
    COMP_LOOP_C_468 = 11'd829,
    COMP_LOOP_C_469 = 11'd830,
    COMP_LOOP_C_470 = 11'd831,
    COMP_LOOP_C_471 = 11'd832,
    COMP_LOOP_C_472 = 11'd833,
    COMP_LOOP_C_473 = 11'd834,
    COMP_LOOP_C_474 = 11'd835,
    COMP_LOOP_C_475 = 11'd836,
    COMP_LOOP_C_476 = 11'd837,
    COMP_LOOP_C_477 = 11'd838,
    COMP_LOOP_C_478 = 11'd839,
    COMP_LOOP_C_479 = 11'd840,
    COMP_LOOP_C_480 = 11'd841,
    COMP_LOOP_C_481 = 11'd842,
    COMP_LOOP_C_482 = 11'd843,
    COMP_LOOP_C_483 = 11'd844,
    COMP_LOOP_C_484 = 11'd845,
    COMP_LOOP_C_485 = 11'd846,
    COMP_LOOP_C_486 = 11'd847,
    COMP_LOOP_C_487 = 11'd848,
    COMP_LOOP_C_488 = 11'd849,
    COMP_LOOP_C_489 = 11'd850,
    COMP_LOOP_C_490 = 11'd851,
    COMP_LOOP_C_491 = 11'd852,
    COMP_LOOP_C_492 = 11'd853,
    COMP_LOOP_C_493 = 11'd854,
    COMP_LOOP_C_494 = 11'd855,
    COMP_LOOP_C_495 = 11'd856,
    COMP_LOOP_C_496 = 11'd857,
    COMP_LOOP_C_497 = 11'd858,
    COMP_LOOP_9_modExp_1_while_C_0 = 11'd859,
    COMP_LOOP_9_modExp_1_while_C_1 = 11'd860,
    COMP_LOOP_9_modExp_1_while_C_2 = 11'd861,
    COMP_LOOP_9_modExp_1_while_C_3 = 11'd862,
    COMP_LOOP_9_modExp_1_while_C_4 = 11'd863,
    COMP_LOOP_9_modExp_1_while_C_5 = 11'd864,
    COMP_LOOP_9_modExp_1_while_C_6 = 11'd865,
    COMP_LOOP_9_modExp_1_while_C_7 = 11'd866,
    COMP_LOOP_9_modExp_1_while_C_8 = 11'd867,
    COMP_LOOP_9_modExp_1_while_C_9 = 11'd868,
    COMP_LOOP_9_modExp_1_while_C_10 = 11'd869,
    COMP_LOOP_9_modExp_1_while_C_11 = 11'd870,
    COMP_LOOP_9_modExp_1_while_C_12 = 11'd871,
    COMP_LOOP_9_modExp_1_while_C_13 = 11'd872,
    COMP_LOOP_9_modExp_1_while_C_14 = 11'd873,
    COMP_LOOP_9_modExp_1_while_C_15 = 11'd874,
    COMP_LOOP_9_modExp_1_while_C_16 = 11'd875,
    COMP_LOOP_9_modExp_1_while_C_17 = 11'd876,
    COMP_LOOP_9_modExp_1_while_C_18 = 11'd877,
    COMP_LOOP_9_modExp_1_while_C_19 = 11'd878,
    COMP_LOOP_9_modExp_1_while_C_20 = 11'd879,
    COMP_LOOP_9_modExp_1_while_C_21 = 11'd880,
    COMP_LOOP_9_modExp_1_while_C_22 = 11'd881,
    COMP_LOOP_9_modExp_1_while_C_23 = 11'd882,
    COMP_LOOP_9_modExp_1_while_C_24 = 11'd883,
    COMP_LOOP_9_modExp_1_while_C_25 = 11'd884,
    COMP_LOOP_9_modExp_1_while_C_26 = 11'd885,
    COMP_LOOP_9_modExp_1_while_C_27 = 11'd886,
    COMP_LOOP_9_modExp_1_while_C_28 = 11'd887,
    COMP_LOOP_9_modExp_1_while_C_29 = 11'd888,
    COMP_LOOP_9_modExp_1_while_C_30 = 11'd889,
    COMP_LOOP_9_modExp_1_while_C_31 = 11'd890,
    COMP_LOOP_9_modExp_1_while_C_32 = 11'd891,
    COMP_LOOP_9_modExp_1_while_C_33 = 11'd892,
    COMP_LOOP_9_modExp_1_while_C_34 = 11'd893,
    COMP_LOOP_9_modExp_1_while_C_35 = 11'd894,
    COMP_LOOP_9_modExp_1_while_C_36 = 11'd895,
    COMP_LOOP_9_modExp_1_while_C_37 = 11'd896,
    COMP_LOOP_9_modExp_1_while_C_38 = 11'd897,
    COMP_LOOP_C_498 = 11'd898,
    COMP_LOOP_C_499 = 11'd899,
    COMP_LOOP_C_500 = 11'd900,
    COMP_LOOP_C_501 = 11'd901,
    COMP_LOOP_C_502 = 11'd902,
    COMP_LOOP_C_503 = 11'd903,
    COMP_LOOP_C_504 = 11'd904,
    COMP_LOOP_C_505 = 11'd905,
    COMP_LOOP_C_506 = 11'd906,
    COMP_LOOP_C_507 = 11'd907,
    COMP_LOOP_C_508 = 11'd908,
    COMP_LOOP_C_509 = 11'd909,
    COMP_LOOP_C_510 = 11'd910,
    COMP_LOOP_C_511 = 11'd911,
    COMP_LOOP_C_512 = 11'd912,
    COMP_LOOP_C_513 = 11'd913,
    COMP_LOOP_C_514 = 11'd914,
    COMP_LOOP_C_515 = 11'd915,
    COMP_LOOP_C_516 = 11'd916,
    COMP_LOOP_C_517 = 11'd917,
    COMP_LOOP_C_518 = 11'd918,
    COMP_LOOP_C_519 = 11'd919,
    COMP_LOOP_C_520 = 11'd920,
    COMP_LOOP_C_521 = 11'd921,
    COMP_LOOP_C_522 = 11'd922,
    COMP_LOOP_C_523 = 11'd923,
    COMP_LOOP_C_524 = 11'd924,
    COMP_LOOP_C_525 = 11'd925,
    COMP_LOOP_C_526 = 11'd926,
    COMP_LOOP_C_527 = 11'd927,
    COMP_LOOP_C_528 = 11'd928,
    COMP_LOOP_C_529 = 11'd929,
    COMP_LOOP_C_530 = 11'd930,
    COMP_LOOP_C_531 = 11'd931,
    COMP_LOOP_C_532 = 11'd932,
    COMP_LOOP_C_533 = 11'd933,
    COMP_LOOP_C_534 = 11'd934,
    COMP_LOOP_C_535 = 11'd935,
    COMP_LOOP_C_536 = 11'd936,
    COMP_LOOP_C_537 = 11'd937,
    COMP_LOOP_C_538 = 11'd938,
    COMP_LOOP_C_539 = 11'd939,
    COMP_LOOP_C_540 = 11'd940,
    COMP_LOOP_C_541 = 11'd941,
    COMP_LOOP_C_542 = 11'd942,
    COMP_LOOP_C_543 = 11'd943,
    COMP_LOOP_C_544 = 11'd944,
    COMP_LOOP_C_545 = 11'd945,
    COMP_LOOP_C_546 = 11'd946,
    COMP_LOOP_C_547 = 11'd947,
    COMP_LOOP_C_548 = 11'd948,
    COMP_LOOP_C_549 = 11'd949,
    COMP_LOOP_C_550 = 11'd950,
    COMP_LOOP_C_551 = 11'd951,
    COMP_LOOP_C_552 = 11'd952,
    COMP_LOOP_C_553 = 11'd953,
    COMP_LOOP_C_554 = 11'd954,
    COMP_LOOP_C_555 = 11'd955,
    COMP_LOOP_C_556 = 11'd956,
    COMP_LOOP_C_557 = 11'd957,
    COMP_LOOP_C_558 = 11'd958,
    COMP_LOOP_C_559 = 11'd959,
    COMP_LOOP_10_modExp_1_while_C_0 = 11'd960,
    COMP_LOOP_10_modExp_1_while_C_1 = 11'd961,
    COMP_LOOP_10_modExp_1_while_C_2 = 11'd962,
    COMP_LOOP_10_modExp_1_while_C_3 = 11'd963,
    COMP_LOOP_10_modExp_1_while_C_4 = 11'd964,
    COMP_LOOP_10_modExp_1_while_C_5 = 11'd965,
    COMP_LOOP_10_modExp_1_while_C_6 = 11'd966,
    COMP_LOOP_10_modExp_1_while_C_7 = 11'd967,
    COMP_LOOP_10_modExp_1_while_C_8 = 11'd968,
    COMP_LOOP_10_modExp_1_while_C_9 = 11'd969,
    COMP_LOOP_10_modExp_1_while_C_10 = 11'd970,
    COMP_LOOP_10_modExp_1_while_C_11 = 11'd971,
    COMP_LOOP_10_modExp_1_while_C_12 = 11'd972,
    COMP_LOOP_10_modExp_1_while_C_13 = 11'd973,
    COMP_LOOP_10_modExp_1_while_C_14 = 11'd974,
    COMP_LOOP_10_modExp_1_while_C_15 = 11'd975,
    COMP_LOOP_10_modExp_1_while_C_16 = 11'd976,
    COMP_LOOP_10_modExp_1_while_C_17 = 11'd977,
    COMP_LOOP_10_modExp_1_while_C_18 = 11'd978,
    COMP_LOOP_10_modExp_1_while_C_19 = 11'd979,
    COMP_LOOP_10_modExp_1_while_C_20 = 11'd980,
    COMP_LOOP_10_modExp_1_while_C_21 = 11'd981,
    COMP_LOOP_10_modExp_1_while_C_22 = 11'd982,
    COMP_LOOP_10_modExp_1_while_C_23 = 11'd983,
    COMP_LOOP_10_modExp_1_while_C_24 = 11'd984,
    COMP_LOOP_10_modExp_1_while_C_25 = 11'd985,
    COMP_LOOP_10_modExp_1_while_C_26 = 11'd986,
    COMP_LOOP_10_modExp_1_while_C_27 = 11'd987,
    COMP_LOOP_10_modExp_1_while_C_28 = 11'd988,
    COMP_LOOP_10_modExp_1_while_C_29 = 11'd989,
    COMP_LOOP_10_modExp_1_while_C_30 = 11'd990,
    COMP_LOOP_10_modExp_1_while_C_31 = 11'd991,
    COMP_LOOP_10_modExp_1_while_C_32 = 11'd992,
    COMP_LOOP_10_modExp_1_while_C_33 = 11'd993,
    COMP_LOOP_10_modExp_1_while_C_34 = 11'd994,
    COMP_LOOP_10_modExp_1_while_C_35 = 11'd995,
    COMP_LOOP_10_modExp_1_while_C_36 = 11'd996,
    COMP_LOOP_10_modExp_1_while_C_37 = 11'd997,
    COMP_LOOP_10_modExp_1_while_C_38 = 11'd998,
    COMP_LOOP_C_560 = 11'd999,
    COMP_LOOP_C_561 = 11'd1000,
    COMP_LOOP_C_562 = 11'd1001,
    COMP_LOOP_C_563 = 11'd1002,
    COMP_LOOP_C_564 = 11'd1003,
    COMP_LOOP_C_565 = 11'd1004,
    COMP_LOOP_C_566 = 11'd1005,
    COMP_LOOP_C_567 = 11'd1006,
    COMP_LOOP_C_568 = 11'd1007,
    COMP_LOOP_C_569 = 11'd1008,
    COMP_LOOP_C_570 = 11'd1009,
    COMP_LOOP_C_571 = 11'd1010,
    COMP_LOOP_C_572 = 11'd1011,
    COMP_LOOP_C_573 = 11'd1012,
    COMP_LOOP_C_574 = 11'd1013,
    COMP_LOOP_C_575 = 11'd1014,
    COMP_LOOP_C_576 = 11'd1015,
    COMP_LOOP_C_577 = 11'd1016,
    COMP_LOOP_C_578 = 11'd1017,
    COMP_LOOP_C_579 = 11'd1018,
    COMP_LOOP_C_580 = 11'd1019,
    COMP_LOOP_C_581 = 11'd1020,
    COMP_LOOP_C_582 = 11'd1021,
    COMP_LOOP_C_583 = 11'd1022,
    COMP_LOOP_C_584 = 11'd1023,
    COMP_LOOP_C_585 = 11'd1024,
    COMP_LOOP_C_586 = 11'd1025,
    COMP_LOOP_C_587 = 11'd1026,
    COMP_LOOP_C_588 = 11'd1027,
    COMP_LOOP_C_589 = 11'd1028,
    COMP_LOOP_C_590 = 11'd1029,
    COMP_LOOP_C_591 = 11'd1030,
    COMP_LOOP_C_592 = 11'd1031,
    COMP_LOOP_C_593 = 11'd1032,
    COMP_LOOP_C_594 = 11'd1033,
    COMP_LOOP_C_595 = 11'd1034,
    COMP_LOOP_C_596 = 11'd1035,
    COMP_LOOP_C_597 = 11'd1036,
    COMP_LOOP_C_598 = 11'd1037,
    COMP_LOOP_C_599 = 11'd1038,
    COMP_LOOP_C_600 = 11'd1039,
    COMP_LOOP_C_601 = 11'd1040,
    COMP_LOOP_C_602 = 11'd1041,
    COMP_LOOP_C_603 = 11'd1042,
    COMP_LOOP_C_604 = 11'd1043,
    COMP_LOOP_C_605 = 11'd1044,
    COMP_LOOP_C_606 = 11'd1045,
    COMP_LOOP_C_607 = 11'd1046,
    COMP_LOOP_C_608 = 11'd1047,
    COMP_LOOP_C_609 = 11'd1048,
    COMP_LOOP_C_610 = 11'd1049,
    COMP_LOOP_C_611 = 11'd1050,
    COMP_LOOP_C_612 = 11'd1051,
    COMP_LOOP_C_613 = 11'd1052,
    COMP_LOOP_C_614 = 11'd1053,
    COMP_LOOP_C_615 = 11'd1054,
    COMP_LOOP_C_616 = 11'd1055,
    COMP_LOOP_C_617 = 11'd1056,
    COMP_LOOP_C_618 = 11'd1057,
    COMP_LOOP_C_619 = 11'd1058,
    COMP_LOOP_C_620 = 11'd1059,
    COMP_LOOP_C_621 = 11'd1060,
    COMP_LOOP_11_modExp_1_while_C_0 = 11'd1061,
    COMP_LOOP_11_modExp_1_while_C_1 = 11'd1062,
    COMP_LOOP_11_modExp_1_while_C_2 = 11'd1063,
    COMP_LOOP_11_modExp_1_while_C_3 = 11'd1064,
    COMP_LOOP_11_modExp_1_while_C_4 = 11'd1065,
    COMP_LOOP_11_modExp_1_while_C_5 = 11'd1066,
    COMP_LOOP_11_modExp_1_while_C_6 = 11'd1067,
    COMP_LOOP_11_modExp_1_while_C_7 = 11'd1068,
    COMP_LOOP_11_modExp_1_while_C_8 = 11'd1069,
    COMP_LOOP_11_modExp_1_while_C_9 = 11'd1070,
    COMP_LOOP_11_modExp_1_while_C_10 = 11'd1071,
    COMP_LOOP_11_modExp_1_while_C_11 = 11'd1072,
    COMP_LOOP_11_modExp_1_while_C_12 = 11'd1073,
    COMP_LOOP_11_modExp_1_while_C_13 = 11'd1074,
    COMP_LOOP_11_modExp_1_while_C_14 = 11'd1075,
    COMP_LOOP_11_modExp_1_while_C_15 = 11'd1076,
    COMP_LOOP_11_modExp_1_while_C_16 = 11'd1077,
    COMP_LOOP_11_modExp_1_while_C_17 = 11'd1078,
    COMP_LOOP_11_modExp_1_while_C_18 = 11'd1079,
    COMP_LOOP_11_modExp_1_while_C_19 = 11'd1080,
    COMP_LOOP_11_modExp_1_while_C_20 = 11'd1081,
    COMP_LOOP_11_modExp_1_while_C_21 = 11'd1082,
    COMP_LOOP_11_modExp_1_while_C_22 = 11'd1083,
    COMP_LOOP_11_modExp_1_while_C_23 = 11'd1084,
    COMP_LOOP_11_modExp_1_while_C_24 = 11'd1085,
    COMP_LOOP_11_modExp_1_while_C_25 = 11'd1086,
    COMP_LOOP_11_modExp_1_while_C_26 = 11'd1087,
    COMP_LOOP_11_modExp_1_while_C_27 = 11'd1088,
    COMP_LOOP_11_modExp_1_while_C_28 = 11'd1089,
    COMP_LOOP_11_modExp_1_while_C_29 = 11'd1090,
    COMP_LOOP_11_modExp_1_while_C_30 = 11'd1091,
    COMP_LOOP_11_modExp_1_while_C_31 = 11'd1092,
    COMP_LOOP_11_modExp_1_while_C_32 = 11'd1093,
    COMP_LOOP_11_modExp_1_while_C_33 = 11'd1094,
    COMP_LOOP_11_modExp_1_while_C_34 = 11'd1095,
    COMP_LOOP_11_modExp_1_while_C_35 = 11'd1096,
    COMP_LOOP_11_modExp_1_while_C_36 = 11'd1097,
    COMP_LOOP_11_modExp_1_while_C_37 = 11'd1098,
    COMP_LOOP_11_modExp_1_while_C_38 = 11'd1099,
    COMP_LOOP_C_622 = 11'd1100,
    COMP_LOOP_C_623 = 11'd1101,
    COMP_LOOP_C_624 = 11'd1102,
    COMP_LOOP_C_625 = 11'd1103,
    COMP_LOOP_C_626 = 11'd1104,
    COMP_LOOP_C_627 = 11'd1105,
    COMP_LOOP_C_628 = 11'd1106,
    COMP_LOOP_C_629 = 11'd1107,
    COMP_LOOP_C_630 = 11'd1108,
    COMP_LOOP_C_631 = 11'd1109,
    COMP_LOOP_C_632 = 11'd1110,
    COMP_LOOP_C_633 = 11'd1111,
    COMP_LOOP_C_634 = 11'd1112,
    COMP_LOOP_C_635 = 11'd1113,
    COMP_LOOP_C_636 = 11'd1114,
    COMP_LOOP_C_637 = 11'd1115,
    COMP_LOOP_C_638 = 11'd1116,
    COMP_LOOP_C_639 = 11'd1117,
    COMP_LOOP_C_640 = 11'd1118,
    COMP_LOOP_C_641 = 11'd1119,
    COMP_LOOP_C_642 = 11'd1120,
    COMP_LOOP_C_643 = 11'd1121,
    COMP_LOOP_C_644 = 11'd1122,
    COMP_LOOP_C_645 = 11'd1123,
    COMP_LOOP_C_646 = 11'd1124,
    COMP_LOOP_C_647 = 11'd1125,
    COMP_LOOP_C_648 = 11'd1126,
    COMP_LOOP_C_649 = 11'd1127,
    COMP_LOOP_C_650 = 11'd1128,
    COMP_LOOP_C_651 = 11'd1129,
    COMP_LOOP_C_652 = 11'd1130,
    COMP_LOOP_C_653 = 11'd1131,
    COMP_LOOP_C_654 = 11'd1132,
    COMP_LOOP_C_655 = 11'd1133,
    COMP_LOOP_C_656 = 11'd1134,
    COMP_LOOP_C_657 = 11'd1135,
    COMP_LOOP_C_658 = 11'd1136,
    COMP_LOOP_C_659 = 11'd1137,
    COMP_LOOP_C_660 = 11'd1138,
    COMP_LOOP_C_661 = 11'd1139,
    COMP_LOOP_C_662 = 11'd1140,
    COMP_LOOP_C_663 = 11'd1141,
    COMP_LOOP_C_664 = 11'd1142,
    COMP_LOOP_C_665 = 11'd1143,
    COMP_LOOP_C_666 = 11'd1144,
    COMP_LOOP_C_667 = 11'd1145,
    COMP_LOOP_C_668 = 11'd1146,
    COMP_LOOP_C_669 = 11'd1147,
    COMP_LOOP_C_670 = 11'd1148,
    COMP_LOOP_C_671 = 11'd1149,
    COMP_LOOP_C_672 = 11'd1150,
    COMP_LOOP_C_673 = 11'd1151,
    COMP_LOOP_C_674 = 11'd1152,
    COMP_LOOP_C_675 = 11'd1153,
    COMP_LOOP_C_676 = 11'd1154,
    COMP_LOOP_C_677 = 11'd1155,
    COMP_LOOP_C_678 = 11'd1156,
    COMP_LOOP_C_679 = 11'd1157,
    COMP_LOOP_C_680 = 11'd1158,
    COMP_LOOP_C_681 = 11'd1159,
    COMP_LOOP_C_682 = 11'd1160,
    COMP_LOOP_C_683 = 11'd1161,
    COMP_LOOP_12_modExp_1_while_C_0 = 11'd1162,
    COMP_LOOP_12_modExp_1_while_C_1 = 11'd1163,
    COMP_LOOP_12_modExp_1_while_C_2 = 11'd1164,
    COMP_LOOP_12_modExp_1_while_C_3 = 11'd1165,
    COMP_LOOP_12_modExp_1_while_C_4 = 11'd1166,
    COMP_LOOP_12_modExp_1_while_C_5 = 11'd1167,
    COMP_LOOP_12_modExp_1_while_C_6 = 11'd1168,
    COMP_LOOP_12_modExp_1_while_C_7 = 11'd1169,
    COMP_LOOP_12_modExp_1_while_C_8 = 11'd1170,
    COMP_LOOP_12_modExp_1_while_C_9 = 11'd1171,
    COMP_LOOP_12_modExp_1_while_C_10 = 11'd1172,
    COMP_LOOP_12_modExp_1_while_C_11 = 11'd1173,
    COMP_LOOP_12_modExp_1_while_C_12 = 11'd1174,
    COMP_LOOP_12_modExp_1_while_C_13 = 11'd1175,
    COMP_LOOP_12_modExp_1_while_C_14 = 11'd1176,
    COMP_LOOP_12_modExp_1_while_C_15 = 11'd1177,
    COMP_LOOP_12_modExp_1_while_C_16 = 11'd1178,
    COMP_LOOP_12_modExp_1_while_C_17 = 11'd1179,
    COMP_LOOP_12_modExp_1_while_C_18 = 11'd1180,
    COMP_LOOP_12_modExp_1_while_C_19 = 11'd1181,
    COMP_LOOP_12_modExp_1_while_C_20 = 11'd1182,
    COMP_LOOP_12_modExp_1_while_C_21 = 11'd1183,
    COMP_LOOP_12_modExp_1_while_C_22 = 11'd1184,
    COMP_LOOP_12_modExp_1_while_C_23 = 11'd1185,
    COMP_LOOP_12_modExp_1_while_C_24 = 11'd1186,
    COMP_LOOP_12_modExp_1_while_C_25 = 11'd1187,
    COMP_LOOP_12_modExp_1_while_C_26 = 11'd1188,
    COMP_LOOP_12_modExp_1_while_C_27 = 11'd1189,
    COMP_LOOP_12_modExp_1_while_C_28 = 11'd1190,
    COMP_LOOP_12_modExp_1_while_C_29 = 11'd1191,
    COMP_LOOP_12_modExp_1_while_C_30 = 11'd1192,
    COMP_LOOP_12_modExp_1_while_C_31 = 11'd1193,
    COMP_LOOP_12_modExp_1_while_C_32 = 11'd1194,
    COMP_LOOP_12_modExp_1_while_C_33 = 11'd1195,
    COMP_LOOP_12_modExp_1_while_C_34 = 11'd1196,
    COMP_LOOP_12_modExp_1_while_C_35 = 11'd1197,
    COMP_LOOP_12_modExp_1_while_C_36 = 11'd1198,
    COMP_LOOP_12_modExp_1_while_C_37 = 11'd1199,
    COMP_LOOP_12_modExp_1_while_C_38 = 11'd1200,
    COMP_LOOP_C_684 = 11'd1201,
    COMP_LOOP_C_685 = 11'd1202,
    COMP_LOOP_C_686 = 11'd1203,
    COMP_LOOP_C_687 = 11'd1204,
    COMP_LOOP_C_688 = 11'd1205,
    COMP_LOOP_C_689 = 11'd1206,
    COMP_LOOP_C_690 = 11'd1207,
    COMP_LOOP_C_691 = 11'd1208,
    COMP_LOOP_C_692 = 11'd1209,
    COMP_LOOP_C_693 = 11'd1210,
    COMP_LOOP_C_694 = 11'd1211,
    COMP_LOOP_C_695 = 11'd1212,
    COMP_LOOP_C_696 = 11'd1213,
    COMP_LOOP_C_697 = 11'd1214,
    COMP_LOOP_C_698 = 11'd1215,
    COMP_LOOP_C_699 = 11'd1216,
    COMP_LOOP_C_700 = 11'd1217,
    COMP_LOOP_C_701 = 11'd1218,
    COMP_LOOP_C_702 = 11'd1219,
    COMP_LOOP_C_703 = 11'd1220,
    COMP_LOOP_C_704 = 11'd1221,
    COMP_LOOP_C_705 = 11'd1222,
    COMP_LOOP_C_706 = 11'd1223,
    COMP_LOOP_C_707 = 11'd1224,
    COMP_LOOP_C_708 = 11'd1225,
    COMP_LOOP_C_709 = 11'd1226,
    COMP_LOOP_C_710 = 11'd1227,
    COMP_LOOP_C_711 = 11'd1228,
    COMP_LOOP_C_712 = 11'd1229,
    COMP_LOOP_C_713 = 11'd1230,
    COMP_LOOP_C_714 = 11'd1231,
    COMP_LOOP_C_715 = 11'd1232,
    COMP_LOOP_C_716 = 11'd1233,
    COMP_LOOP_C_717 = 11'd1234,
    COMP_LOOP_C_718 = 11'd1235,
    COMP_LOOP_C_719 = 11'd1236,
    COMP_LOOP_C_720 = 11'd1237,
    COMP_LOOP_C_721 = 11'd1238,
    COMP_LOOP_C_722 = 11'd1239,
    COMP_LOOP_C_723 = 11'd1240,
    COMP_LOOP_C_724 = 11'd1241,
    COMP_LOOP_C_725 = 11'd1242,
    COMP_LOOP_C_726 = 11'd1243,
    COMP_LOOP_C_727 = 11'd1244,
    COMP_LOOP_C_728 = 11'd1245,
    COMP_LOOP_C_729 = 11'd1246,
    COMP_LOOP_C_730 = 11'd1247,
    COMP_LOOP_C_731 = 11'd1248,
    COMP_LOOP_C_732 = 11'd1249,
    COMP_LOOP_C_733 = 11'd1250,
    COMP_LOOP_C_734 = 11'd1251,
    COMP_LOOP_C_735 = 11'd1252,
    COMP_LOOP_C_736 = 11'd1253,
    COMP_LOOP_C_737 = 11'd1254,
    COMP_LOOP_C_738 = 11'd1255,
    COMP_LOOP_C_739 = 11'd1256,
    COMP_LOOP_C_740 = 11'd1257,
    COMP_LOOP_C_741 = 11'd1258,
    COMP_LOOP_C_742 = 11'd1259,
    COMP_LOOP_C_743 = 11'd1260,
    COMP_LOOP_C_744 = 11'd1261,
    COMP_LOOP_C_745 = 11'd1262,
    COMP_LOOP_13_modExp_1_while_C_0 = 11'd1263,
    COMP_LOOP_13_modExp_1_while_C_1 = 11'd1264,
    COMP_LOOP_13_modExp_1_while_C_2 = 11'd1265,
    COMP_LOOP_13_modExp_1_while_C_3 = 11'd1266,
    COMP_LOOP_13_modExp_1_while_C_4 = 11'd1267,
    COMP_LOOP_13_modExp_1_while_C_5 = 11'd1268,
    COMP_LOOP_13_modExp_1_while_C_6 = 11'd1269,
    COMP_LOOP_13_modExp_1_while_C_7 = 11'd1270,
    COMP_LOOP_13_modExp_1_while_C_8 = 11'd1271,
    COMP_LOOP_13_modExp_1_while_C_9 = 11'd1272,
    COMP_LOOP_13_modExp_1_while_C_10 = 11'd1273,
    COMP_LOOP_13_modExp_1_while_C_11 = 11'd1274,
    COMP_LOOP_13_modExp_1_while_C_12 = 11'd1275,
    COMP_LOOP_13_modExp_1_while_C_13 = 11'd1276,
    COMP_LOOP_13_modExp_1_while_C_14 = 11'd1277,
    COMP_LOOP_13_modExp_1_while_C_15 = 11'd1278,
    COMP_LOOP_13_modExp_1_while_C_16 = 11'd1279,
    COMP_LOOP_13_modExp_1_while_C_17 = 11'd1280,
    COMP_LOOP_13_modExp_1_while_C_18 = 11'd1281,
    COMP_LOOP_13_modExp_1_while_C_19 = 11'd1282,
    COMP_LOOP_13_modExp_1_while_C_20 = 11'd1283,
    COMP_LOOP_13_modExp_1_while_C_21 = 11'd1284,
    COMP_LOOP_13_modExp_1_while_C_22 = 11'd1285,
    COMP_LOOP_13_modExp_1_while_C_23 = 11'd1286,
    COMP_LOOP_13_modExp_1_while_C_24 = 11'd1287,
    COMP_LOOP_13_modExp_1_while_C_25 = 11'd1288,
    COMP_LOOP_13_modExp_1_while_C_26 = 11'd1289,
    COMP_LOOP_13_modExp_1_while_C_27 = 11'd1290,
    COMP_LOOP_13_modExp_1_while_C_28 = 11'd1291,
    COMP_LOOP_13_modExp_1_while_C_29 = 11'd1292,
    COMP_LOOP_13_modExp_1_while_C_30 = 11'd1293,
    COMP_LOOP_13_modExp_1_while_C_31 = 11'd1294,
    COMP_LOOP_13_modExp_1_while_C_32 = 11'd1295,
    COMP_LOOP_13_modExp_1_while_C_33 = 11'd1296,
    COMP_LOOP_13_modExp_1_while_C_34 = 11'd1297,
    COMP_LOOP_13_modExp_1_while_C_35 = 11'd1298,
    COMP_LOOP_13_modExp_1_while_C_36 = 11'd1299,
    COMP_LOOP_13_modExp_1_while_C_37 = 11'd1300,
    COMP_LOOP_13_modExp_1_while_C_38 = 11'd1301,
    COMP_LOOP_C_746 = 11'd1302,
    COMP_LOOP_C_747 = 11'd1303,
    COMP_LOOP_C_748 = 11'd1304,
    COMP_LOOP_C_749 = 11'd1305,
    COMP_LOOP_C_750 = 11'd1306,
    COMP_LOOP_C_751 = 11'd1307,
    COMP_LOOP_C_752 = 11'd1308,
    COMP_LOOP_C_753 = 11'd1309,
    COMP_LOOP_C_754 = 11'd1310,
    COMP_LOOP_C_755 = 11'd1311,
    COMP_LOOP_C_756 = 11'd1312,
    COMP_LOOP_C_757 = 11'd1313,
    COMP_LOOP_C_758 = 11'd1314,
    COMP_LOOP_C_759 = 11'd1315,
    COMP_LOOP_C_760 = 11'd1316,
    COMP_LOOP_C_761 = 11'd1317,
    COMP_LOOP_C_762 = 11'd1318,
    COMP_LOOP_C_763 = 11'd1319,
    COMP_LOOP_C_764 = 11'd1320,
    COMP_LOOP_C_765 = 11'd1321,
    COMP_LOOP_C_766 = 11'd1322,
    COMP_LOOP_C_767 = 11'd1323,
    COMP_LOOP_C_768 = 11'd1324,
    COMP_LOOP_C_769 = 11'd1325,
    COMP_LOOP_C_770 = 11'd1326,
    COMP_LOOP_C_771 = 11'd1327,
    COMP_LOOP_C_772 = 11'd1328,
    COMP_LOOP_C_773 = 11'd1329,
    COMP_LOOP_C_774 = 11'd1330,
    COMP_LOOP_C_775 = 11'd1331,
    COMP_LOOP_C_776 = 11'd1332,
    COMP_LOOP_C_777 = 11'd1333,
    COMP_LOOP_C_778 = 11'd1334,
    COMP_LOOP_C_779 = 11'd1335,
    COMP_LOOP_C_780 = 11'd1336,
    COMP_LOOP_C_781 = 11'd1337,
    COMP_LOOP_C_782 = 11'd1338,
    COMP_LOOP_C_783 = 11'd1339,
    COMP_LOOP_C_784 = 11'd1340,
    COMP_LOOP_C_785 = 11'd1341,
    COMP_LOOP_C_786 = 11'd1342,
    COMP_LOOP_C_787 = 11'd1343,
    COMP_LOOP_C_788 = 11'd1344,
    COMP_LOOP_C_789 = 11'd1345,
    COMP_LOOP_C_790 = 11'd1346,
    COMP_LOOP_C_791 = 11'd1347,
    COMP_LOOP_C_792 = 11'd1348,
    COMP_LOOP_C_793 = 11'd1349,
    COMP_LOOP_C_794 = 11'd1350,
    COMP_LOOP_C_795 = 11'd1351,
    COMP_LOOP_C_796 = 11'd1352,
    COMP_LOOP_C_797 = 11'd1353,
    COMP_LOOP_C_798 = 11'd1354,
    COMP_LOOP_C_799 = 11'd1355,
    COMP_LOOP_C_800 = 11'd1356,
    COMP_LOOP_C_801 = 11'd1357,
    COMP_LOOP_C_802 = 11'd1358,
    COMP_LOOP_C_803 = 11'd1359,
    COMP_LOOP_C_804 = 11'd1360,
    COMP_LOOP_C_805 = 11'd1361,
    COMP_LOOP_C_806 = 11'd1362,
    COMP_LOOP_C_807 = 11'd1363,
    COMP_LOOP_14_modExp_1_while_C_0 = 11'd1364,
    COMP_LOOP_14_modExp_1_while_C_1 = 11'd1365,
    COMP_LOOP_14_modExp_1_while_C_2 = 11'd1366,
    COMP_LOOP_14_modExp_1_while_C_3 = 11'd1367,
    COMP_LOOP_14_modExp_1_while_C_4 = 11'd1368,
    COMP_LOOP_14_modExp_1_while_C_5 = 11'd1369,
    COMP_LOOP_14_modExp_1_while_C_6 = 11'd1370,
    COMP_LOOP_14_modExp_1_while_C_7 = 11'd1371,
    COMP_LOOP_14_modExp_1_while_C_8 = 11'd1372,
    COMP_LOOP_14_modExp_1_while_C_9 = 11'd1373,
    COMP_LOOP_14_modExp_1_while_C_10 = 11'd1374,
    COMP_LOOP_14_modExp_1_while_C_11 = 11'd1375,
    COMP_LOOP_14_modExp_1_while_C_12 = 11'd1376,
    COMP_LOOP_14_modExp_1_while_C_13 = 11'd1377,
    COMP_LOOP_14_modExp_1_while_C_14 = 11'd1378,
    COMP_LOOP_14_modExp_1_while_C_15 = 11'd1379,
    COMP_LOOP_14_modExp_1_while_C_16 = 11'd1380,
    COMP_LOOP_14_modExp_1_while_C_17 = 11'd1381,
    COMP_LOOP_14_modExp_1_while_C_18 = 11'd1382,
    COMP_LOOP_14_modExp_1_while_C_19 = 11'd1383,
    COMP_LOOP_14_modExp_1_while_C_20 = 11'd1384,
    COMP_LOOP_14_modExp_1_while_C_21 = 11'd1385,
    COMP_LOOP_14_modExp_1_while_C_22 = 11'd1386,
    COMP_LOOP_14_modExp_1_while_C_23 = 11'd1387,
    COMP_LOOP_14_modExp_1_while_C_24 = 11'd1388,
    COMP_LOOP_14_modExp_1_while_C_25 = 11'd1389,
    COMP_LOOP_14_modExp_1_while_C_26 = 11'd1390,
    COMP_LOOP_14_modExp_1_while_C_27 = 11'd1391,
    COMP_LOOP_14_modExp_1_while_C_28 = 11'd1392,
    COMP_LOOP_14_modExp_1_while_C_29 = 11'd1393,
    COMP_LOOP_14_modExp_1_while_C_30 = 11'd1394,
    COMP_LOOP_14_modExp_1_while_C_31 = 11'd1395,
    COMP_LOOP_14_modExp_1_while_C_32 = 11'd1396,
    COMP_LOOP_14_modExp_1_while_C_33 = 11'd1397,
    COMP_LOOP_14_modExp_1_while_C_34 = 11'd1398,
    COMP_LOOP_14_modExp_1_while_C_35 = 11'd1399,
    COMP_LOOP_14_modExp_1_while_C_36 = 11'd1400,
    COMP_LOOP_14_modExp_1_while_C_37 = 11'd1401,
    COMP_LOOP_14_modExp_1_while_C_38 = 11'd1402,
    COMP_LOOP_C_808 = 11'd1403,
    COMP_LOOP_C_809 = 11'd1404,
    COMP_LOOP_C_810 = 11'd1405,
    COMP_LOOP_C_811 = 11'd1406,
    COMP_LOOP_C_812 = 11'd1407,
    COMP_LOOP_C_813 = 11'd1408,
    COMP_LOOP_C_814 = 11'd1409,
    COMP_LOOP_C_815 = 11'd1410,
    COMP_LOOP_C_816 = 11'd1411,
    COMP_LOOP_C_817 = 11'd1412,
    COMP_LOOP_C_818 = 11'd1413,
    COMP_LOOP_C_819 = 11'd1414,
    COMP_LOOP_C_820 = 11'd1415,
    COMP_LOOP_C_821 = 11'd1416,
    COMP_LOOP_C_822 = 11'd1417,
    COMP_LOOP_C_823 = 11'd1418,
    COMP_LOOP_C_824 = 11'd1419,
    COMP_LOOP_C_825 = 11'd1420,
    COMP_LOOP_C_826 = 11'd1421,
    COMP_LOOP_C_827 = 11'd1422,
    COMP_LOOP_C_828 = 11'd1423,
    COMP_LOOP_C_829 = 11'd1424,
    COMP_LOOP_C_830 = 11'd1425,
    COMP_LOOP_C_831 = 11'd1426,
    COMP_LOOP_C_832 = 11'd1427,
    COMP_LOOP_C_833 = 11'd1428,
    COMP_LOOP_C_834 = 11'd1429,
    COMP_LOOP_C_835 = 11'd1430,
    COMP_LOOP_C_836 = 11'd1431,
    COMP_LOOP_C_837 = 11'd1432,
    COMP_LOOP_C_838 = 11'd1433,
    COMP_LOOP_C_839 = 11'd1434,
    COMP_LOOP_C_840 = 11'd1435,
    COMP_LOOP_C_841 = 11'd1436,
    COMP_LOOP_C_842 = 11'd1437,
    COMP_LOOP_C_843 = 11'd1438,
    COMP_LOOP_C_844 = 11'd1439,
    COMP_LOOP_C_845 = 11'd1440,
    COMP_LOOP_C_846 = 11'd1441,
    COMP_LOOP_C_847 = 11'd1442,
    COMP_LOOP_C_848 = 11'd1443,
    COMP_LOOP_C_849 = 11'd1444,
    COMP_LOOP_C_850 = 11'd1445,
    COMP_LOOP_C_851 = 11'd1446,
    COMP_LOOP_C_852 = 11'd1447,
    COMP_LOOP_C_853 = 11'd1448,
    COMP_LOOP_C_854 = 11'd1449,
    COMP_LOOP_C_855 = 11'd1450,
    COMP_LOOP_C_856 = 11'd1451,
    COMP_LOOP_C_857 = 11'd1452,
    COMP_LOOP_C_858 = 11'd1453,
    COMP_LOOP_C_859 = 11'd1454,
    COMP_LOOP_C_860 = 11'd1455,
    COMP_LOOP_C_861 = 11'd1456,
    COMP_LOOP_C_862 = 11'd1457,
    COMP_LOOP_C_863 = 11'd1458,
    COMP_LOOP_C_864 = 11'd1459,
    COMP_LOOP_C_865 = 11'd1460,
    COMP_LOOP_C_866 = 11'd1461,
    COMP_LOOP_C_867 = 11'd1462,
    COMP_LOOP_C_868 = 11'd1463,
    COMP_LOOP_C_869 = 11'd1464,
    COMP_LOOP_15_modExp_1_while_C_0 = 11'd1465,
    COMP_LOOP_15_modExp_1_while_C_1 = 11'd1466,
    COMP_LOOP_15_modExp_1_while_C_2 = 11'd1467,
    COMP_LOOP_15_modExp_1_while_C_3 = 11'd1468,
    COMP_LOOP_15_modExp_1_while_C_4 = 11'd1469,
    COMP_LOOP_15_modExp_1_while_C_5 = 11'd1470,
    COMP_LOOP_15_modExp_1_while_C_6 = 11'd1471,
    COMP_LOOP_15_modExp_1_while_C_7 = 11'd1472,
    COMP_LOOP_15_modExp_1_while_C_8 = 11'd1473,
    COMP_LOOP_15_modExp_1_while_C_9 = 11'd1474,
    COMP_LOOP_15_modExp_1_while_C_10 = 11'd1475,
    COMP_LOOP_15_modExp_1_while_C_11 = 11'd1476,
    COMP_LOOP_15_modExp_1_while_C_12 = 11'd1477,
    COMP_LOOP_15_modExp_1_while_C_13 = 11'd1478,
    COMP_LOOP_15_modExp_1_while_C_14 = 11'd1479,
    COMP_LOOP_15_modExp_1_while_C_15 = 11'd1480,
    COMP_LOOP_15_modExp_1_while_C_16 = 11'd1481,
    COMP_LOOP_15_modExp_1_while_C_17 = 11'd1482,
    COMP_LOOP_15_modExp_1_while_C_18 = 11'd1483,
    COMP_LOOP_15_modExp_1_while_C_19 = 11'd1484,
    COMP_LOOP_15_modExp_1_while_C_20 = 11'd1485,
    COMP_LOOP_15_modExp_1_while_C_21 = 11'd1486,
    COMP_LOOP_15_modExp_1_while_C_22 = 11'd1487,
    COMP_LOOP_15_modExp_1_while_C_23 = 11'd1488,
    COMP_LOOP_15_modExp_1_while_C_24 = 11'd1489,
    COMP_LOOP_15_modExp_1_while_C_25 = 11'd1490,
    COMP_LOOP_15_modExp_1_while_C_26 = 11'd1491,
    COMP_LOOP_15_modExp_1_while_C_27 = 11'd1492,
    COMP_LOOP_15_modExp_1_while_C_28 = 11'd1493,
    COMP_LOOP_15_modExp_1_while_C_29 = 11'd1494,
    COMP_LOOP_15_modExp_1_while_C_30 = 11'd1495,
    COMP_LOOP_15_modExp_1_while_C_31 = 11'd1496,
    COMP_LOOP_15_modExp_1_while_C_32 = 11'd1497,
    COMP_LOOP_15_modExp_1_while_C_33 = 11'd1498,
    COMP_LOOP_15_modExp_1_while_C_34 = 11'd1499,
    COMP_LOOP_15_modExp_1_while_C_35 = 11'd1500,
    COMP_LOOP_15_modExp_1_while_C_36 = 11'd1501,
    COMP_LOOP_15_modExp_1_while_C_37 = 11'd1502,
    COMP_LOOP_15_modExp_1_while_C_38 = 11'd1503,
    COMP_LOOP_C_870 = 11'd1504,
    COMP_LOOP_C_871 = 11'd1505,
    COMP_LOOP_C_872 = 11'd1506,
    COMP_LOOP_C_873 = 11'd1507,
    COMP_LOOP_C_874 = 11'd1508,
    COMP_LOOP_C_875 = 11'd1509,
    COMP_LOOP_C_876 = 11'd1510,
    COMP_LOOP_C_877 = 11'd1511,
    COMP_LOOP_C_878 = 11'd1512,
    COMP_LOOP_C_879 = 11'd1513,
    COMP_LOOP_C_880 = 11'd1514,
    COMP_LOOP_C_881 = 11'd1515,
    COMP_LOOP_C_882 = 11'd1516,
    COMP_LOOP_C_883 = 11'd1517,
    COMP_LOOP_C_884 = 11'd1518,
    COMP_LOOP_C_885 = 11'd1519,
    COMP_LOOP_C_886 = 11'd1520,
    COMP_LOOP_C_887 = 11'd1521,
    COMP_LOOP_C_888 = 11'd1522,
    COMP_LOOP_C_889 = 11'd1523,
    COMP_LOOP_C_890 = 11'd1524,
    COMP_LOOP_C_891 = 11'd1525,
    COMP_LOOP_C_892 = 11'd1526,
    COMP_LOOP_C_893 = 11'd1527,
    COMP_LOOP_C_894 = 11'd1528,
    COMP_LOOP_C_895 = 11'd1529,
    COMP_LOOP_C_896 = 11'd1530,
    COMP_LOOP_C_897 = 11'd1531,
    COMP_LOOP_C_898 = 11'd1532,
    COMP_LOOP_C_899 = 11'd1533,
    COMP_LOOP_C_900 = 11'd1534,
    COMP_LOOP_C_901 = 11'd1535,
    COMP_LOOP_C_902 = 11'd1536,
    COMP_LOOP_C_903 = 11'd1537,
    COMP_LOOP_C_904 = 11'd1538,
    COMP_LOOP_C_905 = 11'd1539,
    COMP_LOOP_C_906 = 11'd1540,
    COMP_LOOP_C_907 = 11'd1541,
    COMP_LOOP_C_908 = 11'd1542,
    COMP_LOOP_C_909 = 11'd1543,
    COMP_LOOP_C_910 = 11'd1544,
    COMP_LOOP_C_911 = 11'd1545,
    COMP_LOOP_C_912 = 11'd1546,
    COMP_LOOP_C_913 = 11'd1547,
    COMP_LOOP_C_914 = 11'd1548,
    COMP_LOOP_C_915 = 11'd1549,
    COMP_LOOP_C_916 = 11'd1550,
    COMP_LOOP_C_917 = 11'd1551,
    COMP_LOOP_C_918 = 11'd1552,
    COMP_LOOP_C_919 = 11'd1553,
    COMP_LOOP_C_920 = 11'd1554,
    COMP_LOOP_C_921 = 11'd1555,
    COMP_LOOP_C_922 = 11'd1556,
    COMP_LOOP_C_923 = 11'd1557,
    COMP_LOOP_C_924 = 11'd1558,
    COMP_LOOP_C_925 = 11'd1559,
    COMP_LOOP_C_926 = 11'd1560,
    COMP_LOOP_C_927 = 11'd1561,
    COMP_LOOP_C_928 = 11'd1562,
    COMP_LOOP_C_929 = 11'd1563,
    COMP_LOOP_C_930 = 11'd1564,
    COMP_LOOP_C_931 = 11'd1565,
    COMP_LOOP_16_modExp_1_while_C_0 = 11'd1566,
    COMP_LOOP_16_modExp_1_while_C_1 = 11'd1567,
    COMP_LOOP_16_modExp_1_while_C_2 = 11'd1568,
    COMP_LOOP_16_modExp_1_while_C_3 = 11'd1569,
    COMP_LOOP_16_modExp_1_while_C_4 = 11'd1570,
    COMP_LOOP_16_modExp_1_while_C_5 = 11'd1571,
    COMP_LOOP_16_modExp_1_while_C_6 = 11'd1572,
    COMP_LOOP_16_modExp_1_while_C_7 = 11'd1573,
    COMP_LOOP_16_modExp_1_while_C_8 = 11'd1574,
    COMP_LOOP_16_modExp_1_while_C_9 = 11'd1575,
    COMP_LOOP_16_modExp_1_while_C_10 = 11'd1576,
    COMP_LOOP_16_modExp_1_while_C_11 = 11'd1577,
    COMP_LOOP_16_modExp_1_while_C_12 = 11'd1578,
    COMP_LOOP_16_modExp_1_while_C_13 = 11'd1579,
    COMP_LOOP_16_modExp_1_while_C_14 = 11'd1580,
    COMP_LOOP_16_modExp_1_while_C_15 = 11'd1581,
    COMP_LOOP_16_modExp_1_while_C_16 = 11'd1582,
    COMP_LOOP_16_modExp_1_while_C_17 = 11'd1583,
    COMP_LOOP_16_modExp_1_while_C_18 = 11'd1584,
    COMP_LOOP_16_modExp_1_while_C_19 = 11'd1585,
    COMP_LOOP_16_modExp_1_while_C_20 = 11'd1586,
    COMP_LOOP_16_modExp_1_while_C_21 = 11'd1587,
    COMP_LOOP_16_modExp_1_while_C_22 = 11'd1588,
    COMP_LOOP_16_modExp_1_while_C_23 = 11'd1589,
    COMP_LOOP_16_modExp_1_while_C_24 = 11'd1590,
    COMP_LOOP_16_modExp_1_while_C_25 = 11'd1591,
    COMP_LOOP_16_modExp_1_while_C_26 = 11'd1592,
    COMP_LOOP_16_modExp_1_while_C_27 = 11'd1593,
    COMP_LOOP_16_modExp_1_while_C_28 = 11'd1594,
    COMP_LOOP_16_modExp_1_while_C_29 = 11'd1595,
    COMP_LOOP_16_modExp_1_while_C_30 = 11'd1596,
    COMP_LOOP_16_modExp_1_while_C_31 = 11'd1597,
    COMP_LOOP_16_modExp_1_while_C_32 = 11'd1598,
    COMP_LOOP_16_modExp_1_while_C_33 = 11'd1599,
    COMP_LOOP_16_modExp_1_while_C_34 = 11'd1600,
    COMP_LOOP_16_modExp_1_while_C_35 = 11'd1601,
    COMP_LOOP_16_modExp_1_while_C_36 = 11'd1602,
    COMP_LOOP_16_modExp_1_while_C_37 = 11'd1603,
    COMP_LOOP_16_modExp_1_while_C_38 = 11'd1604,
    COMP_LOOP_C_932 = 11'd1605,
    COMP_LOOP_C_933 = 11'd1606,
    COMP_LOOP_C_934 = 11'd1607,
    COMP_LOOP_C_935 = 11'd1608,
    COMP_LOOP_C_936 = 11'd1609,
    COMP_LOOP_C_937 = 11'd1610,
    COMP_LOOP_C_938 = 11'd1611,
    COMP_LOOP_C_939 = 11'd1612,
    COMP_LOOP_C_940 = 11'd1613,
    COMP_LOOP_C_941 = 11'd1614,
    COMP_LOOP_C_942 = 11'd1615,
    COMP_LOOP_C_943 = 11'd1616,
    COMP_LOOP_C_944 = 11'd1617,
    COMP_LOOP_C_945 = 11'd1618,
    COMP_LOOP_C_946 = 11'd1619,
    COMP_LOOP_C_947 = 11'd1620,
    COMP_LOOP_C_948 = 11'd1621,
    COMP_LOOP_C_949 = 11'd1622,
    COMP_LOOP_C_950 = 11'd1623,
    COMP_LOOP_C_951 = 11'd1624,
    COMP_LOOP_C_952 = 11'd1625,
    COMP_LOOP_C_953 = 11'd1626,
    COMP_LOOP_C_954 = 11'd1627,
    COMP_LOOP_C_955 = 11'd1628,
    COMP_LOOP_C_956 = 11'd1629,
    COMP_LOOP_C_957 = 11'd1630,
    COMP_LOOP_C_958 = 11'd1631,
    COMP_LOOP_C_959 = 11'd1632,
    COMP_LOOP_C_960 = 11'd1633,
    COMP_LOOP_C_961 = 11'd1634,
    COMP_LOOP_C_962 = 11'd1635,
    COMP_LOOP_C_963 = 11'd1636,
    COMP_LOOP_C_964 = 11'd1637,
    COMP_LOOP_C_965 = 11'd1638,
    COMP_LOOP_C_966 = 11'd1639,
    COMP_LOOP_C_967 = 11'd1640,
    COMP_LOOP_C_968 = 11'd1641,
    COMP_LOOP_C_969 = 11'd1642,
    COMP_LOOP_C_970 = 11'd1643,
    COMP_LOOP_C_971 = 11'd1644,
    COMP_LOOP_C_972 = 11'd1645,
    COMP_LOOP_C_973 = 11'd1646,
    COMP_LOOP_C_974 = 11'd1647,
    COMP_LOOP_C_975 = 11'd1648,
    COMP_LOOP_C_976 = 11'd1649,
    COMP_LOOP_C_977 = 11'd1650,
    COMP_LOOP_C_978 = 11'd1651,
    COMP_LOOP_C_979 = 11'd1652,
    COMP_LOOP_C_980 = 11'd1653,
    COMP_LOOP_C_981 = 11'd1654,
    COMP_LOOP_C_982 = 11'd1655,
    COMP_LOOP_C_983 = 11'd1656,
    COMP_LOOP_C_984 = 11'd1657,
    COMP_LOOP_C_985 = 11'd1658,
    COMP_LOOP_C_986 = 11'd1659,
    COMP_LOOP_C_987 = 11'd1660,
    COMP_LOOP_C_988 = 11'd1661,
    COMP_LOOP_C_989 = 11'd1662,
    COMP_LOOP_C_990 = 11'd1663,
    COMP_LOOP_C_991 = 11'd1664,
    COMP_LOOP_C_992 = 11'd1665,
    VEC_LOOP_C_0 = 11'd1666,
    STAGE_LOOP_C_9 = 11'd1667,
    main_C_1 = 11'd1668;

  reg [10:0] state_var;
  reg [10:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : inPlaceNTT_DIT_core_core_fsm_1
    case (state_var)
      STAGE_LOOP_C_0 : begin
        fsm_output = 11'b00000000001;
        state_var_NS = STAGE_LOOP_C_1;
      end
      STAGE_LOOP_C_1 : begin
        fsm_output = 11'b00000000010;
        state_var_NS = STAGE_LOOP_C_2;
      end
      STAGE_LOOP_C_2 : begin
        fsm_output = 11'b00000000011;
        state_var_NS = STAGE_LOOP_C_3;
      end
      STAGE_LOOP_C_3 : begin
        fsm_output = 11'b00000000100;
        state_var_NS = STAGE_LOOP_C_4;
      end
      STAGE_LOOP_C_4 : begin
        fsm_output = 11'b00000000101;
        state_var_NS = STAGE_LOOP_C_5;
      end
      STAGE_LOOP_C_5 : begin
        fsm_output = 11'b00000000110;
        state_var_NS = STAGE_LOOP_C_6;
      end
      STAGE_LOOP_C_6 : begin
        fsm_output = 11'b00000000111;
        state_var_NS = STAGE_LOOP_C_7;
      end
      STAGE_LOOP_C_7 : begin
        fsm_output = 11'b00000001000;
        state_var_NS = STAGE_LOOP_C_8;
      end
      STAGE_LOOP_C_8 : begin
        fsm_output = 11'b00000001001;
        if ( STAGE_LOOP_C_8_tr0 ) begin
          state_var_NS = COMP_LOOP_C_0;
        end
        else begin
          state_var_NS = modExp_while_C_0;
        end
      end
      modExp_while_C_0 : begin
        fsm_output = 11'b00000001010;
        state_var_NS = modExp_while_C_1;
      end
      modExp_while_C_1 : begin
        fsm_output = 11'b00000001011;
        state_var_NS = modExp_while_C_2;
      end
      modExp_while_C_2 : begin
        fsm_output = 11'b00000001100;
        state_var_NS = modExp_while_C_3;
      end
      modExp_while_C_3 : begin
        fsm_output = 11'b00000001101;
        state_var_NS = modExp_while_C_4;
      end
      modExp_while_C_4 : begin
        fsm_output = 11'b00000001110;
        state_var_NS = modExp_while_C_5;
      end
      modExp_while_C_5 : begin
        fsm_output = 11'b00000001111;
        state_var_NS = modExp_while_C_6;
      end
      modExp_while_C_6 : begin
        fsm_output = 11'b00000010000;
        state_var_NS = modExp_while_C_7;
      end
      modExp_while_C_7 : begin
        fsm_output = 11'b00000010001;
        state_var_NS = modExp_while_C_8;
      end
      modExp_while_C_8 : begin
        fsm_output = 11'b00000010010;
        state_var_NS = modExp_while_C_9;
      end
      modExp_while_C_9 : begin
        fsm_output = 11'b00000010011;
        state_var_NS = modExp_while_C_10;
      end
      modExp_while_C_10 : begin
        fsm_output = 11'b00000010100;
        state_var_NS = modExp_while_C_11;
      end
      modExp_while_C_11 : begin
        fsm_output = 11'b00000010101;
        state_var_NS = modExp_while_C_12;
      end
      modExp_while_C_12 : begin
        fsm_output = 11'b00000010110;
        state_var_NS = modExp_while_C_13;
      end
      modExp_while_C_13 : begin
        fsm_output = 11'b00000010111;
        state_var_NS = modExp_while_C_14;
      end
      modExp_while_C_14 : begin
        fsm_output = 11'b00000011000;
        state_var_NS = modExp_while_C_15;
      end
      modExp_while_C_15 : begin
        fsm_output = 11'b00000011001;
        state_var_NS = modExp_while_C_16;
      end
      modExp_while_C_16 : begin
        fsm_output = 11'b00000011010;
        state_var_NS = modExp_while_C_17;
      end
      modExp_while_C_17 : begin
        fsm_output = 11'b00000011011;
        state_var_NS = modExp_while_C_18;
      end
      modExp_while_C_18 : begin
        fsm_output = 11'b00000011100;
        state_var_NS = modExp_while_C_19;
      end
      modExp_while_C_19 : begin
        fsm_output = 11'b00000011101;
        state_var_NS = modExp_while_C_20;
      end
      modExp_while_C_20 : begin
        fsm_output = 11'b00000011110;
        state_var_NS = modExp_while_C_21;
      end
      modExp_while_C_21 : begin
        fsm_output = 11'b00000011111;
        state_var_NS = modExp_while_C_22;
      end
      modExp_while_C_22 : begin
        fsm_output = 11'b00000100000;
        state_var_NS = modExp_while_C_23;
      end
      modExp_while_C_23 : begin
        fsm_output = 11'b00000100001;
        state_var_NS = modExp_while_C_24;
      end
      modExp_while_C_24 : begin
        fsm_output = 11'b00000100010;
        state_var_NS = modExp_while_C_25;
      end
      modExp_while_C_25 : begin
        fsm_output = 11'b00000100011;
        state_var_NS = modExp_while_C_26;
      end
      modExp_while_C_26 : begin
        fsm_output = 11'b00000100100;
        state_var_NS = modExp_while_C_27;
      end
      modExp_while_C_27 : begin
        fsm_output = 11'b00000100101;
        state_var_NS = modExp_while_C_28;
      end
      modExp_while_C_28 : begin
        fsm_output = 11'b00000100110;
        state_var_NS = modExp_while_C_29;
      end
      modExp_while_C_29 : begin
        fsm_output = 11'b00000100111;
        state_var_NS = modExp_while_C_30;
      end
      modExp_while_C_30 : begin
        fsm_output = 11'b00000101000;
        state_var_NS = modExp_while_C_31;
      end
      modExp_while_C_31 : begin
        fsm_output = 11'b00000101001;
        state_var_NS = modExp_while_C_32;
      end
      modExp_while_C_32 : begin
        fsm_output = 11'b00000101010;
        state_var_NS = modExp_while_C_33;
      end
      modExp_while_C_33 : begin
        fsm_output = 11'b00000101011;
        state_var_NS = modExp_while_C_34;
      end
      modExp_while_C_34 : begin
        fsm_output = 11'b00000101100;
        state_var_NS = modExp_while_C_35;
      end
      modExp_while_C_35 : begin
        fsm_output = 11'b00000101101;
        state_var_NS = modExp_while_C_36;
      end
      modExp_while_C_36 : begin
        fsm_output = 11'b00000101110;
        state_var_NS = modExp_while_C_37;
      end
      modExp_while_C_37 : begin
        fsm_output = 11'b00000101111;
        state_var_NS = modExp_while_C_38;
      end
      modExp_while_C_38 : begin
        fsm_output = 11'b00000110000;
        if ( modExp_while_C_38_tr0 ) begin
          state_var_NS = COMP_LOOP_C_0;
        end
        else begin
          state_var_NS = modExp_while_C_0;
        end
      end
      COMP_LOOP_C_0 : begin
        fsm_output = 11'b00000110001;
        state_var_NS = COMP_LOOP_C_1;
      end
      COMP_LOOP_C_1 : begin
        fsm_output = 11'b00000110010;
        if ( COMP_LOOP_C_1_tr0 ) begin
          state_var_NS = COMP_LOOP_C_2;
        end
        else begin
          state_var_NS = COMP_LOOP_1_modExp_1_while_C_0;
        end
      end
      COMP_LOOP_1_modExp_1_while_C_0 : begin
        fsm_output = 11'b00000110011;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_1;
      end
      COMP_LOOP_1_modExp_1_while_C_1 : begin
        fsm_output = 11'b00000110100;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_2;
      end
      COMP_LOOP_1_modExp_1_while_C_2 : begin
        fsm_output = 11'b00000110101;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_3;
      end
      COMP_LOOP_1_modExp_1_while_C_3 : begin
        fsm_output = 11'b00000110110;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_4;
      end
      COMP_LOOP_1_modExp_1_while_C_4 : begin
        fsm_output = 11'b00000110111;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_5;
      end
      COMP_LOOP_1_modExp_1_while_C_5 : begin
        fsm_output = 11'b00000111000;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_6;
      end
      COMP_LOOP_1_modExp_1_while_C_6 : begin
        fsm_output = 11'b00000111001;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_7;
      end
      COMP_LOOP_1_modExp_1_while_C_7 : begin
        fsm_output = 11'b00000111010;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_8;
      end
      COMP_LOOP_1_modExp_1_while_C_8 : begin
        fsm_output = 11'b00000111011;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_9;
      end
      COMP_LOOP_1_modExp_1_while_C_9 : begin
        fsm_output = 11'b00000111100;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_10;
      end
      COMP_LOOP_1_modExp_1_while_C_10 : begin
        fsm_output = 11'b00000111101;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_11;
      end
      COMP_LOOP_1_modExp_1_while_C_11 : begin
        fsm_output = 11'b00000111110;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_12;
      end
      COMP_LOOP_1_modExp_1_while_C_12 : begin
        fsm_output = 11'b00000111111;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_13;
      end
      COMP_LOOP_1_modExp_1_while_C_13 : begin
        fsm_output = 11'b00001000000;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_14;
      end
      COMP_LOOP_1_modExp_1_while_C_14 : begin
        fsm_output = 11'b00001000001;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_15;
      end
      COMP_LOOP_1_modExp_1_while_C_15 : begin
        fsm_output = 11'b00001000010;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_16;
      end
      COMP_LOOP_1_modExp_1_while_C_16 : begin
        fsm_output = 11'b00001000011;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_17;
      end
      COMP_LOOP_1_modExp_1_while_C_17 : begin
        fsm_output = 11'b00001000100;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_18;
      end
      COMP_LOOP_1_modExp_1_while_C_18 : begin
        fsm_output = 11'b00001000101;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_19;
      end
      COMP_LOOP_1_modExp_1_while_C_19 : begin
        fsm_output = 11'b00001000110;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_20;
      end
      COMP_LOOP_1_modExp_1_while_C_20 : begin
        fsm_output = 11'b00001000111;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_21;
      end
      COMP_LOOP_1_modExp_1_while_C_21 : begin
        fsm_output = 11'b00001001000;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_22;
      end
      COMP_LOOP_1_modExp_1_while_C_22 : begin
        fsm_output = 11'b00001001001;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_23;
      end
      COMP_LOOP_1_modExp_1_while_C_23 : begin
        fsm_output = 11'b00001001010;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_24;
      end
      COMP_LOOP_1_modExp_1_while_C_24 : begin
        fsm_output = 11'b00001001011;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_25;
      end
      COMP_LOOP_1_modExp_1_while_C_25 : begin
        fsm_output = 11'b00001001100;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_26;
      end
      COMP_LOOP_1_modExp_1_while_C_26 : begin
        fsm_output = 11'b00001001101;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_27;
      end
      COMP_LOOP_1_modExp_1_while_C_27 : begin
        fsm_output = 11'b00001001110;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_28;
      end
      COMP_LOOP_1_modExp_1_while_C_28 : begin
        fsm_output = 11'b00001001111;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_29;
      end
      COMP_LOOP_1_modExp_1_while_C_29 : begin
        fsm_output = 11'b00001010000;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_30;
      end
      COMP_LOOP_1_modExp_1_while_C_30 : begin
        fsm_output = 11'b00001010001;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_31;
      end
      COMP_LOOP_1_modExp_1_while_C_31 : begin
        fsm_output = 11'b00001010010;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_32;
      end
      COMP_LOOP_1_modExp_1_while_C_32 : begin
        fsm_output = 11'b00001010011;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_33;
      end
      COMP_LOOP_1_modExp_1_while_C_33 : begin
        fsm_output = 11'b00001010100;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_34;
      end
      COMP_LOOP_1_modExp_1_while_C_34 : begin
        fsm_output = 11'b00001010101;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_35;
      end
      COMP_LOOP_1_modExp_1_while_C_35 : begin
        fsm_output = 11'b00001010110;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_36;
      end
      COMP_LOOP_1_modExp_1_while_C_36 : begin
        fsm_output = 11'b00001010111;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_37;
      end
      COMP_LOOP_1_modExp_1_while_C_37 : begin
        fsm_output = 11'b00001011000;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_38;
      end
      COMP_LOOP_1_modExp_1_while_C_38 : begin
        fsm_output = 11'b00001011001;
        if ( COMP_LOOP_1_modExp_1_while_C_38_tr0 ) begin
          state_var_NS = COMP_LOOP_C_2;
        end
        else begin
          state_var_NS = COMP_LOOP_1_modExp_1_while_C_0;
        end
      end
      COMP_LOOP_C_2 : begin
        fsm_output = 11'b00001011010;
        state_var_NS = COMP_LOOP_C_3;
      end
      COMP_LOOP_C_3 : begin
        fsm_output = 11'b00001011011;
        state_var_NS = COMP_LOOP_C_4;
      end
      COMP_LOOP_C_4 : begin
        fsm_output = 11'b00001011100;
        state_var_NS = COMP_LOOP_C_5;
      end
      COMP_LOOP_C_5 : begin
        fsm_output = 11'b00001011101;
        state_var_NS = COMP_LOOP_C_6;
      end
      COMP_LOOP_C_6 : begin
        fsm_output = 11'b00001011110;
        state_var_NS = COMP_LOOP_C_7;
      end
      COMP_LOOP_C_7 : begin
        fsm_output = 11'b00001011111;
        state_var_NS = COMP_LOOP_C_8;
      end
      COMP_LOOP_C_8 : begin
        fsm_output = 11'b00001100000;
        state_var_NS = COMP_LOOP_C_9;
      end
      COMP_LOOP_C_9 : begin
        fsm_output = 11'b00001100001;
        state_var_NS = COMP_LOOP_C_10;
      end
      COMP_LOOP_C_10 : begin
        fsm_output = 11'b00001100010;
        state_var_NS = COMP_LOOP_C_11;
      end
      COMP_LOOP_C_11 : begin
        fsm_output = 11'b00001100011;
        state_var_NS = COMP_LOOP_C_12;
      end
      COMP_LOOP_C_12 : begin
        fsm_output = 11'b00001100100;
        state_var_NS = COMP_LOOP_C_13;
      end
      COMP_LOOP_C_13 : begin
        fsm_output = 11'b00001100101;
        state_var_NS = COMP_LOOP_C_14;
      end
      COMP_LOOP_C_14 : begin
        fsm_output = 11'b00001100110;
        state_var_NS = COMP_LOOP_C_15;
      end
      COMP_LOOP_C_15 : begin
        fsm_output = 11'b00001100111;
        state_var_NS = COMP_LOOP_C_16;
      end
      COMP_LOOP_C_16 : begin
        fsm_output = 11'b00001101000;
        state_var_NS = COMP_LOOP_C_17;
      end
      COMP_LOOP_C_17 : begin
        fsm_output = 11'b00001101001;
        state_var_NS = COMP_LOOP_C_18;
      end
      COMP_LOOP_C_18 : begin
        fsm_output = 11'b00001101010;
        state_var_NS = COMP_LOOP_C_19;
      end
      COMP_LOOP_C_19 : begin
        fsm_output = 11'b00001101011;
        state_var_NS = COMP_LOOP_C_20;
      end
      COMP_LOOP_C_20 : begin
        fsm_output = 11'b00001101100;
        state_var_NS = COMP_LOOP_C_21;
      end
      COMP_LOOP_C_21 : begin
        fsm_output = 11'b00001101101;
        state_var_NS = COMP_LOOP_C_22;
      end
      COMP_LOOP_C_22 : begin
        fsm_output = 11'b00001101110;
        state_var_NS = COMP_LOOP_C_23;
      end
      COMP_LOOP_C_23 : begin
        fsm_output = 11'b00001101111;
        state_var_NS = COMP_LOOP_C_24;
      end
      COMP_LOOP_C_24 : begin
        fsm_output = 11'b00001110000;
        state_var_NS = COMP_LOOP_C_25;
      end
      COMP_LOOP_C_25 : begin
        fsm_output = 11'b00001110001;
        state_var_NS = COMP_LOOP_C_26;
      end
      COMP_LOOP_C_26 : begin
        fsm_output = 11'b00001110010;
        state_var_NS = COMP_LOOP_C_27;
      end
      COMP_LOOP_C_27 : begin
        fsm_output = 11'b00001110011;
        state_var_NS = COMP_LOOP_C_28;
      end
      COMP_LOOP_C_28 : begin
        fsm_output = 11'b00001110100;
        state_var_NS = COMP_LOOP_C_29;
      end
      COMP_LOOP_C_29 : begin
        fsm_output = 11'b00001110101;
        state_var_NS = COMP_LOOP_C_30;
      end
      COMP_LOOP_C_30 : begin
        fsm_output = 11'b00001110110;
        state_var_NS = COMP_LOOP_C_31;
      end
      COMP_LOOP_C_31 : begin
        fsm_output = 11'b00001110111;
        state_var_NS = COMP_LOOP_C_32;
      end
      COMP_LOOP_C_32 : begin
        fsm_output = 11'b00001111000;
        state_var_NS = COMP_LOOP_C_33;
      end
      COMP_LOOP_C_33 : begin
        fsm_output = 11'b00001111001;
        state_var_NS = COMP_LOOP_C_34;
      end
      COMP_LOOP_C_34 : begin
        fsm_output = 11'b00001111010;
        state_var_NS = COMP_LOOP_C_35;
      end
      COMP_LOOP_C_35 : begin
        fsm_output = 11'b00001111011;
        state_var_NS = COMP_LOOP_C_36;
      end
      COMP_LOOP_C_36 : begin
        fsm_output = 11'b00001111100;
        state_var_NS = COMP_LOOP_C_37;
      end
      COMP_LOOP_C_37 : begin
        fsm_output = 11'b00001111101;
        state_var_NS = COMP_LOOP_C_38;
      end
      COMP_LOOP_C_38 : begin
        fsm_output = 11'b00001111110;
        state_var_NS = COMP_LOOP_C_39;
      end
      COMP_LOOP_C_39 : begin
        fsm_output = 11'b00001111111;
        state_var_NS = COMP_LOOP_C_40;
      end
      COMP_LOOP_C_40 : begin
        fsm_output = 11'b00010000000;
        state_var_NS = COMP_LOOP_C_41;
      end
      COMP_LOOP_C_41 : begin
        fsm_output = 11'b00010000001;
        state_var_NS = COMP_LOOP_C_42;
      end
      COMP_LOOP_C_42 : begin
        fsm_output = 11'b00010000010;
        state_var_NS = COMP_LOOP_C_43;
      end
      COMP_LOOP_C_43 : begin
        fsm_output = 11'b00010000011;
        state_var_NS = COMP_LOOP_C_44;
      end
      COMP_LOOP_C_44 : begin
        fsm_output = 11'b00010000100;
        state_var_NS = COMP_LOOP_C_45;
      end
      COMP_LOOP_C_45 : begin
        fsm_output = 11'b00010000101;
        state_var_NS = COMP_LOOP_C_46;
      end
      COMP_LOOP_C_46 : begin
        fsm_output = 11'b00010000110;
        state_var_NS = COMP_LOOP_C_47;
      end
      COMP_LOOP_C_47 : begin
        fsm_output = 11'b00010000111;
        state_var_NS = COMP_LOOP_C_48;
      end
      COMP_LOOP_C_48 : begin
        fsm_output = 11'b00010001000;
        state_var_NS = COMP_LOOP_C_49;
      end
      COMP_LOOP_C_49 : begin
        fsm_output = 11'b00010001001;
        state_var_NS = COMP_LOOP_C_50;
      end
      COMP_LOOP_C_50 : begin
        fsm_output = 11'b00010001010;
        state_var_NS = COMP_LOOP_C_51;
      end
      COMP_LOOP_C_51 : begin
        fsm_output = 11'b00010001011;
        state_var_NS = COMP_LOOP_C_52;
      end
      COMP_LOOP_C_52 : begin
        fsm_output = 11'b00010001100;
        state_var_NS = COMP_LOOP_C_53;
      end
      COMP_LOOP_C_53 : begin
        fsm_output = 11'b00010001101;
        state_var_NS = COMP_LOOP_C_54;
      end
      COMP_LOOP_C_54 : begin
        fsm_output = 11'b00010001110;
        state_var_NS = COMP_LOOP_C_55;
      end
      COMP_LOOP_C_55 : begin
        fsm_output = 11'b00010001111;
        state_var_NS = COMP_LOOP_C_56;
      end
      COMP_LOOP_C_56 : begin
        fsm_output = 11'b00010010000;
        state_var_NS = COMP_LOOP_C_57;
      end
      COMP_LOOP_C_57 : begin
        fsm_output = 11'b00010010001;
        state_var_NS = COMP_LOOP_C_58;
      end
      COMP_LOOP_C_58 : begin
        fsm_output = 11'b00010010010;
        state_var_NS = COMP_LOOP_C_59;
      end
      COMP_LOOP_C_59 : begin
        fsm_output = 11'b00010010011;
        state_var_NS = COMP_LOOP_C_60;
      end
      COMP_LOOP_C_60 : begin
        fsm_output = 11'b00010010100;
        state_var_NS = COMP_LOOP_C_61;
      end
      COMP_LOOP_C_61 : begin
        fsm_output = 11'b00010010101;
        state_var_NS = COMP_LOOP_C_62;
      end
      COMP_LOOP_C_62 : begin
        fsm_output = 11'b00010010110;
        if ( COMP_LOOP_C_62_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_63;
        end
      end
      COMP_LOOP_C_63 : begin
        fsm_output = 11'b00010010111;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_0;
      end
      COMP_LOOP_2_modExp_1_while_C_0 : begin
        fsm_output = 11'b00010011000;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_1;
      end
      COMP_LOOP_2_modExp_1_while_C_1 : begin
        fsm_output = 11'b00010011001;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_2;
      end
      COMP_LOOP_2_modExp_1_while_C_2 : begin
        fsm_output = 11'b00010011010;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_3;
      end
      COMP_LOOP_2_modExp_1_while_C_3 : begin
        fsm_output = 11'b00010011011;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_4;
      end
      COMP_LOOP_2_modExp_1_while_C_4 : begin
        fsm_output = 11'b00010011100;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_5;
      end
      COMP_LOOP_2_modExp_1_while_C_5 : begin
        fsm_output = 11'b00010011101;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_6;
      end
      COMP_LOOP_2_modExp_1_while_C_6 : begin
        fsm_output = 11'b00010011110;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_7;
      end
      COMP_LOOP_2_modExp_1_while_C_7 : begin
        fsm_output = 11'b00010011111;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_8;
      end
      COMP_LOOP_2_modExp_1_while_C_8 : begin
        fsm_output = 11'b00010100000;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_9;
      end
      COMP_LOOP_2_modExp_1_while_C_9 : begin
        fsm_output = 11'b00010100001;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_10;
      end
      COMP_LOOP_2_modExp_1_while_C_10 : begin
        fsm_output = 11'b00010100010;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_11;
      end
      COMP_LOOP_2_modExp_1_while_C_11 : begin
        fsm_output = 11'b00010100011;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_12;
      end
      COMP_LOOP_2_modExp_1_while_C_12 : begin
        fsm_output = 11'b00010100100;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_13;
      end
      COMP_LOOP_2_modExp_1_while_C_13 : begin
        fsm_output = 11'b00010100101;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_14;
      end
      COMP_LOOP_2_modExp_1_while_C_14 : begin
        fsm_output = 11'b00010100110;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_15;
      end
      COMP_LOOP_2_modExp_1_while_C_15 : begin
        fsm_output = 11'b00010100111;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_16;
      end
      COMP_LOOP_2_modExp_1_while_C_16 : begin
        fsm_output = 11'b00010101000;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_17;
      end
      COMP_LOOP_2_modExp_1_while_C_17 : begin
        fsm_output = 11'b00010101001;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_18;
      end
      COMP_LOOP_2_modExp_1_while_C_18 : begin
        fsm_output = 11'b00010101010;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_19;
      end
      COMP_LOOP_2_modExp_1_while_C_19 : begin
        fsm_output = 11'b00010101011;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_20;
      end
      COMP_LOOP_2_modExp_1_while_C_20 : begin
        fsm_output = 11'b00010101100;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_21;
      end
      COMP_LOOP_2_modExp_1_while_C_21 : begin
        fsm_output = 11'b00010101101;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_22;
      end
      COMP_LOOP_2_modExp_1_while_C_22 : begin
        fsm_output = 11'b00010101110;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_23;
      end
      COMP_LOOP_2_modExp_1_while_C_23 : begin
        fsm_output = 11'b00010101111;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_24;
      end
      COMP_LOOP_2_modExp_1_while_C_24 : begin
        fsm_output = 11'b00010110000;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_25;
      end
      COMP_LOOP_2_modExp_1_while_C_25 : begin
        fsm_output = 11'b00010110001;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_26;
      end
      COMP_LOOP_2_modExp_1_while_C_26 : begin
        fsm_output = 11'b00010110010;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_27;
      end
      COMP_LOOP_2_modExp_1_while_C_27 : begin
        fsm_output = 11'b00010110011;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_28;
      end
      COMP_LOOP_2_modExp_1_while_C_28 : begin
        fsm_output = 11'b00010110100;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_29;
      end
      COMP_LOOP_2_modExp_1_while_C_29 : begin
        fsm_output = 11'b00010110101;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_30;
      end
      COMP_LOOP_2_modExp_1_while_C_30 : begin
        fsm_output = 11'b00010110110;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_31;
      end
      COMP_LOOP_2_modExp_1_while_C_31 : begin
        fsm_output = 11'b00010110111;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_32;
      end
      COMP_LOOP_2_modExp_1_while_C_32 : begin
        fsm_output = 11'b00010111000;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_33;
      end
      COMP_LOOP_2_modExp_1_while_C_33 : begin
        fsm_output = 11'b00010111001;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_34;
      end
      COMP_LOOP_2_modExp_1_while_C_34 : begin
        fsm_output = 11'b00010111010;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_35;
      end
      COMP_LOOP_2_modExp_1_while_C_35 : begin
        fsm_output = 11'b00010111011;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_36;
      end
      COMP_LOOP_2_modExp_1_while_C_36 : begin
        fsm_output = 11'b00010111100;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_37;
      end
      COMP_LOOP_2_modExp_1_while_C_37 : begin
        fsm_output = 11'b00010111101;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_38;
      end
      COMP_LOOP_2_modExp_1_while_C_38 : begin
        fsm_output = 11'b00010111110;
        if ( COMP_LOOP_2_modExp_1_while_C_38_tr0 ) begin
          state_var_NS = COMP_LOOP_C_64;
        end
        else begin
          state_var_NS = COMP_LOOP_2_modExp_1_while_C_0;
        end
      end
      COMP_LOOP_C_64 : begin
        fsm_output = 11'b00010111111;
        state_var_NS = COMP_LOOP_C_65;
      end
      COMP_LOOP_C_65 : begin
        fsm_output = 11'b00011000000;
        state_var_NS = COMP_LOOP_C_66;
      end
      COMP_LOOP_C_66 : begin
        fsm_output = 11'b00011000001;
        state_var_NS = COMP_LOOP_C_67;
      end
      COMP_LOOP_C_67 : begin
        fsm_output = 11'b00011000010;
        state_var_NS = COMP_LOOP_C_68;
      end
      COMP_LOOP_C_68 : begin
        fsm_output = 11'b00011000011;
        state_var_NS = COMP_LOOP_C_69;
      end
      COMP_LOOP_C_69 : begin
        fsm_output = 11'b00011000100;
        state_var_NS = COMP_LOOP_C_70;
      end
      COMP_LOOP_C_70 : begin
        fsm_output = 11'b00011000101;
        state_var_NS = COMP_LOOP_C_71;
      end
      COMP_LOOP_C_71 : begin
        fsm_output = 11'b00011000110;
        state_var_NS = COMP_LOOP_C_72;
      end
      COMP_LOOP_C_72 : begin
        fsm_output = 11'b00011000111;
        state_var_NS = COMP_LOOP_C_73;
      end
      COMP_LOOP_C_73 : begin
        fsm_output = 11'b00011001000;
        state_var_NS = COMP_LOOP_C_74;
      end
      COMP_LOOP_C_74 : begin
        fsm_output = 11'b00011001001;
        state_var_NS = COMP_LOOP_C_75;
      end
      COMP_LOOP_C_75 : begin
        fsm_output = 11'b00011001010;
        state_var_NS = COMP_LOOP_C_76;
      end
      COMP_LOOP_C_76 : begin
        fsm_output = 11'b00011001011;
        state_var_NS = COMP_LOOP_C_77;
      end
      COMP_LOOP_C_77 : begin
        fsm_output = 11'b00011001100;
        state_var_NS = COMP_LOOP_C_78;
      end
      COMP_LOOP_C_78 : begin
        fsm_output = 11'b00011001101;
        state_var_NS = COMP_LOOP_C_79;
      end
      COMP_LOOP_C_79 : begin
        fsm_output = 11'b00011001110;
        state_var_NS = COMP_LOOP_C_80;
      end
      COMP_LOOP_C_80 : begin
        fsm_output = 11'b00011001111;
        state_var_NS = COMP_LOOP_C_81;
      end
      COMP_LOOP_C_81 : begin
        fsm_output = 11'b00011010000;
        state_var_NS = COMP_LOOP_C_82;
      end
      COMP_LOOP_C_82 : begin
        fsm_output = 11'b00011010001;
        state_var_NS = COMP_LOOP_C_83;
      end
      COMP_LOOP_C_83 : begin
        fsm_output = 11'b00011010010;
        state_var_NS = COMP_LOOP_C_84;
      end
      COMP_LOOP_C_84 : begin
        fsm_output = 11'b00011010011;
        state_var_NS = COMP_LOOP_C_85;
      end
      COMP_LOOP_C_85 : begin
        fsm_output = 11'b00011010100;
        state_var_NS = COMP_LOOP_C_86;
      end
      COMP_LOOP_C_86 : begin
        fsm_output = 11'b00011010101;
        state_var_NS = COMP_LOOP_C_87;
      end
      COMP_LOOP_C_87 : begin
        fsm_output = 11'b00011010110;
        state_var_NS = COMP_LOOP_C_88;
      end
      COMP_LOOP_C_88 : begin
        fsm_output = 11'b00011010111;
        state_var_NS = COMP_LOOP_C_89;
      end
      COMP_LOOP_C_89 : begin
        fsm_output = 11'b00011011000;
        state_var_NS = COMP_LOOP_C_90;
      end
      COMP_LOOP_C_90 : begin
        fsm_output = 11'b00011011001;
        state_var_NS = COMP_LOOP_C_91;
      end
      COMP_LOOP_C_91 : begin
        fsm_output = 11'b00011011010;
        state_var_NS = COMP_LOOP_C_92;
      end
      COMP_LOOP_C_92 : begin
        fsm_output = 11'b00011011011;
        state_var_NS = COMP_LOOP_C_93;
      end
      COMP_LOOP_C_93 : begin
        fsm_output = 11'b00011011100;
        state_var_NS = COMP_LOOP_C_94;
      end
      COMP_LOOP_C_94 : begin
        fsm_output = 11'b00011011101;
        state_var_NS = COMP_LOOP_C_95;
      end
      COMP_LOOP_C_95 : begin
        fsm_output = 11'b00011011110;
        state_var_NS = COMP_LOOP_C_96;
      end
      COMP_LOOP_C_96 : begin
        fsm_output = 11'b00011011111;
        state_var_NS = COMP_LOOP_C_97;
      end
      COMP_LOOP_C_97 : begin
        fsm_output = 11'b00011100000;
        state_var_NS = COMP_LOOP_C_98;
      end
      COMP_LOOP_C_98 : begin
        fsm_output = 11'b00011100001;
        state_var_NS = COMP_LOOP_C_99;
      end
      COMP_LOOP_C_99 : begin
        fsm_output = 11'b00011100010;
        state_var_NS = COMP_LOOP_C_100;
      end
      COMP_LOOP_C_100 : begin
        fsm_output = 11'b00011100011;
        state_var_NS = COMP_LOOP_C_101;
      end
      COMP_LOOP_C_101 : begin
        fsm_output = 11'b00011100100;
        state_var_NS = COMP_LOOP_C_102;
      end
      COMP_LOOP_C_102 : begin
        fsm_output = 11'b00011100101;
        state_var_NS = COMP_LOOP_C_103;
      end
      COMP_LOOP_C_103 : begin
        fsm_output = 11'b00011100110;
        state_var_NS = COMP_LOOP_C_104;
      end
      COMP_LOOP_C_104 : begin
        fsm_output = 11'b00011100111;
        state_var_NS = COMP_LOOP_C_105;
      end
      COMP_LOOP_C_105 : begin
        fsm_output = 11'b00011101000;
        state_var_NS = COMP_LOOP_C_106;
      end
      COMP_LOOP_C_106 : begin
        fsm_output = 11'b00011101001;
        state_var_NS = COMP_LOOP_C_107;
      end
      COMP_LOOP_C_107 : begin
        fsm_output = 11'b00011101010;
        state_var_NS = COMP_LOOP_C_108;
      end
      COMP_LOOP_C_108 : begin
        fsm_output = 11'b00011101011;
        state_var_NS = COMP_LOOP_C_109;
      end
      COMP_LOOP_C_109 : begin
        fsm_output = 11'b00011101100;
        state_var_NS = COMP_LOOP_C_110;
      end
      COMP_LOOP_C_110 : begin
        fsm_output = 11'b00011101101;
        state_var_NS = COMP_LOOP_C_111;
      end
      COMP_LOOP_C_111 : begin
        fsm_output = 11'b00011101110;
        state_var_NS = COMP_LOOP_C_112;
      end
      COMP_LOOP_C_112 : begin
        fsm_output = 11'b00011101111;
        state_var_NS = COMP_LOOP_C_113;
      end
      COMP_LOOP_C_113 : begin
        fsm_output = 11'b00011110000;
        state_var_NS = COMP_LOOP_C_114;
      end
      COMP_LOOP_C_114 : begin
        fsm_output = 11'b00011110001;
        state_var_NS = COMP_LOOP_C_115;
      end
      COMP_LOOP_C_115 : begin
        fsm_output = 11'b00011110010;
        state_var_NS = COMP_LOOP_C_116;
      end
      COMP_LOOP_C_116 : begin
        fsm_output = 11'b00011110011;
        state_var_NS = COMP_LOOP_C_117;
      end
      COMP_LOOP_C_117 : begin
        fsm_output = 11'b00011110100;
        state_var_NS = COMP_LOOP_C_118;
      end
      COMP_LOOP_C_118 : begin
        fsm_output = 11'b00011110101;
        state_var_NS = COMP_LOOP_C_119;
      end
      COMP_LOOP_C_119 : begin
        fsm_output = 11'b00011110110;
        state_var_NS = COMP_LOOP_C_120;
      end
      COMP_LOOP_C_120 : begin
        fsm_output = 11'b00011110111;
        state_var_NS = COMP_LOOP_C_121;
      end
      COMP_LOOP_C_121 : begin
        fsm_output = 11'b00011111000;
        state_var_NS = COMP_LOOP_C_122;
      end
      COMP_LOOP_C_122 : begin
        fsm_output = 11'b00011111001;
        state_var_NS = COMP_LOOP_C_123;
      end
      COMP_LOOP_C_123 : begin
        fsm_output = 11'b00011111010;
        state_var_NS = COMP_LOOP_C_124;
      end
      COMP_LOOP_C_124 : begin
        fsm_output = 11'b00011111011;
        if ( COMP_LOOP_C_124_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_125;
        end
      end
      COMP_LOOP_C_125 : begin
        fsm_output = 11'b00011111100;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_0;
      end
      COMP_LOOP_3_modExp_1_while_C_0 : begin
        fsm_output = 11'b00011111101;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_1;
      end
      COMP_LOOP_3_modExp_1_while_C_1 : begin
        fsm_output = 11'b00011111110;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_2;
      end
      COMP_LOOP_3_modExp_1_while_C_2 : begin
        fsm_output = 11'b00011111111;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_3;
      end
      COMP_LOOP_3_modExp_1_while_C_3 : begin
        fsm_output = 11'b00100000000;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_4;
      end
      COMP_LOOP_3_modExp_1_while_C_4 : begin
        fsm_output = 11'b00100000001;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_5;
      end
      COMP_LOOP_3_modExp_1_while_C_5 : begin
        fsm_output = 11'b00100000010;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_6;
      end
      COMP_LOOP_3_modExp_1_while_C_6 : begin
        fsm_output = 11'b00100000011;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_7;
      end
      COMP_LOOP_3_modExp_1_while_C_7 : begin
        fsm_output = 11'b00100000100;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_8;
      end
      COMP_LOOP_3_modExp_1_while_C_8 : begin
        fsm_output = 11'b00100000101;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_9;
      end
      COMP_LOOP_3_modExp_1_while_C_9 : begin
        fsm_output = 11'b00100000110;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_10;
      end
      COMP_LOOP_3_modExp_1_while_C_10 : begin
        fsm_output = 11'b00100000111;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_11;
      end
      COMP_LOOP_3_modExp_1_while_C_11 : begin
        fsm_output = 11'b00100001000;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_12;
      end
      COMP_LOOP_3_modExp_1_while_C_12 : begin
        fsm_output = 11'b00100001001;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_13;
      end
      COMP_LOOP_3_modExp_1_while_C_13 : begin
        fsm_output = 11'b00100001010;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_14;
      end
      COMP_LOOP_3_modExp_1_while_C_14 : begin
        fsm_output = 11'b00100001011;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_15;
      end
      COMP_LOOP_3_modExp_1_while_C_15 : begin
        fsm_output = 11'b00100001100;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_16;
      end
      COMP_LOOP_3_modExp_1_while_C_16 : begin
        fsm_output = 11'b00100001101;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_17;
      end
      COMP_LOOP_3_modExp_1_while_C_17 : begin
        fsm_output = 11'b00100001110;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_18;
      end
      COMP_LOOP_3_modExp_1_while_C_18 : begin
        fsm_output = 11'b00100001111;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_19;
      end
      COMP_LOOP_3_modExp_1_while_C_19 : begin
        fsm_output = 11'b00100010000;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_20;
      end
      COMP_LOOP_3_modExp_1_while_C_20 : begin
        fsm_output = 11'b00100010001;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_21;
      end
      COMP_LOOP_3_modExp_1_while_C_21 : begin
        fsm_output = 11'b00100010010;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_22;
      end
      COMP_LOOP_3_modExp_1_while_C_22 : begin
        fsm_output = 11'b00100010011;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_23;
      end
      COMP_LOOP_3_modExp_1_while_C_23 : begin
        fsm_output = 11'b00100010100;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_24;
      end
      COMP_LOOP_3_modExp_1_while_C_24 : begin
        fsm_output = 11'b00100010101;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_25;
      end
      COMP_LOOP_3_modExp_1_while_C_25 : begin
        fsm_output = 11'b00100010110;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_26;
      end
      COMP_LOOP_3_modExp_1_while_C_26 : begin
        fsm_output = 11'b00100010111;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_27;
      end
      COMP_LOOP_3_modExp_1_while_C_27 : begin
        fsm_output = 11'b00100011000;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_28;
      end
      COMP_LOOP_3_modExp_1_while_C_28 : begin
        fsm_output = 11'b00100011001;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_29;
      end
      COMP_LOOP_3_modExp_1_while_C_29 : begin
        fsm_output = 11'b00100011010;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_30;
      end
      COMP_LOOP_3_modExp_1_while_C_30 : begin
        fsm_output = 11'b00100011011;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_31;
      end
      COMP_LOOP_3_modExp_1_while_C_31 : begin
        fsm_output = 11'b00100011100;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_32;
      end
      COMP_LOOP_3_modExp_1_while_C_32 : begin
        fsm_output = 11'b00100011101;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_33;
      end
      COMP_LOOP_3_modExp_1_while_C_33 : begin
        fsm_output = 11'b00100011110;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_34;
      end
      COMP_LOOP_3_modExp_1_while_C_34 : begin
        fsm_output = 11'b00100011111;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_35;
      end
      COMP_LOOP_3_modExp_1_while_C_35 : begin
        fsm_output = 11'b00100100000;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_36;
      end
      COMP_LOOP_3_modExp_1_while_C_36 : begin
        fsm_output = 11'b00100100001;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_37;
      end
      COMP_LOOP_3_modExp_1_while_C_37 : begin
        fsm_output = 11'b00100100010;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_38;
      end
      COMP_LOOP_3_modExp_1_while_C_38 : begin
        fsm_output = 11'b00100100011;
        if ( COMP_LOOP_3_modExp_1_while_C_38_tr0 ) begin
          state_var_NS = COMP_LOOP_C_126;
        end
        else begin
          state_var_NS = COMP_LOOP_3_modExp_1_while_C_0;
        end
      end
      COMP_LOOP_C_126 : begin
        fsm_output = 11'b00100100100;
        state_var_NS = COMP_LOOP_C_127;
      end
      COMP_LOOP_C_127 : begin
        fsm_output = 11'b00100100101;
        state_var_NS = COMP_LOOP_C_128;
      end
      COMP_LOOP_C_128 : begin
        fsm_output = 11'b00100100110;
        state_var_NS = COMP_LOOP_C_129;
      end
      COMP_LOOP_C_129 : begin
        fsm_output = 11'b00100100111;
        state_var_NS = COMP_LOOP_C_130;
      end
      COMP_LOOP_C_130 : begin
        fsm_output = 11'b00100101000;
        state_var_NS = COMP_LOOP_C_131;
      end
      COMP_LOOP_C_131 : begin
        fsm_output = 11'b00100101001;
        state_var_NS = COMP_LOOP_C_132;
      end
      COMP_LOOP_C_132 : begin
        fsm_output = 11'b00100101010;
        state_var_NS = COMP_LOOP_C_133;
      end
      COMP_LOOP_C_133 : begin
        fsm_output = 11'b00100101011;
        state_var_NS = COMP_LOOP_C_134;
      end
      COMP_LOOP_C_134 : begin
        fsm_output = 11'b00100101100;
        state_var_NS = COMP_LOOP_C_135;
      end
      COMP_LOOP_C_135 : begin
        fsm_output = 11'b00100101101;
        state_var_NS = COMP_LOOP_C_136;
      end
      COMP_LOOP_C_136 : begin
        fsm_output = 11'b00100101110;
        state_var_NS = COMP_LOOP_C_137;
      end
      COMP_LOOP_C_137 : begin
        fsm_output = 11'b00100101111;
        state_var_NS = COMP_LOOP_C_138;
      end
      COMP_LOOP_C_138 : begin
        fsm_output = 11'b00100110000;
        state_var_NS = COMP_LOOP_C_139;
      end
      COMP_LOOP_C_139 : begin
        fsm_output = 11'b00100110001;
        state_var_NS = COMP_LOOP_C_140;
      end
      COMP_LOOP_C_140 : begin
        fsm_output = 11'b00100110010;
        state_var_NS = COMP_LOOP_C_141;
      end
      COMP_LOOP_C_141 : begin
        fsm_output = 11'b00100110011;
        state_var_NS = COMP_LOOP_C_142;
      end
      COMP_LOOP_C_142 : begin
        fsm_output = 11'b00100110100;
        state_var_NS = COMP_LOOP_C_143;
      end
      COMP_LOOP_C_143 : begin
        fsm_output = 11'b00100110101;
        state_var_NS = COMP_LOOP_C_144;
      end
      COMP_LOOP_C_144 : begin
        fsm_output = 11'b00100110110;
        state_var_NS = COMP_LOOP_C_145;
      end
      COMP_LOOP_C_145 : begin
        fsm_output = 11'b00100110111;
        state_var_NS = COMP_LOOP_C_146;
      end
      COMP_LOOP_C_146 : begin
        fsm_output = 11'b00100111000;
        state_var_NS = COMP_LOOP_C_147;
      end
      COMP_LOOP_C_147 : begin
        fsm_output = 11'b00100111001;
        state_var_NS = COMP_LOOP_C_148;
      end
      COMP_LOOP_C_148 : begin
        fsm_output = 11'b00100111010;
        state_var_NS = COMP_LOOP_C_149;
      end
      COMP_LOOP_C_149 : begin
        fsm_output = 11'b00100111011;
        state_var_NS = COMP_LOOP_C_150;
      end
      COMP_LOOP_C_150 : begin
        fsm_output = 11'b00100111100;
        state_var_NS = COMP_LOOP_C_151;
      end
      COMP_LOOP_C_151 : begin
        fsm_output = 11'b00100111101;
        state_var_NS = COMP_LOOP_C_152;
      end
      COMP_LOOP_C_152 : begin
        fsm_output = 11'b00100111110;
        state_var_NS = COMP_LOOP_C_153;
      end
      COMP_LOOP_C_153 : begin
        fsm_output = 11'b00100111111;
        state_var_NS = COMP_LOOP_C_154;
      end
      COMP_LOOP_C_154 : begin
        fsm_output = 11'b00101000000;
        state_var_NS = COMP_LOOP_C_155;
      end
      COMP_LOOP_C_155 : begin
        fsm_output = 11'b00101000001;
        state_var_NS = COMP_LOOP_C_156;
      end
      COMP_LOOP_C_156 : begin
        fsm_output = 11'b00101000010;
        state_var_NS = COMP_LOOP_C_157;
      end
      COMP_LOOP_C_157 : begin
        fsm_output = 11'b00101000011;
        state_var_NS = COMP_LOOP_C_158;
      end
      COMP_LOOP_C_158 : begin
        fsm_output = 11'b00101000100;
        state_var_NS = COMP_LOOP_C_159;
      end
      COMP_LOOP_C_159 : begin
        fsm_output = 11'b00101000101;
        state_var_NS = COMP_LOOP_C_160;
      end
      COMP_LOOP_C_160 : begin
        fsm_output = 11'b00101000110;
        state_var_NS = COMP_LOOP_C_161;
      end
      COMP_LOOP_C_161 : begin
        fsm_output = 11'b00101000111;
        state_var_NS = COMP_LOOP_C_162;
      end
      COMP_LOOP_C_162 : begin
        fsm_output = 11'b00101001000;
        state_var_NS = COMP_LOOP_C_163;
      end
      COMP_LOOP_C_163 : begin
        fsm_output = 11'b00101001001;
        state_var_NS = COMP_LOOP_C_164;
      end
      COMP_LOOP_C_164 : begin
        fsm_output = 11'b00101001010;
        state_var_NS = COMP_LOOP_C_165;
      end
      COMP_LOOP_C_165 : begin
        fsm_output = 11'b00101001011;
        state_var_NS = COMP_LOOP_C_166;
      end
      COMP_LOOP_C_166 : begin
        fsm_output = 11'b00101001100;
        state_var_NS = COMP_LOOP_C_167;
      end
      COMP_LOOP_C_167 : begin
        fsm_output = 11'b00101001101;
        state_var_NS = COMP_LOOP_C_168;
      end
      COMP_LOOP_C_168 : begin
        fsm_output = 11'b00101001110;
        state_var_NS = COMP_LOOP_C_169;
      end
      COMP_LOOP_C_169 : begin
        fsm_output = 11'b00101001111;
        state_var_NS = COMP_LOOP_C_170;
      end
      COMP_LOOP_C_170 : begin
        fsm_output = 11'b00101010000;
        state_var_NS = COMP_LOOP_C_171;
      end
      COMP_LOOP_C_171 : begin
        fsm_output = 11'b00101010001;
        state_var_NS = COMP_LOOP_C_172;
      end
      COMP_LOOP_C_172 : begin
        fsm_output = 11'b00101010010;
        state_var_NS = COMP_LOOP_C_173;
      end
      COMP_LOOP_C_173 : begin
        fsm_output = 11'b00101010011;
        state_var_NS = COMP_LOOP_C_174;
      end
      COMP_LOOP_C_174 : begin
        fsm_output = 11'b00101010100;
        state_var_NS = COMP_LOOP_C_175;
      end
      COMP_LOOP_C_175 : begin
        fsm_output = 11'b00101010101;
        state_var_NS = COMP_LOOP_C_176;
      end
      COMP_LOOP_C_176 : begin
        fsm_output = 11'b00101010110;
        state_var_NS = COMP_LOOP_C_177;
      end
      COMP_LOOP_C_177 : begin
        fsm_output = 11'b00101010111;
        state_var_NS = COMP_LOOP_C_178;
      end
      COMP_LOOP_C_178 : begin
        fsm_output = 11'b00101011000;
        state_var_NS = COMP_LOOP_C_179;
      end
      COMP_LOOP_C_179 : begin
        fsm_output = 11'b00101011001;
        state_var_NS = COMP_LOOP_C_180;
      end
      COMP_LOOP_C_180 : begin
        fsm_output = 11'b00101011010;
        state_var_NS = COMP_LOOP_C_181;
      end
      COMP_LOOP_C_181 : begin
        fsm_output = 11'b00101011011;
        state_var_NS = COMP_LOOP_C_182;
      end
      COMP_LOOP_C_182 : begin
        fsm_output = 11'b00101011100;
        state_var_NS = COMP_LOOP_C_183;
      end
      COMP_LOOP_C_183 : begin
        fsm_output = 11'b00101011101;
        state_var_NS = COMP_LOOP_C_184;
      end
      COMP_LOOP_C_184 : begin
        fsm_output = 11'b00101011110;
        state_var_NS = COMP_LOOP_C_185;
      end
      COMP_LOOP_C_185 : begin
        fsm_output = 11'b00101011111;
        state_var_NS = COMP_LOOP_C_186;
      end
      COMP_LOOP_C_186 : begin
        fsm_output = 11'b00101100000;
        if ( COMP_LOOP_C_186_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_187;
        end
      end
      COMP_LOOP_C_187 : begin
        fsm_output = 11'b00101100001;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_0;
      end
      COMP_LOOP_4_modExp_1_while_C_0 : begin
        fsm_output = 11'b00101100010;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_1;
      end
      COMP_LOOP_4_modExp_1_while_C_1 : begin
        fsm_output = 11'b00101100011;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_2;
      end
      COMP_LOOP_4_modExp_1_while_C_2 : begin
        fsm_output = 11'b00101100100;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_3;
      end
      COMP_LOOP_4_modExp_1_while_C_3 : begin
        fsm_output = 11'b00101100101;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_4;
      end
      COMP_LOOP_4_modExp_1_while_C_4 : begin
        fsm_output = 11'b00101100110;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_5;
      end
      COMP_LOOP_4_modExp_1_while_C_5 : begin
        fsm_output = 11'b00101100111;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_6;
      end
      COMP_LOOP_4_modExp_1_while_C_6 : begin
        fsm_output = 11'b00101101000;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_7;
      end
      COMP_LOOP_4_modExp_1_while_C_7 : begin
        fsm_output = 11'b00101101001;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_8;
      end
      COMP_LOOP_4_modExp_1_while_C_8 : begin
        fsm_output = 11'b00101101010;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_9;
      end
      COMP_LOOP_4_modExp_1_while_C_9 : begin
        fsm_output = 11'b00101101011;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_10;
      end
      COMP_LOOP_4_modExp_1_while_C_10 : begin
        fsm_output = 11'b00101101100;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_11;
      end
      COMP_LOOP_4_modExp_1_while_C_11 : begin
        fsm_output = 11'b00101101101;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_12;
      end
      COMP_LOOP_4_modExp_1_while_C_12 : begin
        fsm_output = 11'b00101101110;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_13;
      end
      COMP_LOOP_4_modExp_1_while_C_13 : begin
        fsm_output = 11'b00101101111;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_14;
      end
      COMP_LOOP_4_modExp_1_while_C_14 : begin
        fsm_output = 11'b00101110000;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_15;
      end
      COMP_LOOP_4_modExp_1_while_C_15 : begin
        fsm_output = 11'b00101110001;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_16;
      end
      COMP_LOOP_4_modExp_1_while_C_16 : begin
        fsm_output = 11'b00101110010;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_17;
      end
      COMP_LOOP_4_modExp_1_while_C_17 : begin
        fsm_output = 11'b00101110011;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_18;
      end
      COMP_LOOP_4_modExp_1_while_C_18 : begin
        fsm_output = 11'b00101110100;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_19;
      end
      COMP_LOOP_4_modExp_1_while_C_19 : begin
        fsm_output = 11'b00101110101;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_20;
      end
      COMP_LOOP_4_modExp_1_while_C_20 : begin
        fsm_output = 11'b00101110110;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_21;
      end
      COMP_LOOP_4_modExp_1_while_C_21 : begin
        fsm_output = 11'b00101110111;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_22;
      end
      COMP_LOOP_4_modExp_1_while_C_22 : begin
        fsm_output = 11'b00101111000;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_23;
      end
      COMP_LOOP_4_modExp_1_while_C_23 : begin
        fsm_output = 11'b00101111001;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_24;
      end
      COMP_LOOP_4_modExp_1_while_C_24 : begin
        fsm_output = 11'b00101111010;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_25;
      end
      COMP_LOOP_4_modExp_1_while_C_25 : begin
        fsm_output = 11'b00101111011;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_26;
      end
      COMP_LOOP_4_modExp_1_while_C_26 : begin
        fsm_output = 11'b00101111100;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_27;
      end
      COMP_LOOP_4_modExp_1_while_C_27 : begin
        fsm_output = 11'b00101111101;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_28;
      end
      COMP_LOOP_4_modExp_1_while_C_28 : begin
        fsm_output = 11'b00101111110;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_29;
      end
      COMP_LOOP_4_modExp_1_while_C_29 : begin
        fsm_output = 11'b00101111111;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_30;
      end
      COMP_LOOP_4_modExp_1_while_C_30 : begin
        fsm_output = 11'b00110000000;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_31;
      end
      COMP_LOOP_4_modExp_1_while_C_31 : begin
        fsm_output = 11'b00110000001;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_32;
      end
      COMP_LOOP_4_modExp_1_while_C_32 : begin
        fsm_output = 11'b00110000010;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_33;
      end
      COMP_LOOP_4_modExp_1_while_C_33 : begin
        fsm_output = 11'b00110000011;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_34;
      end
      COMP_LOOP_4_modExp_1_while_C_34 : begin
        fsm_output = 11'b00110000100;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_35;
      end
      COMP_LOOP_4_modExp_1_while_C_35 : begin
        fsm_output = 11'b00110000101;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_36;
      end
      COMP_LOOP_4_modExp_1_while_C_36 : begin
        fsm_output = 11'b00110000110;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_37;
      end
      COMP_LOOP_4_modExp_1_while_C_37 : begin
        fsm_output = 11'b00110000111;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_38;
      end
      COMP_LOOP_4_modExp_1_while_C_38 : begin
        fsm_output = 11'b00110001000;
        if ( COMP_LOOP_4_modExp_1_while_C_38_tr0 ) begin
          state_var_NS = COMP_LOOP_C_188;
        end
        else begin
          state_var_NS = COMP_LOOP_4_modExp_1_while_C_0;
        end
      end
      COMP_LOOP_C_188 : begin
        fsm_output = 11'b00110001001;
        state_var_NS = COMP_LOOP_C_189;
      end
      COMP_LOOP_C_189 : begin
        fsm_output = 11'b00110001010;
        state_var_NS = COMP_LOOP_C_190;
      end
      COMP_LOOP_C_190 : begin
        fsm_output = 11'b00110001011;
        state_var_NS = COMP_LOOP_C_191;
      end
      COMP_LOOP_C_191 : begin
        fsm_output = 11'b00110001100;
        state_var_NS = COMP_LOOP_C_192;
      end
      COMP_LOOP_C_192 : begin
        fsm_output = 11'b00110001101;
        state_var_NS = COMP_LOOP_C_193;
      end
      COMP_LOOP_C_193 : begin
        fsm_output = 11'b00110001110;
        state_var_NS = COMP_LOOP_C_194;
      end
      COMP_LOOP_C_194 : begin
        fsm_output = 11'b00110001111;
        state_var_NS = COMP_LOOP_C_195;
      end
      COMP_LOOP_C_195 : begin
        fsm_output = 11'b00110010000;
        state_var_NS = COMP_LOOP_C_196;
      end
      COMP_LOOP_C_196 : begin
        fsm_output = 11'b00110010001;
        state_var_NS = COMP_LOOP_C_197;
      end
      COMP_LOOP_C_197 : begin
        fsm_output = 11'b00110010010;
        state_var_NS = COMP_LOOP_C_198;
      end
      COMP_LOOP_C_198 : begin
        fsm_output = 11'b00110010011;
        state_var_NS = COMP_LOOP_C_199;
      end
      COMP_LOOP_C_199 : begin
        fsm_output = 11'b00110010100;
        state_var_NS = COMP_LOOP_C_200;
      end
      COMP_LOOP_C_200 : begin
        fsm_output = 11'b00110010101;
        state_var_NS = COMP_LOOP_C_201;
      end
      COMP_LOOP_C_201 : begin
        fsm_output = 11'b00110010110;
        state_var_NS = COMP_LOOP_C_202;
      end
      COMP_LOOP_C_202 : begin
        fsm_output = 11'b00110010111;
        state_var_NS = COMP_LOOP_C_203;
      end
      COMP_LOOP_C_203 : begin
        fsm_output = 11'b00110011000;
        state_var_NS = COMP_LOOP_C_204;
      end
      COMP_LOOP_C_204 : begin
        fsm_output = 11'b00110011001;
        state_var_NS = COMP_LOOP_C_205;
      end
      COMP_LOOP_C_205 : begin
        fsm_output = 11'b00110011010;
        state_var_NS = COMP_LOOP_C_206;
      end
      COMP_LOOP_C_206 : begin
        fsm_output = 11'b00110011011;
        state_var_NS = COMP_LOOP_C_207;
      end
      COMP_LOOP_C_207 : begin
        fsm_output = 11'b00110011100;
        state_var_NS = COMP_LOOP_C_208;
      end
      COMP_LOOP_C_208 : begin
        fsm_output = 11'b00110011101;
        state_var_NS = COMP_LOOP_C_209;
      end
      COMP_LOOP_C_209 : begin
        fsm_output = 11'b00110011110;
        state_var_NS = COMP_LOOP_C_210;
      end
      COMP_LOOP_C_210 : begin
        fsm_output = 11'b00110011111;
        state_var_NS = COMP_LOOP_C_211;
      end
      COMP_LOOP_C_211 : begin
        fsm_output = 11'b00110100000;
        state_var_NS = COMP_LOOP_C_212;
      end
      COMP_LOOP_C_212 : begin
        fsm_output = 11'b00110100001;
        state_var_NS = COMP_LOOP_C_213;
      end
      COMP_LOOP_C_213 : begin
        fsm_output = 11'b00110100010;
        state_var_NS = COMP_LOOP_C_214;
      end
      COMP_LOOP_C_214 : begin
        fsm_output = 11'b00110100011;
        state_var_NS = COMP_LOOP_C_215;
      end
      COMP_LOOP_C_215 : begin
        fsm_output = 11'b00110100100;
        state_var_NS = COMP_LOOP_C_216;
      end
      COMP_LOOP_C_216 : begin
        fsm_output = 11'b00110100101;
        state_var_NS = COMP_LOOP_C_217;
      end
      COMP_LOOP_C_217 : begin
        fsm_output = 11'b00110100110;
        state_var_NS = COMP_LOOP_C_218;
      end
      COMP_LOOP_C_218 : begin
        fsm_output = 11'b00110100111;
        state_var_NS = COMP_LOOP_C_219;
      end
      COMP_LOOP_C_219 : begin
        fsm_output = 11'b00110101000;
        state_var_NS = COMP_LOOP_C_220;
      end
      COMP_LOOP_C_220 : begin
        fsm_output = 11'b00110101001;
        state_var_NS = COMP_LOOP_C_221;
      end
      COMP_LOOP_C_221 : begin
        fsm_output = 11'b00110101010;
        state_var_NS = COMP_LOOP_C_222;
      end
      COMP_LOOP_C_222 : begin
        fsm_output = 11'b00110101011;
        state_var_NS = COMP_LOOP_C_223;
      end
      COMP_LOOP_C_223 : begin
        fsm_output = 11'b00110101100;
        state_var_NS = COMP_LOOP_C_224;
      end
      COMP_LOOP_C_224 : begin
        fsm_output = 11'b00110101101;
        state_var_NS = COMP_LOOP_C_225;
      end
      COMP_LOOP_C_225 : begin
        fsm_output = 11'b00110101110;
        state_var_NS = COMP_LOOP_C_226;
      end
      COMP_LOOP_C_226 : begin
        fsm_output = 11'b00110101111;
        state_var_NS = COMP_LOOP_C_227;
      end
      COMP_LOOP_C_227 : begin
        fsm_output = 11'b00110110000;
        state_var_NS = COMP_LOOP_C_228;
      end
      COMP_LOOP_C_228 : begin
        fsm_output = 11'b00110110001;
        state_var_NS = COMP_LOOP_C_229;
      end
      COMP_LOOP_C_229 : begin
        fsm_output = 11'b00110110010;
        state_var_NS = COMP_LOOP_C_230;
      end
      COMP_LOOP_C_230 : begin
        fsm_output = 11'b00110110011;
        state_var_NS = COMP_LOOP_C_231;
      end
      COMP_LOOP_C_231 : begin
        fsm_output = 11'b00110110100;
        state_var_NS = COMP_LOOP_C_232;
      end
      COMP_LOOP_C_232 : begin
        fsm_output = 11'b00110110101;
        state_var_NS = COMP_LOOP_C_233;
      end
      COMP_LOOP_C_233 : begin
        fsm_output = 11'b00110110110;
        state_var_NS = COMP_LOOP_C_234;
      end
      COMP_LOOP_C_234 : begin
        fsm_output = 11'b00110110111;
        state_var_NS = COMP_LOOP_C_235;
      end
      COMP_LOOP_C_235 : begin
        fsm_output = 11'b00110111000;
        state_var_NS = COMP_LOOP_C_236;
      end
      COMP_LOOP_C_236 : begin
        fsm_output = 11'b00110111001;
        state_var_NS = COMP_LOOP_C_237;
      end
      COMP_LOOP_C_237 : begin
        fsm_output = 11'b00110111010;
        state_var_NS = COMP_LOOP_C_238;
      end
      COMP_LOOP_C_238 : begin
        fsm_output = 11'b00110111011;
        state_var_NS = COMP_LOOP_C_239;
      end
      COMP_LOOP_C_239 : begin
        fsm_output = 11'b00110111100;
        state_var_NS = COMP_LOOP_C_240;
      end
      COMP_LOOP_C_240 : begin
        fsm_output = 11'b00110111101;
        state_var_NS = COMP_LOOP_C_241;
      end
      COMP_LOOP_C_241 : begin
        fsm_output = 11'b00110111110;
        state_var_NS = COMP_LOOP_C_242;
      end
      COMP_LOOP_C_242 : begin
        fsm_output = 11'b00110111111;
        state_var_NS = COMP_LOOP_C_243;
      end
      COMP_LOOP_C_243 : begin
        fsm_output = 11'b00111000000;
        state_var_NS = COMP_LOOP_C_244;
      end
      COMP_LOOP_C_244 : begin
        fsm_output = 11'b00111000001;
        state_var_NS = COMP_LOOP_C_245;
      end
      COMP_LOOP_C_245 : begin
        fsm_output = 11'b00111000010;
        state_var_NS = COMP_LOOP_C_246;
      end
      COMP_LOOP_C_246 : begin
        fsm_output = 11'b00111000011;
        state_var_NS = COMP_LOOP_C_247;
      end
      COMP_LOOP_C_247 : begin
        fsm_output = 11'b00111000100;
        state_var_NS = COMP_LOOP_C_248;
      end
      COMP_LOOP_C_248 : begin
        fsm_output = 11'b00111000101;
        if ( COMP_LOOP_C_248_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_249;
        end
      end
      COMP_LOOP_C_249 : begin
        fsm_output = 11'b00111000110;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_0;
      end
      COMP_LOOP_5_modExp_1_while_C_0 : begin
        fsm_output = 11'b00111000111;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_1;
      end
      COMP_LOOP_5_modExp_1_while_C_1 : begin
        fsm_output = 11'b00111001000;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_2;
      end
      COMP_LOOP_5_modExp_1_while_C_2 : begin
        fsm_output = 11'b00111001001;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_3;
      end
      COMP_LOOP_5_modExp_1_while_C_3 : begin
        fsm_output = 11'b00111001010;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_4;
      end
      COMP_LOOP_5_modExp_1_while_C_4 : begin
        fsm_output = 11'b00111001011;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_5;
      end
      COMP_LOOP_5_modExp_1_while_C_5 : begin
        fsm_output = 11'b00111001100;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_6;
      end
      COMP_LOOP_5_modExp_1_while_C_6 : begin
        fsm_output = 11'b00111001101;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_7;
      end
      COMP_LOOP_5_modExp_1_while_C_7 : begin
        fsm_output = 11'b00111001110;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_8;
      end
      COMP_LOOP_5_modExp_1_while_C_8 : begin
        fsm_output = 11'b00111001111;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_9;
      end
      COMP_LOOP_5_modExp_1_while_C_9 : begin
        fsm_output = 11'b00111010000;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_10;
      end
      COMP_LOOP_5_modExp_1_while_C_10 : begin
        fsm_output = 11'b00111010001;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_11;
      end
      COMP_LOOP_5_modExp_1_while_C_11 : begin
        fsm_output = 11'b00111010010;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_12;
      end
      COMP_LOOP_5_modExp_1_while_C_12 : begin
        fsm_output = 11'b00111010011;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_13;
      end
      COMP_LOOP_5_modExp_1_while_C_13 : begin
        fsm_output = 11'b00111010100;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_14;
      end
      COMP_LOOP_5_modExp_1_while_C_14 : begin
        fsm_output = 11'b00111010101;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_15;
      end
      COMP_LOOP_5_modExp_1_while_C_15 : begin
        fsm_output = 11'b00111010110;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_16;
      end
      COMP_LOOP_5_modExp_1_while_C_16 : begin
        fsm_output = 11'b00111010111;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_17;
      end
      COMP_LOOP_5_modExp_1_while_C_17 : begin
        fsm_output = 11'b00111011000;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_18;
      end
      COMP_LOOP_5_modExp_1_while_C_18 : begin
        fsm_output = 11'b00111011001;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_19;
      end
      COMP_LOOP_5_modExp_1_while_C_19 : begin
        fsm_output = 11'b00111011010;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_20;
      end
      COMP_LOOP_5_modExp_1_while_C_20 : begin
        fsm_output = 11'b00111011011;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_21;
      end
      COMP_LOOP_5_modExp_1_while_C_21 : begin
        fsm_output = 11'b00111011100;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_22;
      end
      COMP_LOOP_5_modExp_1_while_C_22 : begin
        fsm_output = 11'b00111011101;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_23;
      end
      COMP_LOOP_5_modExp_1_while_C_23 : begin
        fsm_output = 11'b00111011110;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_24;
      end
      COMP_LOOP_5_modExp_1_while_C_24 : begin
        fsm_output = 11'b00111011111;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_25;
      end
      COMP_LOOP_5_modExp_1_while_C_25 : begin
        fsm_output = 11'b00111100000;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_26;
      end
      COMP_LOOP_5_modExp_1_while_C_26 : begin
        fsm_output = 11'b00111100001;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_27;
      end
      COMP_LOOP_5_modExp_1_while_C_27 : begin
        fsm_output = 11'b00111100010;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_28;
      end
      COMP_LOOP_5_modExp_1_while_C_28 : begin
        fsm_output = 11'b00111100011;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_29;
      end
      COMP_LOOP_5_modExp_1_while_C_29 : begin
        fsm_output = 11'b00111100100;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_30;
      end
      COMP_LOOP_5_modExp_1_while_C_30 : begin
        fsm_output = 11'b00111100101;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_31;
      end
      COMP_LOOP_5_modExp_1_while_C_31 : begin
        fsm_output = 11'b00111100110;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_32;
      end
      COMP_LOOP_5_modExp_1_while_C_32 : begin
        fsm_output = 11'b00111100111;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_33;
      end
      COMP_LOOP_5_modExp_1_while_C_33 : begin
        fsm_output = 11'b00111101000;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_34;
      end
      COMP_LOOP_5_modExp_1_while_C_34 : begin
        fsm_output = 11'b00111101001;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_35;
      end
      COMP_LOOP_5_modExp_1_while_C_35 : begin
        fsm_output = 11'b00111101010;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_36;
      end
      COMP_LOOP_5_modExp_1_while_C_36 : begin
        fsm_output = 11'b00111101011;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_37;
      end
      COMP_LOOP_5_modExp_1_while_C_37 : begin
        fsm_output = 11'b00111101100;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_38;
      end
      COMP_LOOP_5_modExp_1_while_C_38 : begin
        fsm_output = 11'b00111101101;
        if ( COMP_LOOP_5_modExp_1_while_C_38_tr0 ) begin
          state_var_NS = COMP_LOOP_C_250;
        end
        else begin
          state_var_NS = COMP_LOOP_5_modExp_1_while_C_0;
        end
      end
      COMP_LOOP_C_250 : begin
        fsm_output = 11'b00111101110;
        state_var_NS = COMP_LOOP_C_251;
      end
      COMP_LOOP_C_251 : begin
        fsm_output = 11'b00111101111;
        state_var_NS = COMP_LOOP_C_252;
      end
      COMP_LOOP_C_252 : begin
        fsm_output = 11'b00111110000;
        state_var_NS = COMP_LOOP_C_253;
      end
      COMP_LOOP_C_253 : begin
        fsm_output = 11'b00111110001;
        state_var_NS = COMP_LOOP_C_254;
      end
      COMP_LOOP_C_254 : begin
        fsm_output = 11'b00111110010;
        state_var_NS = COMP_LOOP_C_255;
      end
      COMP_LOOP_C_255 : begin
        fsm_output = 11'b00111110011;
        state_var_NS = COMP_LOOP_C_256;
      end
      COMP_LOOP_C_256 : begin
        fsm_output = 11'b00111110100;
        state_var_NS = COMP_LOOP_C_257;
      end
      COMP_LOOP_C_257 : begin
        fsm_output = 11'b00111110101;
        state_var_NS = COMP_LOOP_C_258;
      end
      COMP_LOOP_C_258 : begin
        fsm_output = 11'b00111110110;
        state_var_NS = COMP_LOOP_C_259;
      end
      COMP_LOOP_C_259 : begin
        fsm_output = 11'b00111110111;
        state_var_NS = COMP_LOOP_C_260;
      end
      COMP_LOOP_C_260 : begin
        fsm_output = 11'b00111111000;
        state_var_NS = COMP_LOOP_C_261;
      end
      COMP_LOOP_C_261 : begin
        fsm_output = 11'b00111111001;
        state_var_NS = COMP_LOOP_C_262;
      end
      COMP_LOOP_C_262 : begin
        fsm_output = 11'b00111111010;
        state_var_NS = COMP_LOOP_C_263;
      end
      COMP_LOOP_C_263 : begin
        fsm_output = 11'b00111111011;
        state_var_NS = COMP_LOOP_C_264;
      end
      COMP_LOOP_C_264 : begin
        fsm_output = 11'b00111111100;
        state_var_NS = COMP_LOOP_C_265;
      end
      COMP_LOOP_C_265 : begin
        fsm_output = 11'b00111111101;
        state_var_NS = COMP_LOOP_C_266;
      end
      COMP_LOOP_C_266 : begin
        fsm_output = 11'b00111111110;
        state_var_NS = COMP_LOOP_C_267;
      end
      COMP_LOOP_C_267 : begin
        fsm_output = 11'b00111111111;
        state_var_NS = COMP_LOOP_C_268;
      end
      COMP_LOOP_C_268 : begin
        fsm_output = 11'b01000000000;
        state_var_NS = COMP_LOOP_C_269;
      end
      COMP_LOOP_C_269 : begin
        fsm_output = 11'b01000000001;
        state_var_NS = COMP_LOOP_C_270;
      end
      COMP_LOOP_C_270 : begin
        fsm_output = 11'b01000000010;
        state_var_NS = COMP_LOOP_C_271;
      end
      COMP_LOOP_C_271 : begin
        fsm_output = 11'b01000000011;
        state_var_NS = COMP_LOOP_C_272;
      end
      COMP_LOOP_C_272 : begin
        fsm_output = 11'b01000000100;
        state_var_NS = COMP_LOOP_C_273;
      end
      COMP_LOOP_C_273 : begin
        fsm_output = 11'b01000000101;
        state_var_NS = COMP_LOOP_C_274;
      end
      COMP_LOOP_C_274 : begin
        fsm_output = 11'b01000000110;
        state_var_NS = COMP_LOOP_C_275;
      end
      COMP_LOOP_C_275 : begin
        fsm_output = 11'b01000000111;
        state_var_NS = COMP_LOOP_C_276;
      end
      COMP_LOOP_C_276 : begin
        fsm_output = 11'b01000001000;
        state_var_NS = COMP_LOOP_C_277;
      end
      COMP_LOOP_C_277 : begin
        fsm_output = 11'b01000001001;
        state_var_NS = COMP_LOOP_C_278;
      end
      COMP_LOOP_C_278 : begin
        fsm_output = 11'b01000001010;
        state_var_NS = COMP_LOOP_C_279;
      end
      COMP_LOOP_C_279 : begin
        fsm_output = 11'b01000001011;
        state_var_NS = COMP_LOOP_C_280;
      end
      COMP_LOOP_C_280 : begin
        fsm_output = 11'b01000001100;
        state_var_NS = COMP_LOOP_C_281;
      end
      COMP_LOOP_C_281 : begin
        fsm_output = 11'b01000001101;
        state_var_NS = COMP_LOOP_C_282;
      end
      COMP_LOOP_C_282 : begin
        fsm_output = 11'b01000001110;
        state_var_NS = COMP_LOOP_C_283;
      end
      COMP_LOOP_C_283 : begin
        fsm_output = 11'b01000001111;
        state_var_NS = COMP_LOOP_C_284;
      end
      COMP_LOOP_C_284 : begin
        fsm_output = 11'b01000010000;
        state_var_NS = COMP_LOOP_C_285;
      end
      COMP_LOOP_C_285 : begin
        fsm_output = 11'b01000010001;
        state_var_NS = COMP_LOOP_C_286;
      end
      COMP_LOOP_C_286 : begin
        fsm_output = 11'b01000010010;
        state_var_NS = COMP_LOOP_C_287;
      end
      COMP_LOOP_C_287 : begin
        fsm_output = 11'b01000010011;
        state_var_NS = COMP_LOOP_C_288;
      end
      COMP_LOOP_C_288 : begin
        fsm_output = 11'b01000010100;
        state_var_NS = COMP_LOOP_C_289;
      end
      COMP_LOOP_C_289 : begin
        fsm_output = 11'b01000010101;
        state_var_NS = COMP_LOOP_C_290;
      end
      COMP_LOOP_C_290 : begin
        fsm_output = 11'b01000010110;
        state_var_NS = COMP_LOOP_C_291;
      end
      COMP_LOOP_C_291 : begin
        fsm_output = 11'b01000010111;
        state_var_NS = COMP_LOOP_C_292;
      end
      COMP_LOOP_C_292 : begin
        fsm_output = 11'b01000011000;
        state_var_NS = COMP_LOOP_C_293;
      end
      COMP_LOOP_C_293 : begin
        fsm_output = 11'b01000011001;
        state_var_NS = COMP_LOOP_C_294;
      end
      COMP_LOOP_C_294 : begin
        fsm_output = 11'b01000011010;
        state_var_NS = COMP_LOOP_C_295;
      end
      COMP_LOOP_C_295 : begin
        fsm_output = 11'b01000011011;
        state_var_NS = COMP_LOOP_C_296;
      end
      COMP_LOOP_C_296 : begin
        fsm_output = 11'b01000011100;
        state_var_NS = COMP_LOOP_C_297;
      end
      COMP_LOOP_C_297 : begin
        fsm_output = 11'b01000011101;
        state_var_NS = COMP_LOOP_C_298;
      end
      COMP_LOOP_C_298 : begin
        fsm_output = 11'b01000011110;
        state_var_NS = COMP_LOOP_C_299;
      end
      COMP_LOOP_C_299 : begin
        fsm_output = 11'b01000011111;
        state_var_NS = COMP_LOOP_C_300;
      end
      COMP_LOOP_C_300 : begin
        fsm_output = 11'b01000100000;
        state_var_NS = COMP_LOOP_C_301;
      end
      COMP_LOOP_C_301 : begin
        fsm_output = 11'b01000100001;
        state_var_NS = COMP_LOOP_C_302;
      end
      COMP_LOOP_C_302 : begin
        fsm_output = 11'b01000100010;
        state_var_NS = COMP_LOOP_C_303;
      end
      COMP_LOOP_C_303 : begin
        fsm_output = 11'b01000100011;
        state_var_NS = COMP_LOOP_C_304;
      end
      COMP_LOOP_C_304 : begin
        fsm_output = 11'b01000100100;
        state_var_NS = COMP_LOOP_C_305;
      end
      COMP_LOOP_C_305 : begin
        fsm_output = 11'b01000100101;
        state_var_NS = COMP_LOOP_C_306;
      end
      COMP_LOOP_C_306 : begin
        fsm_output = 11'b01000100110;
        state_var_NS = COMP_LOOP_C_307;
      end
      COMP_LOOP_C_307 : begin
        fsm_output = 11'b01000100111;
        state_var_NS = COMP_LOOP_C_308;
      end
      COMP_LOOP_C_308 : begin
        fsm_output = 11'b01000101000;
        state_var_NS = COMP_LOOP_C_309;
      end
      COMP_LOOP_C_309 : begin
        fsm_output = 11'b01000101001;
        state_var_NS = COMP_LOOP_C_310;
      end
      COMP_LOOP_C_310 : begin
        fsm_output = 11'b01000101010;
        if ( COMP_LOOP_C_310_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_311;
        end
      end
      COMP_LOOP_C_311 : begin
        fsm_output = 11'b01000101011;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_0;
      end
      COMP_LOOP_6_modExp_1_while_C_0 : begin
        fsm_output = 11'b01000101100;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_1;
      end
      COMP_LOOP_6_modExp_1_while_C_1 : begin
        fsm_output = 11'b01000101101;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_2;
      end
      COMP_LOOP_6_modExp_1_while_C_2 : begin
        fsm_output = 11'b01000101110;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_3;
      end
      COMP_LOOP_6_modExp_1_while_C_3 : begin
        fsm_output = 11'b01000101111;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_4;
      end
      COMP_LOOP_6_modExp_1_while_C_4 : begin
        fsm_output = 11'b01000110000;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_5;
      end
      COMP_LOOP_6_modExp_1_while_C_5 : begin
        fsm_output = 11'b01000110001;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_6;
      end
      COMP_LOOP_6_modExp_1_while_C_6 : begin
        fsm_output = 11'b01000110010;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_7;
      end
      COMP_LOOP_6_modExp_1_while_C_7 : begin
        fsm_output = 11'b01000110011;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_8;
      end
      COMP_LOOP_6_modExp_1_while_C_8 : begin
        fsm_output = 11'b01000110100;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_9;
      end
      COMP_LOOP_6_modExp_1_while_C_9 : begin
        fsm_output = 11'b01000110101;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_10;
      end
      COMP_LOOP_6_modExp_1_while_C_10 : begin
        fsm_output = 11'b01000110110;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_11;
      end
      COMP_LOOP_6_modExp_1_while_C_11 : begin
        fsm_output = 11'b01000110111;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_12;
      end
      COMP_LOOP_6_modExp_1_while_C_12 : begin
        fsm_output = 11'b01000111000;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_13;
      end
      COMP_LOOP_6_modExp_1_while_C_13 : begin
        fsm_output = 11'b01000111001;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_14;
      end
      COMP_LOOP_6_modExp_1_while_C_14 : begin
        fsm_output = 11'b01000111010;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_15;
      end
      COMP_LOOP_6_modExp_1_while_C_15 : begin
        fsm_output = 11'b01000111011;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_16;
      end
      COMP_LOOP_6_modExp_1_while_C_16 : begin
        fsm_output = 11'b01000111100;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_17;
      end
      COMP_LOOP_6_modExp_1_while_C_17 : begin
        fsm_output = 11'b01000111101;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_18;
      end
      COMP_LOOP_6_modExp_1_while_C_18 : begin
        fsm_output = 11'b01000111110;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_19;
      end
      COMP_LOOP_6_modExp_1_while_C_19 : begin
        fsm_output = 11'b01000111111;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_20;
      end
      COMP_LOOP_6_modExp_1_while_C_20 : begin
        fsm_output = 11'b01001000000;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_21;
      end
      COMP_LOOP_6_modExp_1_while_C_21 : begin
        fsm_output = 11'b01001000001;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_22;
      end
      COMP_LOOP_6_modExp_1_while_C_22 : begin
        fsm_output = 11'b01001000010;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_23;
      end
      COMP_LOOP_6_modExp_1_while_C_23 : begin
        fsm_output = 11'b01001000011;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_24;
      end
      COMP_LOOP_6_modExp_1_while_C_24 : begin
        fsm_output = 11'b01001000100;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_25;
      end
      COMP_LOOP_6_modExp_1_while_C_25 : begin
        fsm_output = 11'b01001000101;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_26;
      end
      COMP_LOOP_6_modExp_1_while_C_26 : begin
        fsm_output = 11'b01001000110;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_27;
      end
      COMP_LOOP_6_modExp_1_while_C_27 : begin
        fsm_output = 11'b01001000111;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_28;
      end
      COMP_LOOP_6_modExp_1_while_C_28 : begin
        fsm_output = 11'b01001001000;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_29;
      end
      COMP_LOOP_6_modExp_1_while_C_29 : begin
        fsm_output = 11'b01001001001;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_30;
      end
      COMP_LOOP_6_modExp_1_while_C_30 : begin
        fsm_output = 11'b01001001010;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_31;
      end
      COMP_LOOP_6_modExp_1_while_C_31 : begin
        fsm_output = 11'b01001001011;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_32;
      end
      COMP_LOOP_6_modExp_1_while_C_32 : begin
        fsm_output = 11'b01001001100;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_33;
      end
      COMP_LOOP_6_modExp_1_while_C_33 : begin
        fsm_output = 11'b01001001101;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_34;
      end
      COMP_LOOP_6_modExp_1_while_C_34 : begin
        fsm_output = 11'b01001001110;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_35;
      end
      COMP_LOOP_6_modExp_1_while_C_35 : begin
        fsm_output = 11'b01001001111;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_36;
      end
      COMP_LOOP_6_modExp_1_while_C_36 : begin
        fsm_output = 11'b01001010000;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_37;
      end
      COMP_LOOP_6_modExp_1_while_C_37 : begin
        fsm_output = 11'b01001010001;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_38;
      end
      COMP_LOOP_6_modExp_1_while_C_38 : begin
        fsm_output = 11'b01001010010;
        if ( COMP_LOOP_6_modExp_1_while_C_38_tr0 ) begin
          state_var_NS = COMP_LOOP_C_312;
        end
        else begin
          state_var_NS = COMP_LOOP_6_modExp_1_while_C_0;
        end
      end
      COMP_LOOP_C_312 : begin
        fsm_output = 11'b01001010011;
        state_var_NS = COMP_LOOP_C_313;
      end
      COMP_LOOP_C_313 : begin
        fsm_output = 11'b01001010100;
        state_var_NS = COMP_LOOP_C_314;
      end
      COMP_LOOP_C_314 : begin
        fsm_output = 11'b01001010101;
        state_var_NS = COMP_LOOP_C_315;
      end
      COMP_LOOP_C_315 : begin
        fsm_output = 11'b01001010110;
        state_var_NS = COMP_LOOP_C_316;
      end
      COMP_LOOP_C_316 : begin
        fsm_output = 11'b01001010111;
        state_var_NS = COMP_LOOP_C_317;
      end
      COMP_LOOP_C_317 : begin
        fsm_output = 11'b01001011000;
        state_var_NS = COMP_LOOP_C_318;
      end
      COMP_LOOP_C_318 : begin
        fsm_output = 11'b01001011001;
        state_var_NS = COMP_LOOP_C_319;
      end
      COMP_LOOP_C_319 : begin
        fsm_output = 11'b01001011010;
        state_var_NS = COMP_LOOP_C_320;
      end
      COMP_LOOP_C_320 : begin
        fsm_output = 11'b01001011011;
        state_var_NS = COMP_LOOP_C_321;
      end
      COMP_LOOP_C_321 : begin
        fsm_output = 11'b01001011100;
        state_var_NS = COMP_LOOP_C_322;
      end
      COMP_LOOP_C_322 : begin
        fsm_output = 11'b01001011101;
        state_var_NS = COMP_LOOP_C_323;
      end
      COMP_LOOP_C_323 : begin
        fsm_output = 11'b01001011110;
        state_var_NS = COMP_LOOP_C_324;
      end
      COMP_LOOP_C_324 : begin
        fsm_output = 11'b01001011111;
        state_var_NS = COMP_LOOP_C_325;
      end
      COMP_LOOP_C_325 : begin
        fsm_output = 11'b01001100000;
        state_var_NS = COMP_LOOP_C_326;
      end
      COMP_LOOP_C_326 : begin
        fsm_output = 11'b01001100001;
        state_var_NS = COMP_LOOP_C_327;
      end
      COMP_LOOP_C_327 : begin
        fsm_output = 11'b01001100010;
        state_var_NS = COMP_LOOP_C_328;
      end
      COMP_LOOP_C_328 : begin
        fsm_output = 11'b01001100011;
        state_var_NS = COMP_LOOP_C_329;
      end
      COMP_LOOP_C_329 : begin
        fsm_output = 11'b01001100100;
        state_var_NS = COMP_LOOP_C_330;
      end
      COMP_LOOP_C_330 : begin
        fsm_output = 11'b01001100101;
        state_var_NS = COMP_LOOP_C_331;
      end
      COMP_LOOP_C_331 : begin
        fsm_output = 11'b01001100110;
        state_var_NS = COMP_LOOP_C_332;
      end
      COMP_LOOP_C_332 : begin
        fsm_output = 11'b01001100111;
        state_var_NS = COMP_LOOP_C_333;
      end
      COMP_LOOP_C_333 : begin
        fsm_output = 11'b01001101000;
        state_var_NS = COMP_LOOP_C_334;
      end
      COMP_LOOP_C_334 : begin
        fsm_output = 11'b01001101001;
        state_var_NS = COMP_LOOP_C_335;
      end
      COMP_LOOP_C_335 : begin
        fsm_output = 11'b01001101010;
        state_var_NS = COMP_LOOP_C_336;
      end
      COMP_LOOP_C_336 : begin
        fsm_output = 11'b01001101011;
        state_var_NS = COMP_LOOP_C_337;
      end
      COMP_LOOP_C_337 : begin
        fsm_output = 11'b01001101100;
        state_var_NS = COMP_LOOP_C_338;
      end
      COMP_LOOP_C_338 : begin
        fsm_output = 11'b01001101101;
        state_var_NS = COMP_LOOP_C_339;
      end
      COMP_LOOP_C_339 : begin
        fsm_output = 11'b01001101110;
        state_var_NS = COMP_LOOP_C_340;
      end
      COMP_LOOP_C_340 : begin
        fsm_output = 11'b01001101111;
        state_var_NS = COMP_LOOP_C_341;
      end
      COMP_LOOP_C_341 : begin
        fsm_output = 11'b01001110000;
        state_var_NS = COMP_LOOP_C_342;
      end
      COMP_LOOP_C_342 : begin
        fsm_output = 11'b01001110001;
        state_var_NS = COMP_LOOP_C_343;
      end
      COMP_LOOP_C_343 : begin
        fsm_output = 11'b01001110010;
        state_var_NS = COMP_LOOP_C_344;
      end
      COMP_LOOP_C_344 : begin
        fsm_output = 11'b01001110011;
        state_var_NS = COMP_LOOP_C_345;
      end
      COMP_LOOP_C_345 : begin
        fsm_output = 11'b01001110100;
        state_var_NS = COMP_LOOP_C_346;
      end
      COMP_LOOP_C_346 : begin
        fsm_output = 11'b01001110101;
        state_var_NS = COMP_LOOP_C_347;
      end
      COMP_LOOP_C_347 : begin
        fsm_output = 11'b01001110110;
        state_var_NS = COMP_LOOP_C_348;
      end
      COMP_LOOP_C_348 : begin
        fsm_output = 11'b01001110111;
        state_var_NS = COMP_LOOP_C_349;
      end
      COMP_LOOP_C_349 : begin
        fsm_output = 11'b01001111000;
        state_var_NS = COMP_LOOP_C_350;
      end
      COMP_LOOP_C_350 : begin
        fsm_output = 11'b01001111001;
        state_var_NS = COMP_LOOP_C_351;
      end
      COMP_LOOP_C_351 : begin
        fsm_output = 11'b01001111010;
        state_var_NS = COMP_LOOP_C_352;
      end
      COMP_LOOP_C_352 : begin
        fsm_output = 11'b01001111011;
        state_var_NS = COMP_LOOP_C_353;
      end
      COMP_LOOP_C_353 : begin
        fsm_output = 11'b01001111100;
        state_var_NS = COMP_LOOP_C_354;
      end
      COMP_LOOP_C_354 : begin
        fsm_output = 11'b01001111101;
        state_var_NS = COMP_LOOP_C_355;
      end
      COMP_LOOP_C_355 : begin
        fsm_output = 11'b01001111110;
        state_var_NS = COMP_LOOP_C_356;
      end
      COMP_LOOP_C_356 : begin
        fsm_output = 11'b01001111111;
        state_var_NS = COMP_LOOP_C_357;
      end
      COMP_LOOP_C_357 : begin
        fsm_output = 11'b01010000000;
        state_var_NS = COMP_LOOP_C_358;
      end
      COMP_LOOP_C_358 : begin
        fsm_output = 11'b01010000001;
        state_var_NS = COMP_LOOP_C_359;
      end
      COMP_LOOP_C_359 : begin
        fsm_output = 11'b01010000010;
        state_var_NS = COMP_LOOP_C_360;
      end
      COMP_LOOP_C_360 : begin
        fsm_output = 11'b01010000011;
        state_var_NS = COMP_LOOP_C_361;
      end
      COMP_LOOP_C_361 : begin
        fsm_output = 11'b01010000100;
        state_var_NS = COMP_LOOP_C_362;
      end
      COMP_LOOP_C_362 : begin
        fsm_output = 11'b01010000101;
        state_var_NS = COMP_LOOP_C_363;
      end
      COMP_LOOP_C_363 : begin
        fsm_output = 11'b01010000110;
        state_var_NS = COMP_LOOP_C_364;
      end
      COMP_LOOP_C_364 : begin
        fsm_output = 11'b01010000111;
        state_var_NS = COMP_LOOP_C_365;
      end
      COMP_LOOP_C_365 : begin
        fsm_output = 11'b01010001000;
        state_var_NS = COMP_LOOP_C_366;
      end
      COMP_LOOP_C_366 : begin
        fsm_output = 11'b01010001001;
        state_var_NS = COMP_LOOP_C_367;
      end
      COMP_LOOP_C_367 : begin
        fsm_output = 11'b01010001010;
        state_var_NS = COMP_LOOP_C_368;
      end
      COMP_LOOP_C_368 : begin
        fsm_output = 11'b01010001011;
        state_var_NS = COMP_LOOP_C_369;
      end
      COMP_LOOP_C_369 : begin
        fsm_output = 11'b01010001100;
        state_var_NS = COMP_LOOP_C_370;
      end
      COMP_LOOP_C_370 : begin
        fsm_output = 11'b01010001101;
        state_var_NS = COMP_LOOP_C_371;
      end
      COMP_LOOP_C_371 : begin
        fsm_output = 11'b01010001110;
        state_var_NS = COMP_LOOP_C_372;
      end
      COMP_LOOP_C_372 : begin
        fsm_output = 11'b01010001111;
        if ( COMP_LOOP_C_372_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_373;
        end
      end
      COMP_LOOP_C_373 : begin
        fsm_output = 11'b01010010000;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_0;
      end
      COMP_LOOP_7_modExp_1_while_C_0 : begin
        fsm_output = 11'b01010010001;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_1;
      end
      COMP_LOOP_7_modExp_1_while_C_1 : begin
        fsm_output = 11'b01010010010;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_2;
      end
      COMP_LOOP_7_modExp_1_while_C_2 : begin
        fsm_output = 11'b01010010011;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_3;
      end
      COMP_LOOP_7_modExp_1_while_C_3 : begin
        fsm_output = 11'b01010010100;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_4;
      end
      COMP_LOOP_7_modExp_1_while_C_4 : begin
        fsm_output = 11'b01010010101;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_5;
      end
      COMP_LOOP_7_modExp_1_while_C_5 : begin
        fsm_output = 11'b01010010110;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_6;
      end
      COMP_LOOP_7_modExp_1_while_C_6 : begin
        fsm_output = 11'b01010010111;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_7;
      end
      COMP_LOOP_7_modExp_1_while_C_7 : begin
        fsm_output = 11'b01010011000;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_8;
      end
      COMP_LOOP_7_modExp_1_while_C_8 : begin
        fsm_output = 11'b01010011001;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_9;
      end
      COMP_LOOP_7_modExp_1_while_C_9 : begin
        fsm_output = 11'b01010011010;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_10;
      end
      COMP_LOOP_7_modExp_1_while_C_10 : begin
        fsm_output = 11'b01010011011;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_11;
      end
      COMP_LOOP_7_modExp_1_while_C_11 : begin
        fsm_output = 11'b01010011100;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_12;
      end
      COMP_LOOP_7_modExp_1_while_C_12 : begin
        fsm_output = 11'b01010011101;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_13;
      end
      COMP_LOOP_7_modExp_1_while_C_13 : begin
        fsm_output = 11'b01010011110;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_14;
      end
      COMP_LOOP_7_modExp_1_while_C_14 : begin
        fsm_output = 11'b01010011111;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_15;
      end
      COMP_LOOP_7_modExp_1_while_C_15 : begin
        fsm_output = 11'b01010100000;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_16;
      end
      COMP_LOOP_7_modExp_1_while_C_16 : begin
        fsm_output = 11'b01010100001;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_17;
      end
      COMP_LOOP_7_modExp_1_while_C_17 : begin
        fsm_output = 11'b01010100010;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_18;
      end
      COMP_LOOP_7_modExp_1_while_C_18 : begin
        fsm_output = 11'b01010100011;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_19;
      end
      COMP_LOOP_7_modExp_1_while_C_19 : begin
        fsm_output = 11'b01010100100;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_20;
      end
      COMP_LOOP_7_modExp_1_while_C_20 : begin
        fsm_output = 11'b01010100101;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_21;
      end
      COMP_LOOP_7_modExp_1_while_C_21 : begin
        fsm_output = 11'b01010100110;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_22;
      end
      COMP_LOOP_7_modExp_1_while_C_22 : begin
        fsm_output = 11'b01010100111;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_23;
      end
      COMP_LOOP_7_modExp_1_while_C_23 : begin
        fsm_output = 11'b01010101000;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_24;
      end
      COMP_LOOP_7_modExp_1_while_C_24 : begin
        fsm_output = 11'b01010101001;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_25;
      end
      COMP_LOOP_7_modExp_1_while_C_25 : begin
        fsm_output = 11'b01010101010;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_26;
      end
      COMP_LOOP_7_modExp_1_while_C_26 : begin
        fsm_output = 11'b01010101011;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_27;
      end
      COMP_LOOP_7_modExp_1_while_C_27 : begin
        fsm_output = 11'b01010101100;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_28;
      end
      COMP_LOOP_7_modExp_1_while_C_28 : begin
        fsm_output = 11'b01010101101;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_29;
      end
      COMP_LOOP_7_modExp_1_while_C_29 : begin
        fsm_output = 11'b01010101110;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_30;
      end
      COMP_LOOP_7_modExp_1_while_C_30 : begin
        fsm_output = 11'b01010101111;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_31;
      end
      COMP_LOOP_7_modExp_1_while_C_31 : begin
        fsm_output = 11'b01010110000;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_32;
      end
      COMP_LOOP_7_modExp_1_while_C_32 : begin
        fsm_output = 11'b01010110001;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_33;
      end
      COMP_LOOP_7_modExp_1_while_C_33 : begin
        fsm_output = 11'b01010110010;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_34;
      end
      COMP_LOOP_7_modExp_1_while_C_34 : begin
        fsm_output = 11'b01010110011;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_35;
      end
      COMP_LOOP_7_modExp_1_while_C_35 : begin
        fsm_output = 11'b01010110100;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_36;
      end
      COMP_LOOP_7_modExp_1_while_C_36 : begin
        fsm_output = 11'b01010110101;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_37;
      end
      COMP_LOOP_7_modExp_1_while_C_37 : begin
        fsm_output = 11'b01010110110;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_38;
      end
      COMP_LOOP_7_modExp_1_while_C_38 : begin
        fsm_output = 11'b01010110111;
        if ( COMP_LOOP_7_modExp_1_while_C_38_tr0 ) begin
          state_var_NS = COMP_LOOP_C_374;
        end
        else begin
          state_var_NS = COMP_LOOP_7_modExp_1_while_C_0;
        end
      end
      COMP_LOOP_C_374 : begin
        fsm_output = 11'b01010111000;
        state_var_NS = COMP_LOOP_C_375;
      end
      COMP_LOOP_C_375 : begin
        fsm_output = 11'b01010111001;
        state_var_NS = COMP_LOOP_C_376;
      end
      COMP_LOOP_C_376 : begin
        fsm_output = 11'b01010111010;
        state_var_NS = COMP_LOOP_C_377;
      end
      COMP_LOOP_C_377 : begin
        fsm_output = 11'b01010111011;
        state_var_NS = COMP_LOOP_C_378;
      end
      COMP_LOOP_C_378 : begin
        fsm_output = 11'b01010111100;
        state_var_NS = COMP_LOOP_C_379;
      end
      COMP_LOOP_C_379 : begin
        fsm_output = 11'b01010111101;
        state_var_NS = COMP_LOOP_C_380;
      end
      COMP_LOOP_C_380 : begin
        fsm_output = 11'b01010111110;
        state_var_NS = COMP_LOOP_C_381;
      end
      COMP_LOOP_C_381 : begin
        fsm_output = 11'b01010111111;
        state_var_NS = COMP_LOOP_C_382;
      end
      COMP_LOOP_C_382 : begin
        fsm_output = 11'b01011000000;
        state_var_NS = COMP_LOOP_C_383;
      end
      COMP_LOOP_C_383 : begin
        fsm_output = 11'b01011000001;
        state_var_NS = COMP_LOOP_C_384;
      end
      COMP_LOOP_C_384 : begin
        fsm_output = 11'b01011000010;
        state_var_NS = COMP_LOOP_C_385;
      end
      COMP_LOOP_C_385 : begin
        fsm_output = 11'b01011000011;
        state_var_NS = COMP_LOOP_C_386;
      end
      COMP_LOOP_C_386 : begin
        fsm_output = 11'b01011000100;
        state_var_NS = COMP_LOOP_C_387;
      end
      COMP_LOOP_C_387 : begin
        fsm_output = 11'b01011000101;
        state_var_NS = COMP_LOOP_C_388;
      end
      COMP_LOOP_C_388 : begin
        fsm_output = 11'b01011000110;
        state_var_NS = COMP_LOOP_C_389;
      end
      COMP_LOOP_C_389 : begin
        fsm_output = 11'b01011000111;
        state_var_NS = COMP_LOOP_C_390;
      end
      COMP_LOOP_C_390 : begin
        fsm_output = 11'b01011001000;
        state_var_NS = COMP_LOOP_C_391;
      end
      COMP_LOOP_C_391 : begin
        fsm_output = 11'b01011001001;
        state_var_NS = COMP_LOOP_C_392;
      end
      COMP_LOOP_C_392 : begin
        fsm_output = 11'b01011001010;
        state_var_NS = COMP_LOOP_C_393;
      end
      COMP_LOOP_C_393 : begin
        fsm_output = 11'b01011001011;
        state_var_NS = COMP_LOOP_C_394;
      end
      COMP_LOOP_C_394 : begin
        fsm_output = 11'b01011001100;
        state_var_NS = COMP_LOOP_C_395;
      end
      COMP_LOOP_C_395 : begin
        fsm_output = 11'b01011001101;
        state_var_NS = COMP_LOOP_C_396;
      end
      COMP_LOOP_C_396 : begin
        fsm_output = 11'b01011001110;
        state_var_NS = COMP_LOOP_C_397;
      end
      COMP_LOOP_C_397 : begin
        fsm_output = 11'b01011001111;
        state_var_NS = COMP_LOOP_C_398;
      end
      COMP_LOOP_C_398 : begin
        fsm_output = 11'b01011010000;
        state_var_NS = COMP_LOOP_C_399;
      end
      COMP_LOOP_C_399 : begin
        fsm_output = 11'b01011010001;
        state_var_NS = COMP_LOOP_C_400;
      end
      COMP_LOOP_C_400 : begin
        fsm_output = 11'b01011010010;
        state_var_NS = COMP_LOOP_C_401;
      end
      COMP_LOOP_C_401 : begin
        fsm_output = 11'b01011010011;
        state_var_NS = COMP_LOOP_C_402;
      end
      COMP_LOOP_C_402 : begin
        fsm_output = 11'b01011010100;
        state_var_NS = COMP_LOOP_C_403;
      end
      COMP_LOOP_C_403 : begin
        fsm_output = 11'b01011010101;
        state_var_NS = COMP_LOOP_C_404;
      end
      COMP_LOOP_C_404 : begin
        fsm_output = 11'b01011010110;
        state_var_NS = COMP_LOOP_C_405;
      end
      COMP_LOOP_C_405 : begin
        fsm_output = 11'b01011010111;
        state_var_NS = COMP_LOOP_C_406;
      end
      COMP_LOOP_C_406 : begin
        fsm_output = 11'b01011011000;
        state_var_NS = COMP_LOOP_C_407;
      end
      COMP_LOOP_C_407 : begin
        fsm_output = 11'b01011011001;
        state_var_NS = COMP_LOOP_C_408;
      end
      COMP_LOOP_C_408 : begin
        fsm_output = 11'b01011011010;
        state_var_NS = COMP_LOOP_C_409;
      end
      COMP_LOOP_C_409 : begin
        fsm_output = 11'b01011011011;
        state_var_NS = COMP_LOOP_C_410;
      end
      COMP_LOOP_C_410 : begin
        fsm_output = 11'b01011011100;
        state_var_NS = COMP_LOOP_C_411;
      end
      COMP_LOOP_C_411 : begin
        fsm_output = 11'b01011011101;
        state_var_NS = COMP_LOOP_C_412;
      end
      COMP_LOOP_C_412 : begin
        fsm_output = 11'b01011011110;
        state_var_NS = COMP_LOOP_C_413;
      end
      COMP_LOOP_C_413 : begin
        fsm_output = 11'b01011011111;
        state_var_NS = COMP_LOOP_C_414;
      end
      COMP_LOOP_C_414 : begin
        fsm_output = 11'b01011100000;
        state_var_NS = COMP_LOOP_C_415;
      end
      COMP_LOOP_C_415 : begin
        fsm_output = 11'b01011100001;
        state_var_NS = COMP_LOOP_C_416;
      end
      COMP_LOOP_C_416 : begin
        fsm_output = 11'b01011100010;
        state_var_NS = COMP_LOOP_C_417;
      end
      COMP_LOOP_C_417 : begin
        fsm_output = 11'b01011100011;
        state_var_NS = COMP_LOOP_C_418;
      end
      COMP_LOOP_C_418 : begin
        fsm_output = 11'b01011100100;
        state_var_NS = COMP_LOOP_C_419;
      end
      COMP_LOOP_C_419 : begin
        fsm_output = 11'b01011100101;
        state_var_NS = COMP_LOOP_C_420;
      end
      COMP_LOOP_C_420 : begin
        fsm_output = 11'b01011100110;
        state_var_NS = COMP_LOOP_C_421;
      end
      COMP_LOOP_C_421 : begin
        fsm_output = 11'b01011100111;
        state_var_NS = COMP_LOOP_C_422;
      end
      COMP_LOOP_C_422 : begin
        fsm_output = 11'b01011101000;
        state_var_NS = COMP_LOOP_C_423;
      end
      COMP_LOOP_C_423 : begin
        fsm_output = 11'b01011101001;
        state_var_NS = COMP_LOOP_C_424;
      end
      COMP_LOOP_C_424 : begin
        fsm_output = 11'b01011101010;
        state_var_NS = COMP_LOOP_C_425;
      end
      COMP_LOOP_C_425 : begin
        fsm_output = 11'b01011101011;
        state_var_NS = COMP_LOOP_C_426;
      end
      COMP_LOOP_C_426 : begin
        fsm_output = 11'b01011101100;
        state_var_NS = COMP_LOOP_C_427;
      end
      COMP_LOOP_C_427 : begin
        fsm_output = 11'b01011101101;
        state_var_NS = COMP_LOOP_C_428;
      end
      COMP_LOOP_C_428 : begin
        fsm_output = 11'b01011101110;
        state_var_NS = COMP_LOOP_C_429;
      end
      COMP_LOOP_C_429 : begin
        fsm_output = 11'b01011101111;
        state_var_NS = COMP_LOOP_C_430;
      end
      COMP_LOOP_C_430 : begin
        fsm_output = 11'b01011110000;
        state_var_NS = COMP_LOOP_C_431;
      end
      COMP_LOOP_C_431 : begin
        fsm_output = 11'b01011110001;
        state_var_NS = COMP_LOOP_C_432;
      end
      COMP_LOOP_C_432 : begin
        fsm_output = 11'b01011110010;
        state_var_NS = COMP_LOOP_C_433;
      end
      COMP_LOOP_C_433 : begin
        fsm_output = 11'b01011110011;
        state_var_NS = COMP_LOOP_C_434;
      end
      COMP_LOOP_C_434 : begin
        fsm_output = 11'b01011110100;
        if ( COMP_LOOP_C_434_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_435;
        end
      end
      COMP_LOOP_C_435 : begin
        fsm_output = 11'b01011110101;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_0;
      end
      COMP_LOOP_8_modExp_1_while_C_0 : begin
        fsm_output = 11'b01011110110;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_1;
      end
      COMP_LOOP_8_modExp_1_while_C_1 : begin
        fsm_output = 11'b01011110111;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_2;
      end
      COMP_LOOP_8_modExp_1_while_C_2 : begin
        fsm_output = 11'b01011111000;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_3;
      end
      COMP_LOOP_8_modExp_1_while_C_3 : begin
        fsm_output = 11'b01011111001;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_4;
      end
      COMP_LOOP_8_modExp_1_while_C_4 : begin
        fsm_output = 11'b01011111010;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_5;
      end
      COMP_LOOP_8_modExp_1_while_C_5 : begin
        fsm_output = 11'b01011111011;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_6;
      end
      COMP_LOOP_8_modExp_1_while_C_6 : begin
        fsm_output = 11'b01011111100;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_7;
      end
      COMP_LOOP_8_modExp_1_while_C_7 : begin
        fsm_output = 11'b01011111101;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_8;
      end
      COMP_LOOP_8_modExp_1_while_C_8 : begin
        fsm_output = 11'b01011111110;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_9;
      end
      COMP_LOOP_8_modExp_1_while_C_9 : begin
        fsm_output = 11'b01011111111;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_10;
      end
      COMP_LOOP_8_modExp_1_while_C_10 : begin
        fsm_output = 11'b01100000000;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_11;
      end
      COMP_LOOP_8_modExp_1_while_C_11 : begin
        fsm_output = 11'b01100000001;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_12;
      end
      COMP_LOOP_8_modExp_1_while_C_12 : begin
        fsm_output = 11'b01100000010;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_13;
      end
      COMP_LOOP_8_modExp_1_while_C_13 : begin
        fsm_output = 11'b01100000011;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_14;
      end
      COMP_LOOP_8_modExp_1_while_C_14 : begin
        fsm_output = 11'b01100000100;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_15;
      end
      COMP_LOOP_8_modExp_1_while_C_15 : begin
        fsm_output = 11'b01100000101;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_16;
      end
      COMP_LOOP_8_modExp_1_while_C_16 : begin
        fsm_output = 11'b01100000110;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_17;
      end
      COMP_LOOP_8_modExp_1_while_C_17 : begin
        fsm_output = 11'b01100000111;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_18;
      end
      COMP_LOOP_8_modExp_1_while_C_18 : begin
        fsm_output = 11'b01100001000;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_19;
      end
      COMP_LOOP_8_modExp_1_while_C_19 : begin
        fsm_output = 11'b01100001001;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_20;
      end
      COMP_LOOP_8_modExp_1_while_C_20 : begin
        fsm_output = 11'b01100001010;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_21;
      end
      COMP_LOOP_8_modExp_1_while_C_21 : begin
        fsm_output = 11'b01100001011;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_22;
      end
      COMP_LOOP_8_modExp_1_while_C_22 : begin
        fsm_output = 11'b01100001100;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_23;
      end
      COMP_LOOP_8_modExp_1_while_C_23 : begin
        fsm_output = 11'b01100001101;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_24;
      end
      COMP_LOOP_8_modExp_1_while_C_24 : begin
        fsm_output = 11'b01100001110;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_25;
      end
      COMP_LOOP_8_modExp_1_while_C_25 : begin
        fsm_output = 11'b01100001111;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_26;
      end
      COMP_LOOP_8_modExp_1_while_C_26 : begin
        fsm_output = 11'b01100010000;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_27;
      end
      COMP_LOOP_8_modExp_1_while_C_27 : begin
        fsm_output = 11'b01100010001;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_28;
      end
      COMP_LOOP_8_modExp_1_while_C_28 : begin
        fsm_output = 11'b01100010010;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_29;
      end
      COMP_LOOP_8_modExp_1_while_C_29 : begin
        fsm_output = 11'b01100010011;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_30;
      end
      COMP_LOOP_8_modExp_1_while_C_30 : begin
        fsm_output = 11'b01100010100;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_31;
      end
      COMP_LOOP_8_modExp_1_while_C_31 : begin
        fsm_output = 11'b01100010101;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_32;
      end
      COMP_LOOP_8_modExp_1_while_C_32 : begin
        fsm_output = 11'b01100010110;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_33;
      end
      COMP_LOOP_8_modExp_1_while_C_33 : begin
        fsm_output = 11'b01100010111;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_34;
      end
      COMP_LOOP_8_modExp_1_while_C_34 : begin
        fsm_output = 11'b01100011000;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_35;
      end
      COMP_LOOP_8_modExp_1_while_C_35 : begin
        fsm_output = 11'b01100011001;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_36;
      end
      COMP_LOOP_8_modExp_1_while_C_36 : begin
        fsm_output = 11'b01100011010;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_37;
      end
      COMP_LOOP_8_modExp_1_while_C_37 : begin
        fsm_output = 11'b01100011011;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_38;
      end
      COMP_LOOP_8_modExp_1_while_C_38 : begin
        fsm_output = 11'b01100011100;
        if ( COMP_LOOP_8_modExp_1_while_C_38_tr0 ) begin
          state_var_NS = COMP_LOOP_C_436;
        end
        else begin
          state_var_NS = COMP_LOOP_8_modExp_1_while_C_0;
        end
      end
      COMP_LOOP_C_436 : begin
        fsm_output = 11'b01100011101;
        state_var_NS = COMP_LOOP_C_437;
      end
      COMP_LOOP_C_437 : begin
        fsm_output = 11'b01100011110;
        state_var_NS = COMP_LOOP_C_438;
      end
      COMP_LOOP_C_438 : begin
        fsm_output = 11'b01100011111;
        state_var_NS = COMP_LOOP_C_439;
      end
      COMP_LOOP_C_439 : begin
        fsm_output = 11'b01100100000;
        state_var_NS = COMP_LOOP_C_440;
      end
      COMP_LOOP_C_440 : begin
        fsm_output = 11'b01100100001;
        state_var_NS = COMP_LOOP_C_441;
      end
      COMP_LOOP_C_441 : begin
        fsm_output = 11'b01100100010;
        state_var_NS = COMP_LOOP_C_442;
      end
      COMP_LOOP_C_442 : begin
        fsm_output = 11'b01100100011;
        state_var_NS = COMP_LOOP_C_443;
      end
      COMP_LOOP_C_443 : begin
        fsm_output = 11'b01100100100;
        state_var_NS = COMP_LOOP_C_444;
      end
      COMP_LOOP_C_444 : begin
        fsm_output = 11'b01100100101;
        state_var_NS = COMP_LOOP_C_445;
      end
      COMP_LOOP_C_445 : begin
        fsm_output = 11'b01100100110;
        state_var_NS = COMP_LOOP_C_446;
      end
      COMP_LOOP_C_446 : begin
        fsm_output = 11'b01100100111;
        state_var_NS = COMP_LOOP_C_447;
      end
      COMP_LOOP_C_447 : begin
        fsm_output = 11'b01100101000;
        state_var_NS = COMP_LOOP_C_448;
      end
      COMP_LOOP_C_448 : begin
        fsm_output = 11'b01100101001;
        state_var_NS = COMP_LOOP_C_449;
      end
      COMP_LOOP_C_449 : begin
        fsm_output = 11'b01100101010;
        state_var_NS = COMP_LOOP_C_450;
      end
      COMP_LOOP_C_450 : begin
        fsm_output = 11'b01100101011;
        state_var_NS = COMP_LOOP_C_451;
      end
      COMP_LOOP_C_451 : begin
        fsm_output = 11'b01100101100;
        state_var_NS = COMP_LOOP_C_452;
      end
      COMP_LOOP_C_452 : begin
        fsm_output = 11'b01100101101;
        state_var_NS = COMP_LOOP_C_453;
      end
      COMP_LOOP_C_453 : begin
        fsm_output = 11'b01100101110;
        state_var_NS = COMP_LOOP_C_454;
      end
      COMP_LOOP_C_454 : begin
        fsm_output = 11'b01100101111;
        state_var_NS = COMP_LOOP_C_455;
      end
      COMP_LOOP_C_455 : begin
        fsm_output = 11'b01100110000;
        state_var_NS = COMP_LOOP_C_456;
      end
      COMP_LOOP_C_456 : begin
        fsm_output = 11'b01100110001;
        state_var_NS = COMP_LOOP_C_457;
      end
      COMP_LOOP_C_457 : begin
        fsm_output = 11'b01100110010;
        state_var_NS = COMP_LOOP_C_458;
      end
      COMP_LOOP_C_458 : begin
        fsm_output = 11'b01100110011;
        state_var_NS = COMP_LOOP_C_459;
      end
      COMP_LOOP_C_459 : begin
        fsm_output = 11'b01100110100;
        state_var_NS = COMP_LOOP_C_460;
      end
      COMP_LOOP_C_460 : begin
        fsm_output = 11'b01100110101;
        state_var_NS = COMP_LOOP_C_461;
      end
      COMP_LOOP_C_461 : begin
        fsm_output = 11'b01100110110;
        state_var_NS = COMP_LOOP_C_462;
      end
      COMP_LOOP_C_462 : begin
        fsm_output = 11'b01100110111;
        state_var_NS = COMP_LOOP_C_463;
      end
      COMP_LOOP_C_463 : begin
        fsm_output = 11'b01100111000;
        state_var_NS = COMP_LOOP_C_464;
      end
      COMP_LOOP_C_464 : begin
        fsm_output = 11'b01100111001;
        state_var_NS = COMP_LOOP_C_465;
      end
      COMP_LOOP_C_465 : begin
        fsm_output = 11'b01100111010;
        state_var_NS = COMP_LOOP_C_466;
      end
      COMP_LOOP_C_466 : begin
        fsm_output = 11'b01100111011;
        state_var_NS = COMP_LOOP_C_467;
      end
      COMP_LOOP_C_467 : begin
        fsm_output = 11'b01100111100;
        state_var_NS = COMP_LOOP_C_468;
      end
      COMP_LOOP_C_468 : begin
        fsm_output = 11'b01100111101;
        state_var_NS = COMP_LOOP_C_469;
      end
      COMP_LOOP_C_469 : begin
        fsm_output = 11'b01100111110;
        state_var_NS = COMP_LOOP_C_470;
      end
      COMP_LOOP_C_470 : begin
        fsm_output = 11'b01100111111;
        state_var_NS = COMP_LOOP_C_471;
      end
      COMP_LOOP_C_471 : begin
        fsm_output = 11'b01101000000;
        state_var_NS = COMP_LOOP_C_472;
      end
      COMP_LOOP_C_472 : begin
        fsm_output = 11'b01101000001;
        state_var_NS = COMP_LOOP_C_473;
      end
      COMP_LOOP_C_473 : begin
        fsm_output = 11'b01101000010;
        state_var_NS = COMP_LOOP_C_474;
      end
      COMP_LOOP_C_474 : begin
        fsm_output = 11'b01101000011;
        state_var_NS = COMP_LOOP_C_475;
      end
      COMP_LOOP_C_475 : begin
        fsm_output = 11'b01101000100;
        state_var_NS = COMP_LOOP_C_476;
      end
      COMP_LOOP_C_476 : begin
        fsm_output = 11'b01101000101;
        state_var_NS = COMP_LOOP_C_477;
      end
      COMP_LOOP_C_477 : begin
        fsm_output = 11'b01101000110;
        state_var_NS = COMP_LOOP_C_478;
      end
      COMP_LOOP_C_478 : begin
        fsm_output = 11'b01101000111;
        state_var_NS = COMP_LOOP_C_479;
      end
      COMP_LOOP_C_479 : begin
        fsm_output = 11'b01101001000;
        state_var_NS = COMP_LOOP_C_480;
      end
      COMP_LOOP_C_480 : begin
        fsm_output = 11'b01101001001;
        state_var_NS = COMP_LOOP_C_481;
      end
      COMP_LOOP_C_481 : begin
        fsm_output = 11'b01101001010;
        state_var_NS = COMP_LOOP_C_482;
      end
      COMP_LOOP_C_482 : begin
        fsm_output = 11'b01101001011;
        state_var_NS = COMP_LOOP_C_483;
      end
      COMP_LOOP_C_483 : begin
        fsm_output = 11'b01101001100;
        state_var_NS = COMP_LOOP_C_484;
      end
      COMP_LOOP_C_484 : begin
        fsm_output = 11'b01101001101;
        state_var_NS = COMP_LOOP_C_485;
      end
      COMP_LOOP_C_485 : begin
        fsm_output = 11'b01101001110;
        state_var_NS = COMP_LOOP_C_486;
      end
      COMP_LOOP_C_486 : begin
        fsm_output = 11'b01101001111;
        state_var_NS = COMP_LOOP_C_487;
      end
      COMP_LOOP_C_487 : begin
        fsm_output = 11'b01101010000;
        state_var_NS = COMP_LOOP_C_488;
      end
      COMP_LOOP_C_488 : begin
        fsm_output = 11'b01101010001;
        state_var_NS = COMP_LOOP_C_489;
      end
      COMP_LOOP_C_489 : begin
        fsm_output = 11'b01101010010;
        state_var_NS = COMP_LOOP_C_490;
      end
      COMP_LOOP_C_490 : begin
        fsm_output = 11'b01101010011;
        state_var_NS = COMP_LOOP_C_491;
      end
      COMP_LOOP_C_491 : begin
        fsm_output = 11'b01101010100;
        state_var_NS = COMP_LOOP_C_492;
      end
      COMP_LOOP_C_492 : begin
        fsm_output = 11'b01101010101;
        state_var_NS = COMP_LOOP_C_493;
      end
      COMP_LOOP_C_493 : begin
        fsm_output = 11'b01101010110;
        state_var_NS = COMP_LOOP_C_494;
      end
      COMP_LOOP_C_494 : begin
        fsm_output = 11'b01101010111;
        state_var_NS = COMP_LOOP_C_495;
      end
      COMP_LOOP_C_495 : begin
        fsm_output = 11'b01101011000;
        state_var_NS = COMP_LOOP_C_496;
      end
      COMP_LOOP_C_496 : begin
        fsm_output = 11'b01101011001;
        if ( COMP_LOOP_C_496_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_497;
        end
      end
      COMP_LOOP_C_497 : begin
        fsm_output = 11'b01101011010;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_0;
      end
      COMP_LOOP_9_modExp_1_while_C_0 : begin
        fsm_output = 11'b01101011011;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_1;
      end
      COMP_LOOP_9_modExp_1_while_C_1 : begin
        fsm_output = 11'b01101011100;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_2;
      end
      COMP_LOOP_9_modExp_1_while_C_2 : begin
        fsm_output = 11'b01101011101;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_3;
      end
      COMP_LOOP_9_modExp_1_while_C_3 : begin
        fsm_output = 11'b01101011110;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_4;
      end
      COMP_LOOP_9_modExp_1_while_C_4 : begin
        fsm_output = 11'b01101011111;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_5;
      end
      COMP_LOOP_9_modExp_1_while_C_5 : begin
        fsm_output = 11'b01101100000;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_6;
      end
      COMP_LOOP_9_modExp_1_while_C_6 : begin
        fsm_output = 11'b01101100001;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_7;
      end
      COMP_LOOP_9_modExp_1_while_C_7 : begin
        fsm_output = 11'b01101100010;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_8;
      end
      COMP_LOOP_9_modExp_1_while_C_8 : begin
        fsm_output = 11'b01101100011;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_9;
      end
      COMP_LOOP_9_modExp_1_while_C_9 : begin
        fsm_output = 11'b01101100100;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_10;
      end
      COMP_LOOP_9_modExp_1_while_C_10 : begin
        fsm_output = 11'b01101100101;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_11;
      end
      COMP_LOOP_9_modExp_1_while_C_11 : begin
        fsm_output = 11'b01101100110;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_12;
      end
      COMP_LOOP_9_modExp_1_while_C_12 : begin
        fsm_output = 11'b01101100111;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_13;
      end
      COMP_LOOP_9_modExp_1_while_C_13 : begin
        fsm_output = 11'b01101101000;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_14;
      end
      COMP_LOOP_9_modExp_1_while_C_14 : begin
        fsm_output = 11'b01101101001;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_15;
      end
      COMP_LOOP_9_modExp_1_while_C_15 : begin
        fsm_output = 11'b01101101010;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_16;
      end
      COMP_LOOP_9_modExp_1_while_C_16 : begin
        fsm_output = 11'b01101101011;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_17;
      end
      COMP_LOOP_9_modExp_1_while_C_17 : begin
        fsm_output = 11'b01101101100;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_18;
      end
      COMP_LOOP_9_modExp_1_while_C_18 : begin
        fsm_output = 11'b01101101101;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_19;
      end
      COMP_LOOP_9_modExp_1_while_C_19 : begin
        fsm_output = 11'b01101101110;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_20;
      end
      COMP_LOOP_9_modExp_1_while_C_20 : begin
        fsm_output = 11'b01101101111;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_21;
      end
      COMP_LOOP_9_modExp_1_while_C_21 : begin
        fsm_output = 11'b01101110000;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_22;
      end
      COMP_LOOP_9_modExp_1_while_C_22 : begin
        fsm_output = 11'b01101110001;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_23;
      end
      COMP_LOOP_9_modExp_1_while_C_23 : begin
        fsm_output = 11'b01101110010;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_24;
      end
      COMP_LOOP_9_modExp_1_while_C_24 : begin
        fsm_output = 11'b01101110011;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_25;
      end
      COMP_LOOP_9_modExp_1_while_C_25 : begin
        fsm_output = 11'b01101110100;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_26;
      end
      COMP_LOOP_9_modExp_1_while_C_26 : begin
        fsm_output = 11'b01101110101;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_27;
      end
      COMP_LOOP_9_modExp_1_while_C_27 : begin
        fsm_output = 11'b01101110110;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_28;
      end
      COMP_LOOP_9_modExp_1_while_C_28 : begin
        fsm_output = 11'b01101110111;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_29;
      end
      COMP_LOOP_9_modExp_1_while_C_29 : begin
        fsm_output = 11'b01101111000;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_30;
      end
      COMP_LOOP_9_modExp_1_while_C_30 : begin
        fsm_output = 11'b01101111001;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_31;
      end
      COMP_LOOP_9_modExp_1_while_C_31 : begin
        fsm_output = 11'b01101111010;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_32;
      end
      COMP_LOOP_9_modExp_1_while_C_32 : begin
        fsm_output = 11'b01101111011;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_33;
      end
      COMP_LOOP_9_modExp_1_while_C_33 : begin
        fsm_output = 11'b01101111100;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_34;
      end
      COMP_LOOP_9_modExp_1_while_C_34 : begin
        fsm_output = 11'b01101111101;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_35;
      end
      COMP_LOOP_9_modExp_1_while_C_35 : begin
        fsm_output = 11'b01101111110;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_36;
      end
      COMP_LOOP_9_modExp_1_while_C_36 : begin
        fsm_output = 11'b01101111111;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_37;
      end
      COMP_LOOP_9_modExp_1_while_C_37 : begin
        fsm_output = 11'b01110000000;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_38;
      end
      COMP_LOOP_9_modExp_1_while_C_38 : begin
        fsm_output = 11'b01110000001;
        if ( COMP_LOOP_9_modExp_1_while_C_38_tr0 ) begin
          state_var_NS = COMP_LOOP_C_498;
        end
        else begin
          state_var_NS = COMP_LOOP_9_modExp_1_while_C_0;
        end
      end
      COMP_LOOP_C_498 : begin
        fsm_output = 11'b01110000010;
        state_var_NS = COMP_LOOP_C_499;
      end
      COMP_LOOP_C_499 : begin
        fsm_output = 11'b01110000011;
        state_var_NS = COMP_LOOP_C_500;
      end
      COMP_LOOP_C_500 : begin
        fsm_output = 11'b01110000100;
        state_var_NS = COMP_LOOP_C_501;
      end
      COMP_LOOP_C_501 : begin
        fsm_output = 11'b01110000101;
        state_var_NS = COMP_LOOP_C_502;
      end
      COMP_LOOP_C_502 : begin
        fsm_output = 11'b01110000110;
        state_var_NS = COMP_LOOP_C_503;
      end
      COMP_LOOP_C_503 : begin
        fsm_output = 11'b01110000111;
        state_var_NS = COMP_LOOP_C_504;
      end
      COMP_LOOP_C_504 : begin
        fsm_output = 11'b01110001000;
        state_var_NS = COMP_LOOP_C_505;
      end
      COMP_LOOP_C_505 : begin
        fsm_output = 11'b01110001001;
        state_var_NS = COMP_LOOP_C_506;
      end
      COMP_LOOP_C_506 : begin
        fsm_output = 11'b01110001010;
        state_var_NS = COMP_LOOP_C_507;
      end
      COMP_LOOP_C_507 : begin
        fsm_output = 11'b01110001011;
        state_var_NS = COMP_LOOP_C_508;
      end
      COMP_LOOP_C_508 : begin
        fsm_output = 11'b01110001100;
        state_var_NS = COMP_LOOP_C_509;
      end
      COMP_LOOP_C_509 : begin
        fsm_output = 11'b01110001101;
        state_var_NS = COMP_LOOP_C_510;
      end
      COMP_LOOP_C_510 : begin
        fsm_output = 11'b01110001110;
        state_var_NS = COMP_LOOP_C_511;
      end
      COMP_LOOP_C_511 : begin
        fsm_output = 11'b01110001111;
        state_var_NS = COMP_LOOP_C_512;
      end
      COMP_LOOP_C_512 : begin
        fsm_output = 11'b01110010000;
        state_var_NS = COMP_LOOP_C_513;
      end
      COMP_LOOP_C_513 : begin
        fsm_output = 11'b01110010001;
        state_var_NS = COMP_LOOP_C_514;
      end
      COMP_LOOP_C_514 : begin
        fsm_output = 11'b01110010010;
        state_var_NS = COMP_LOOP_C_515;
      end
      COMP_LOOP_C_515 : begin
        fsm_output = 11'b01110010011;
        state_var_NS = COMP_LOOP_C_516;
      end
      COMP_LOOP_C_516 : begin
        fsm_output = 11'b01110010100;
        state_var_NS = COMP_LOOP_C_517;
      end
      COMP_LOOP_C_517 : begin
        fsm_output = 11'b01110010101;
        state_var_NS = COMP_LOOP_C_518;
      end
      COMP_LOOP_C_518 : begin
        fsm_output = 11'b01110010110;
        state_var_NS = COMP_LOOP_C_519;
      end
      COMP_LOOP_C_519 : begin
        fsm_output = 11'b01110010111;
        state_var_NS = COMP_LOOP_C_520;
      end
      COMP_LOOP_C_520 : begin
        fsm_output = 11'b01110011000;
        state_var_NS = COMP_LOOP_C_521;
      end
      COMP_LOOP_C_521 : begin
        fsm_output = 11'b01110011001;
        state_var_NS = COMP_LOOP_C_522;
      end
      COMP_LOOP_C_522 : begin
        fsm_output = 11'b01110011010;
        state_var_NS = COMP_LOOP_C_523;
      end
      COMP_LOOP_C_523 : begin
        fsm_output = 11'b01110011011;
        state_var_NS = COMP_LOOP_C_524;
      end
      COMP_LOOP_C_524 : begin
        fsm_output = 11'b01110011100;
        state_var_NS = COMP_LOOP_C_525;
      end
      COMP_LOOP_C_525 : begin
        fsm_output = 11'b01110011101;
        state_var_NS = COMP_LOOP_C_526;
      end
      COMP_LOOP_C_526 : begin
        fsm_output = 11'b01110011110;
        state_var_NS = COMP_LOOP_C_527;
      end
      COMP_LOOP_C_527 : begin
        fsm_output = 11'b01110011111;
        state_var_NS = COMP_LOOP_C_528;
      end
      COMP_LOOP_C_528 : begin
        fsm_output = 11'b01110100000;
        state_var_NS = COMP_LOOP_C_529;
      end
      COMP_LOOP_C_529 : begin
        fsm_output = 11'b01110100001;
        state_var_NS = COMP_LOOP_C_530;
      end
      COMP_LOOP_C_530 : begin
        fsm_output = 11'b01110100010;
        state_var_NS = COMP_LOOP_C_531;
      end
      COMP_LOOP_C_531 : begin
        fsm_output = 11'b01110100011;
        state_var_NS = COMP_LOOP_C_532;
      end
      COMP_LOOP_C_532 : begin
        fsm_output = 11'b01110100100;
        state_var_NS = COMP_LOOP_C_533;
      end
      COMP_LOOP_C_533 : begin
        fsm_output = 11'b01110100101;
        state_var_NS = COMP_LOOP_C_534;
      end
      COMP_LOOP_C_534 : begin
        fsm_output = 11'b01110100110;
        state_var_NS = COMP_LOOP_C_535;
      end
      COMP_LOOP_C_535 : begin
        fsm_output = 11'b01110100111;
        state_var_NS = COMP_LOOP_C_536;
      end
      COMP_LOOP_C_536 : begin
        fsm_output = 11'b01110101000;
        state_var_NS = COMP_LOOP_C_537;
      end
      COMP_LOOP_C_537 : begin
        fsm_output = 11'b01110101001;
        state_var_NS = COMP_LOOP_C_538;
      end
      COMP_LOOP_C_538 : begin
        fsm_output = 11'b01110101010;
        state_var_NS = COMP_LOOP_C_539;
      end
      COMP_LOOP_C_539 : begin
        fsm_output = 11'b01110101011;
        state_var_NS = COMP_LOOP_C_540;
      end
      COMP_LOOP_C_540 : begin
        fsm_output = 11'b01110101100;
        state_var_NS = COMP_LOOP_C_541;
      end
      COMP_LOOP_C_541 : begin
        fsm_output = 11'b01110101101;
        state_var_NS = COMP_LOOP_C_542;
      end
      COMP_LOOP_C_542 : begin
        fsm_output = 11'b01110101110;
        state_var_NS = COMP_LOOP_C_543;
      end
      COMP_LOOP_C_543 : begin
        fsm_output = 11'b01110101111;
        state_var_NS = COMP_LOOP_C_544;
      end
      COMP_LOOP_C_544 : begin
        fsm_output = 11'b01110110000;
        state_var_NS = COMP_LOOP_C_545;
      end
      COMP_LOOP_C_545 : begin
        fsm_output = 11'b01110110001;
        state_var_NS = COMP_LOOP_C_546;
      end
      COMP_LOOP_C_546 : begin
        fsm_output = 11'b01110110010;
        state_var_NS = COMP_LOOP_C_547;
      end
      COMP_LOOP_C_547 : begin
        fsm_output = 11'b01110110011;
        state_var_NS = COMP_LOOP_C_548;
      end
      COMP_LOOP_C_548 : begin
        fsm_output = 11'b01110110100;
        state_var_NS = COMP_LOOP_C_549;
      end
      COMP_LOOP_C_549 : begin
        fsm_output = 11'b01110110101;
        state_var_NS = COMP_LOOP_C_550;
      end
      COMP_LOOP_C_550 : begin
        fsm_output = 11'b01110110110;
        state_var_NS = COMP_LOOP_C_551;
      end
      COMP_LOOP_C_551 : begin
        fsm_output = 11'b01110110111;
        state_var_NS = COMP_LOOP_C_552;
      end
      COMP_LOOP_C_552 : begin
        fsm_output = 11'b01110111000;
        state_var_NS = COMP_LOOP_C_553;
      end
      COMP_LOOP_C_553 : begin
        fsm_output = 11'b01110111001;
        state_var_NS = COMP_LOOP_C_554;
      end
      COMP_LOOP_C_554 : begin
        fsm_output = 11'b01110111010;
        state_var_NS = COMP_LOOP_C_555;
      end
      COMP_LOOP_C_555 : begin
        fsm_output = 11'b01110111011;
        state_var_NS = COMP_LOOP_C_556;
      end
      COMP_LOOP_C_556 : begin
        fsm_output = 11'b01110111100;
        state_var_NS = COMP_LOOP_C_557;
      end
      COMP_LOOP_C_557 : begin
        fsm_output = 11'b01110111101;
        state_var_NS = COMP_LOOP_C_558;
      end
      COMP_LOOP_C_558 : begin
        fsm_output = 11'b01110111110;
        if ( COMP_LOOP_C_558_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_559;
        end
      end
      COMP_LOOP_C_559 : begin
        fsm_output = 11'b01110111111;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_0;
      end
      COMP_LOOP_10_modExp_1_while_C_0 : begin
        fsm_output = 11'b01111000000;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_1;
      end
      COMP_LOOP_10_modExp_1_while_C_1 : begin
        fsm_output = 11'b01111000001;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_2;
      end
      COMP_LOOP_10_modExp_1_while_C_2 : begin
        fsm_output = 11'b01111000010;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_3;
      end
      COMP_LOOP_10_modExp_1_while_C_3 : begin
        fsm_output = 11'b01111000011;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_4;
      end
      COMP_LOOP_10_modExp_1_while_C_4 : begin
        fsm_output = 11'b01111000100;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_5;
      end
      COMP_LOOP_10_modExp_1_while_C_5 : begin
        fsm_output = 11'b01111000101;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_6;
      end
      COMP_LOOP_10_modExp_1_while_C_6 : begin
        fsm_output = 11'b01111000110;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_7;
      end
      COMP_LOOP_10_modExp_1_while_C_7 : begin
        fsm_output = 11'b01111000111;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_8;
      end
      COMP_LOOP_10_modExp_1_while_C_8 : begin
        fsm_output = 11'b01111001000;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_9;
      end
      COMP_LOOP_10_modExp_1_while_C_9 : begin
        fsm_output = 11'b01111001001;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_10;
      end
      COMP_LOOP_10_modExp_1_while_C_10 : begin
        fsm_output = 11'b01111001010;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_11;
      end
      COMP_LOOP_10_modExp_1_while_C_11 : begin
        fsm_output = 11'b01111001011;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_12;
      end
      COMP_LOOP_10_modExp_1_while_C_12 : begin
        fsm_output = 11'b01111001100;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_13;
      end
      COMP_LOOP_10_modExp_1_while_C_13 : begin
        fsm_output = 11'b01111001101;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_14;
      end
      COMP_LOOP_10_modExp_1_while_C_14 : begin
        fsm_output = 11'b01111001110;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_15;
      end
      COMP_LOOP_10_modExp_1_while_C_15 : begin
        fsm_output = 11'b01111001111;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_16;
      end
      COMP_LOOP_10_modExp_1_while_C_16 : begin
        fsm_output = 11'b01111010000;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_17;
      end
      COMP_LOOP_10_modExp_1_while_C_17 : begin
        fsm_output = 11'b01111010001;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_18;
      end
      COMP_LOOP_10_modExp_1_while_C_18 : begin
        fsm_output = 11'b01111010010;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_19;
      end
      COMP_LOOP_10_modExp_1_while_C_19 : begin
        fsm_output = 11'b01111010011;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_20;
      end
      COMP_LOOP_10_modExp_1_while_C_20 : begin
        fsm_output = 11'b01111010100;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_21;
      end
      COMP_LOOP_10_modExp_1_while_C_21 : begin
        fsm_output = 11'b01111010101;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_22;
      end
      COMP_LOOP_10_modExp_1_while_C_22 : begin
        fsm_output = 11'b01111010110;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_23;
      end
      COMP_LOOP_10_modExp_1_while_C_23 : begin
        fsm_output = 11'b01111010111;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_24;
      end
      COMP_LOOP_10_modExp_1_while_C_24 : begin
        fsm_output = 11'b01111011000;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_25;
      end
      COMP_LOOP_10_modExp_1_while_C_25 : begin
        fsm_output = 11'b01111011001;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_26;
      end
      COMP_LOOP_10_modExp_1_while_C_26 : begin
        fsm_output = 11'b01111011010;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_27;
      end
      COMP_LOOP_10_modExp_1_while_C_27 : begin
        fsm_output = 11'b01111011011;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_28;
      end
      COMP_LOOP_10_modExp_1_while_C_28 : begin
        fsm_output = 11'b01111011100;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_29;
      end
      COMP_LOOP_10_modExp_1_while_C_29 : begin
        fsm_output = 11'b01111011101;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_30;
      end
      COMP_LOOP_10_modExp_1_while_C_30 : begin
        fsm_output = 11'b01111011110;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_31;
      end
      COMP_LOOP_10_modExp_1_while_C_31 : begin
        fsm_output = 11'b01111011111;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_32;
      end
      COMP_LOOP_10_modExp_1_while_C_32 : begin
        fsm_output = 11'b01111100000;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_33;
      end
      COMP_LOOP_10_modExp_1_while_C_33 : begin
        fsm_output = 11'b01111100001;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_34;
      end
      COMP_LOOP_10_modExp_1_while_C_34 : begin
        fsm_output = 11'b01111100010;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_35;
      end
      COMP_LOOP_10_modExp_1_while_C_35 : begin
        fsm_output = 11'b01111100011;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_36;
      end
      COMP_LOOP_10_modExp_1_while_C_36 : begin
        fsm_output = 11'b01111100100;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_37;
      end
      COMP_LOOP_10_modExp_1_while_C_37 : begin
        fsm_output = 11'b01111100101;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_38;
      end
      COMP_LOOP_10_modExp_1_while_C_38 : begin
        fsm_output = 11'b01111100110;
        if ( COMP_LOOP_10_modExp_1_while_C_38_tr0 ) begin
          state_var_NS = COMP_LOOP_C_560;
        end
        else begin
          state_var_NS = COMP_LOOP_10_modExp_1_while_C_0;
        end
      end
      COMP_LOOP_C_560 : begin
        fsm_output = 11'b01111100111;
        state_var_NS = COMP_LOOP_C_561;
      end
      COMP_LOOP_C_561 : begin
        fsm_output = 11'b01111101000;
        state_var_NS = COMP_LOOP_C_562;
      end
      COMP_LOOP_C_562 : begin
        fsm_output = 11'b01111101001;
        state_var_NS = COMP_LOOP_C_563;
      end
      COMP_LOOP_C_563 : begin
        fsm_output = 11'b01111101010;
        state_var_NS = COMP_LOOP_C_564;
      end
      COMP_LOOP_C_564 : begin
        fsm_output = 11'b01111101011;
        state_var_NS = COMP_LOOP_C_565;
      end
      COMP_LOOP_C_565 : begin
        fsm_output = 11'b01111101100;
        state_var_NS = COMP_LOOP_C_566;
      end
      COMP_LOOP_C_566 : begin
        fsm_output = 11'b01111101101;
        state_var_NS = COMP_LOOP_C_567;
      end
      COMP_LOOP_C_567 : begin
        fsm_output = 11'b01111101110;
        state_var_NS = COMP_LOOP_C_568;
      end
      COMP_LOOP_C_568 : begin
        fsm_output = 11'b01111101111;
        state_var_NS = COMP_LOOP_C_569;
      end
      COMP_LOOP_C_569 : begin
        fsm_output = 11'b01111110000;
        state_var_NS = COMP_LOOP_C_570;
      end
      COMP_LOOP_C_570 : begin
        fsm_output = 11'b01111110001;
        state_var_NS = COMP_LOOP_C_571;
      end
      COMP_LOOP_C_571 : begin
        fsm_output = 11'b01111110010;
        state_var_NS = COMP_LOOP_C_572;
      end
      COMP_LOOP_C_572 : begin
        fsm_output = 11'b01111110011;
        state_var_NS = COMP_LOOP_C_573;
      end
      COMP_LOOP_C_573 : begin
        fsm_output = 11'b01111110100;
        state_var_NS = COMP_LOOP_C_574;
      end
      COMP_LOOP_C_574 : begin
        fsm_output = 11'b01111110101;
        state_var_NS = COMP_LOOP_C_575;
      end
      COMP_LOOP_C_575 : begin
        fsm_output = 11'b01111110110;
        state_var_NS = COMP_LOOP_C_576;
      end
      COMP_LOOP_C_576 : begin
        fsm_output = 11'b01111110111;
        state_var_NS = COMP_LOOP_C_577;
      end
      COMP_LOOP_C_577 : begin
        fsm_output = 11'b01111111000;
        state_var_NS = COMP_LOOP_C_578;
      end
      COMP_LOOP_C_578 : begin
        fsm_output = 11'b01111111001;
        state_var_NS = COMP_LOOP_C_579;
      end
      COMP_LOOP_C_579 : begin
        fsm_output = 11'b01111111010;
        state_var_NS = COMP_LOOP_C_580;
      end
      COMP_LOOP_C_580 : begin
        fsm_output = 11'b01111111011;
        state_var_NS = COMP_LOOP_C_581;
      end
      COMP_LOOP_C_581 : begin
        fsm_output = 11'b01111111100;
        state_var_NS = COMP_LOOP_C_582;
      end
      COMP_LOOP_C_582 : begin
        fsm_output = 11'b01111111101;
        state_var_NS = COMP_LOOP_C_583;
      end
      COMP_LOOP_C_583 : begin
        fsm_output = 11'b01111111110;
        state_var_NS = COMP_LOOP_C_584;
      end
      COMP_LOOP_C_584 : begin
        fsm_output = 11'b01111111111;
        state_var_NS = COMP_LOOP_C_585;
      end
      COMP_LOOP_C_585 : begin
        fsm_output = 11'b10000000000;
        state_var_NS = COMP_LOOP_C_586;
      end
      COMP_LOOP_C_586 : begin
        fsm_output = 11'b10000000001;
        state_var_NS = COMP_LOOP_C_587;
      end
      COMP_LOOP_C_587 : begin
        fsm_output = 11'b10000000010;
        state_var_NS = COMP_LOOP_C_588;
      end
      COMP_LOOP_C_588 : begin
        fsm_output = 11'b10000000011;
        state_var_NS = COMP_LOOP_C_589;
      end
      COMP_LOOP_C_589 : begin
        fsm_output = 11'b10000000100;
        state_var_NS = COMP_LOOP_C_590;
      end
      COMP_LOOP_C_590 : begin
        fsm_output = 11'b10000000101;
        state_var_NS = COMP_LOOP_C_591;
      end
      COMP_LOOP_C_591 : begin
        fsm_output = 11'b10000000110;
        state_var_NS = COMP_LOOP_C_592;
      end
      COMP_LOOP_C_592 : begin
        fsm_output = 11'b10000000111;
        state_var_NS = COMP_LOOP_C_593;
      end
      COMP_LOOP_C_593 : begin
        fsm_output = 11'b10000001000;
        state_var_NS = COMP_LOOP_C_594;
      end
      COMP_LOOP_C_594 : begin
        fsm_output = 11'b10000001001;
        state_var_NS = COMP_LOOP_C_595;
      end
      COMP_LOOP_C_595 : begin
        fsm_output = 11'b10000001010;
        state_var_NS = COMP_LOOP_C_596;
      end
      COMP_LOOP_C_596 : begin
        fsm_output = 11'b10000001011;
        state_var_NS = COMP_LOOP_C_597;
      end
      COMP_LOOP_C_597 : begin
        fsm_output = 11'b10000001100;
        state_var_NS = COMP_LOOP_C_598;
      end
      COMP_LOOP_C_598 : begin
        fsm_output = 11'b10000001101;
        state_var_NS = COMP_LOOP_C_599;
      end
      COMP_LOOP_C_599 : begin
        fsm_output = 11'b10000001110;
        state_var_NS = COMP_LOOP_C_600;
      end
      COMP_LOOP_C_600 : begin
        fsm_output = 11'b10000001111;
        state_var_NS = COMP_LOOP_C_601;
      end
      COMP_LOOP_C_601 : begin
        fsm_output = 11'b10000010000;
        state_var_NS = COMP_LOOP_C_602;
      end
      COMP_LOOP_C_602 : begin
        fsm_output = 11'b10000010001;
        state_var_NS = COMP_LOOP_C_603;
      end
      COMP_LOOP_C_603 : begin
        fsm_output = 11'b10000010010;
        state_var_NS = COMP_LOOP_C_604;
      end
      COMP_LOOP_C_604 : begin
        fsm_output = 11'b10000010011;
        state_var_NS = COMP_LOOP_C_605;
      end
      COMP_LOOP_C_605 : begin
        fsm_output = 11'b10000010100;
        state_var_NS = COMP_LOOP_C_606;
      end
      COMP_LOOP_C_606 : begin
        fsm_output = 11'b10000010101;
        state_var_NS = COMP_LOOP_C_607;
      end
      COMP_LOOP_C_607 : begin
        fsm_output = 11'b10000010110;
        state_var_NS = COMP_LOOP_C_608;
      end
      COMP_LOOP_C_608 : begin
        fsm_output = 11'b10000010111;
        state_var_NS = COMP_LOOP_C_609;
      end
      COMP_LOOP_C_609 : begin
        fsm_output = 11'b10000011000;
        state_var_NS = COMP_LOOP_C_610;
      end
      COMP_LOOP_C_610 : begin
        fsm_output = 11'b10000011001;
        state_var_NS = COMP_LOOP_C_611;
      end
      COMP_LOOP_C_611 : begin
        fsm_output = 11'b10000011010;
        state_var_NS = COMP_LOOP_C_612;
      end
      COMP_LOOP_C_612 : begin
        fsm_output = 11'b10000011011;
        state_var_NS = COMP_LOOP_C_613;
      end
      COMP_LOOP_C_613 : begin
        fsm_output = 11'b10000011100;
        state_var_NS = COMP_LOOP_C_614;
      end
      COMP_LOOP_C_614 : begin
        fsm_output = 11'b10000011101;
        state_var_NS = COMP_LOOP_C_615;
      end
      COMP_LOOP_C_615 : begin
        fsm_output = 11'b10000011110;
        state_var_NS = COMP_LOOP_C_616;
      end
      COMP_LOOP_C_616 : begin
        fsm_output = 11'b10000011111;
        state_var_NS = COMP_LOOP_C_617;
      end
      COMP_LOOP_C_617 : begin
        fsm_output = 11'b10000100000;
        state_var_NS = COMP_LOOP_C_618;
      end
      COMP_LOOP_C_618 : begin
        fsm_output = 11'b10000100001;
        state_var_NS = COMP_LOOP_C_619;
      end
      COMP_LOOP_C_619 : begin
        fsm_output = 11'b10000100010;
        state_var_NS = COMP_LOOP_C_620;
      end
      COMP_LOOP_C_620 : begin
        fsm_output = 11'b10000100011;
        if ( COMP_LOOP_C_620_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_621;
        end
      end
      COMP_LOOP_C_621 : begin
        fsm_output = 11'b10000100100;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_0;
      end
      COMP_LOOP_11_modExp_1_while_C_0 : begin
        fsm_output = 11'b10000100101;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_1;
      end
      COMP_LOOP_11_modExp_1_while_C_1 : begin
        fsm_output = 11'b10000100110;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_2;
      end
      COMP_LOOP_11_modExp_1_while_C_2 : begin
        fsm_output = 11'b10000100111;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_3;
      end
      COMP_LOOP_11_modExp_1_while_C_3 : begin
        fsm_output = 11'b10000101000;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_4;
      end
      COMP_LOOP_11_modExp_1_while_C_4 : begin
        fsm_output = 11'b10000101001;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_5;
      end
      COMP_LOOP_11_modExp_1_while_C_5 : begin
        fsm_output = 11'b10000101010;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_6;
      end
      COMP_LOOP_11_modExp_1_while_C_6 : begin
        fsm_output = 11'b10000101011;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_7;
      end
      COMP_LOOP_11_modExp_1_while_C_7 : begin
        fsm_output = 11'b10000101100;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_8;
      end
      COMP_LOOP_11_modExp_1_while_C_8 : begin
        fsm_output = 11'b10000101101;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_9;
      end
      COMP_LOOP_11_modExp_1_while_C_9 : begin
        fsm_output = 11'b10000101110;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_10;
      end
      COMP_LOOP_11_modExp_1_while_C_10 : begin
        fsm_output = 11'b10000101111;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_11;
      end
      COMP_LOOP_11_modExp_1_while_C_11 : begin
        fsm_output = 11'b10000110000;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_12;
      end
      COMP_LOOP_11_modExp_1_while_C_12 : begin
        fsm_output = 11'b10000110001;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_13;
      end
      COMP_LOOP_11_modExp_1_while_C_13 : begin
        fsm_output = 11'b10000110010;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_14;
      end
      COMP_LOOP_11_modExp_1_while_C_14 : begin
        fsm_output = 11'b10000110011;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_15;
      end
      COMP_LOOP_11_modExp_1_while_C_15 : begin
        fsm_output = 11'b10000110100;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_16;
      end
      COMP_LOOP_11_modExp_1_while_C_16 : begin
        fsm_output = 11'b10000110101;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_17;
      end
      COMP_LOOP_11_modExp_1_while_C_17 : begin
        fsm_output = 11'b10000110110;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_18;
      end
      COMP_LOOP_11_modExp_1_while_C_18 : begin
        fsm_output = 11'b10000110111;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_19;
      end
      COMP_LOOP_11_modExp_1_while_C_19 : begin
        fsm_output = 11'b10000111000;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_20;
      end
      COMP_LOOP_11_modExp_1_while_C_20 : begin
        fsm_output = 11'b10000111001;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_21;
      end
      COMP_LOOP_11_modExp_1_while_C_21 : begin
        fsm_output = 11'b10000111010;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_22;
      end
      COMP_LOOP_11_modExp_1_while_C_22 : begin
        fsm_output = 11'b10000111011;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_23;
      end
      COMP_LOOP_11_modExp_1_while_C_23 : begin
        fsm_output = 11'b10000111100;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_24;
      end
      COMP_LOOP_11_modExp_1_while_C_24 : begin
        fsm_output = 11'b10000111101;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_25;
      end
      COMP_LOOP_11_modExp_1_while_C_25 : begin
        fsm_output = 11'b10000111110;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_26;
      end
      COMP_LOOP_11_modExp_1_while_C_26 : begin
        fsm_output = 11'b10000111111;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_27;
      end
      COMP_LOOP_11_modExp_1_while_C_27 : begin
        fsm_output = 11'b10001000000;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_28;
      end
      COMP_LOOP_11_modExp_1_while_C_28 : begin
        fsm_output = 11'b10001000001;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_29;
      end
      COMP_LOOP_11_modExp_1_while_C_29 : begin
        fsm_output = 11'b10001000010;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_30;
      end
      COMP_LOOP_11_modExp_1_while_C_30 : begin
        fsm_output = 11'b10001000011;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_31;
      end
      COMP_LOOP_11_modExp_1_while_C_31 : begin
        fsm_output = 11'b10001000100;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_32;
      end
      COMP_LOOP_11_modExp_1_while_C_32 : begin
        fsm_output = 11'b10001000101;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_33;
      end
      COMP_LOOP_11_modExp_1_while_C_33 : begin
        fsm_output = 11'b10001000110;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_34;
      end
      COMP_LOOP_11_modExp_1_while_C_34 : begin
        fsm_output = 11'b10001000111;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_35;
      end
      COMP_LOOP_11_modExp_1_while_C_35 : begin
        fsm_output = 11'b10001001000;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_36;
      end
      COMP_LOOP_11_modExp_1_while_C_36 : begin
        fsm_output = 11'b10001001001;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_37;
      end
      COMP_LOOP_11_modExp_1_while_C_37 : begin
        fsm_output = 11'b10001001010;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_38;
      end
      COMP_LOOP_11_modExp_1_while_C_38 : begin
        fsm_output = 11'b10001001011;
        if ( COMP_LOOP_11_modExp_1_while_C_38_tr0 ) begin
          state_var_NS = COMP_LOOP_C_622;
        end
        else begin
          state_var_NS = COMP_LOOP_11_modExp_1_while_C_0;
        end
      end
      COMP_LOOP_C_622 : begin
        fsm_output = 11'b10001001100;
        state_var_NS = COMP_LOOP_C_623;
      end
      COMP_LOOP_C_623 : begin
        fsm_output = 11'b10001001101;
        state_var_NS = COMP_LOOP_C_624;
      end
      COMP_LOOP_C_624 : begin
        fsm_output = 11'b10001001110;
        state_var_NS = COMP_LOOP_C_625;
      end
      COMP_LOOP_C_625 : begin
        fsm_output = 11'b10001001111;
        state_var_NS = COMP_LOOP_C_626;
      end
      COMP_LOOP_C_626 : begin
        fsm_output = 11'b10001010000;
        state_var_NS = COMP_LOOP_C_627;
      end
      COMP_LOOP_C_627 : begin
        fsm_output = 11'b10001010001;
        state_var_NS = COMP_LOOP_C_628;
      end
      COMP_LOOP_C_628 : begin
        fsm_output = 11'b10001010010;
        state_var_NS = COMP_LOOP_C_629;
      end
      COMP_LOOP_C_629 : begin
        fsm_output = 11'b10001010011;
        state_var_NS = COMP_LOOP_C_630;
      end
      COMP_LOOP_C_630 : begin
        fsm_output = 11'b10001010100;
        state_var_NS = COMP_LOOP_C_631;
      end
      COMP_LOOP_C_631 : begin
        fsm_output = 11'b10001010101;
        state_var_NS = COMP_LOOP_C_632;
      end
      COMP_LOOP_C_632 : begin
        fsm_output = 11'b10001010110;
        state_var_NS = COMP_LOOP_C_633;
      end
      COMP_LOOP_C_633 : begin
        fsm_output = 11'b10001010111;
        state_var_NS = COMP_LOOP_C_634;
      end
      COMP_LOOP_C_634 : begin
        fsm_output = 11'b10001011000;
        state_var_NS = COMP_LOOP_C_635;
      end
      COMP_LOOP_C_635 : begin
        fsm_output = 11'b10001011001;
        state_var_NS = COMP_LOOP_C_636;
      end
      COMP_LOOP_C_636 : begin
        fsm_output = 11'b10001011010;
        state_var_NS = COMP_LOOP_C_637;
      end
      COMP_LOOP_C_637 : begin
        fsm_output = 11'b10001011011;
        state_var_NS = COMP_LOOP_C_638;
      end
      COMP_LOOP_C_638 : begin
        fsm_output = 11'b10001011100;
        state_var_NS = COMP_LOOP_C_639;
      end
      COMP_LOOP_C_639 : begin
        fsm_output = 11'b10001011101;
        state_var_NS = COMP_LOOP_C_640;
      end
      COMP_LOOP_C_640 : begin
        fsm_output = 11'b10001011110;
        state_var_NS = COMP_LOOP_C_641;
      end
      COMP_LOOP_C_641 : begin
        fsm_output = 11'b10001011111;
        state_var_NS = COMP_LOOP_C_642;
      end
      COMP_LOOP_C_642 : begin
        fsm_output = 11'b10001100000;
        state_var_NS = COMP_LOOP_C_643;
      end
      COMP_LOOP_C_643 : begin
        fsm_output = 11'b10001100001;
        state_var_NS = COMP_LOOP_C_644;
      end
      COMP_LOOP_C_644 : begin
        fsm_output = 11'b10001100010;
        state_var_NS = COMP_LOOP_C_645;
      end
      COMP_LOOP_C_645 : begin
        fsm_output = 11'b10001100011;
        state_var_NS = COMP_LOOP_C_646;
      end
      COMP_LOOP_C_646 : begin
        fsm_output = 11'b10001100100;
        state_var_NS = COMP_LOOP_C_647;
      end
      COMP_LOOP_C_647 : begin
        fsm_output = 11'b10001100101;
        state_var_NS = COMP_LOOP_C_648;
      end
      COMP_LOOP_C_648 : begin
        fsm_output = 11'b10001100110;
        state_var_NS = COMP_LOOP_C_649;
      end
      COMP_LOOP_C_649 : begin
        fsm_output = 11'b10001100111;
        state_var_NS = COMP_LOOP_C_650;
      end
      COMP_LOOP_C_650 : begin
        fsm_output = 11'b10001101000;
        state_var_NS = COMP_LOOP_C_651;
      end
      COMP_LOOP_C_651 : begin
        fsm_output = 11'b10001101001;
        state_var_NS = COMP_LOOP_C_652;
      end
      COMP_LOOP_C_652 : begin
        fsm_output = 11'b10001101010;
        state_var_NS = COMP_LOOP_C_653;
      end
      COMP_LOOP_C_653 : begin
        fsm_output = 11'b10001101011;
        state_var_NS = COMP_LOOP_C_654;
      end
      COMP_LOOP_C_654 : begin
        fsm_output = 11'b10001101100;
        state_var_NS = COMP_LOOP_C_655;
      end
      COMP_LOOP_C_655 : begin
        fsm_output = 11'b10001101101;
        state_var_NS = COMP_LOOP_C_656;
      end
      COMP_LOOP_C_656 : begin
        fsm_output = 11'b10001101110;
        state_var_NS = COMP_LOOP_C_657;
      end
      COMP_LOOP_C_657 : begin
        fsm_output = 11'b10001101111;
        state_var_NS = COMP_LOOP_C_658;
      end
      COMP_LOOP_C_658 : begin
        fsm_output = 11'b10001110000;
        state_var_NS = COMP_LOOP_C_659;
      end
      COMP_LOOP_C_659 : begin
        fsm_output = 11'b10001110001;
        state_var_NS = COMP_LOOP_C_660;
      end
      COMP_LOOP_C_660 : begin
        fsm_output = 11'b10001110010;
        state_var_NS = COMP_LOOP_C_661;
      end
      COMP_LOOP_C_661 : begin
        fsm_output = 11'b10001110011;
        state_var_NS = COMP_LOOP_C_662;
      end
      COMP_LOOP_C_662 : begin
        fsm_output = 11'b10001110100;
        state_var_NS = COMP_LOOP_C_663;
      end
      COMP_LOOP_C_663 : begin
        fsm_output = 11'b10001110101;
        state_var_NS = COMP_LOOP_C_664;
      end
      COMP_LOOP_C_664 : begin
        fsm_output = 11'b10001110110;
        state_var_NS = COMP_LOOP_C_665;
      end
      COMP_LOOP_C_665 : begin
        fsm_output = 11'b10001110111;
        state_var_NS = COMP_LOOP_C_666;
      end
      COMP_LOOP_C_666 : begin
        fsm_output = 11'b10001111000;
        state_var_NS = COMP_LOOP_C_667;
      end
      COMP_LOOP_C_667 : begin
        fsm_output = 11'b10001111001;
        state_var_NS = COMP_LOOP_C_668;
      end
      COMP_LOOP_C_668 : begin
        fsm_output = 11'b10001111010;
        state_var_NS = COMP_LOOP_C_669;
      end
      COMP_LOOP_C_669 : begin
        fsm_output = 11'b10001111011;
        state_var_NS = COMP_LOOP_C_670;
      end
      COMP_LOOP_C_670 : begin
        fsm_output = 11'b10001111100;
        state_var_NS = COMP_LOOP_C_671;
      end
      COMP_LOOP_C_671 : begin
        fsm_output = 11'b10001111101;
        state_var_NS = COMP_LOOP_C_672;
      end
      COMP_LOOP_C_672 : begin
        fsm_output = 11'b10001111110;
        state_var_NS = COMP_LOOP_C_673;
      end
      COMP_LOOP_C_673 : begin
        fsm_output = 11'b10001111111;
        state_var_NS = COMP_LOOP_C_674;
      end
      COMP_LOOP_C_674 : begin
        fsm_output = 11'b10010000000;
        state_var_NS = COMP_LOOP_C_675;
      end
      COMP_LOOP_C_675 : begin
        fsm_output = 11'b10010000001;
        state_var_NS = COMP_LOOP_C_676;
      end
      COMP_LOOP_C_676 : begin
        fsm_output = 11'b10010000010;
        state_var_NS = COMP_LOOP_C_677;
      end
      COMP_LOOP_C_677 : begin
        fsm_output = 11'b10010000011;
        state_var_NS = COMP_LOOP_C_678;
      end
      COMP_LOOP_C_678 : begin
        fsm_output = 11'b10010000100;
        state_var_NS = COMP_LOOP_C_679;
      end
      COMP_LOOP_C_679 : begin
        fsm_output = 11'b10010000101;
        state_var_NS = COMP_LOOP_C_680;
      end
      COMP_LOOP_C_680 : begin
        fsm_output = 11'b10010000110;
        state_var_NS = COMP_LOOP_C_681;
      end
      COMP_LOOP_C_681 : begin
        fsm_output = 11'b10010000111;
        state_var_NS = COMP_LOOP_C_682;
      end
      COMP_LOOP_C_682 : begin
        fsm_output = 11'b10010001000;
        if ( COMP_LOOP_C_682_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_683;
        end
      end
      COMP_LOOP_C_683 : begin
        fsm_output = 11'b10010001001;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_0;
      end
      COMP_LOOP_12_modExp_1_while_C_0 : begin
        fsm_output = 11'b10010001010;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_1;
      end
      COMP_LOOP_12_modExp_1_while_C_1 : begin
        fsm_output = 11'b10010001011;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_2;
      end
      COMP_LOOP_12_modExp_1_while_C_2 : begin
        fsm_output = 11'b10010001100;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_3;
      end
      COMP_LOOP_12_modExp_1_while_C_3 : begin
        fsm_output = 11'b10010001101;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_4;
      end
      COMP_LOOP_12_modExp_1_while_C_4 : begin
        fsm_output = 11'b10010001110;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_5;
      end
      COMP_LOOP_12_modExp_1_while_C_5 : begin
        fsm_output = 11'b10010001111;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_6;
      end
      COMP_LOOP_12_modExp_1_while_C_6 : begin
        fsm_output = 11'b10010010000;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_7;
      end
      COMP_LOOP_12_modExp_1_while_C_7 : begin
        fsm_output = 11'b10010010001;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_8;
      end
      COMP_LOOP_12_modExp_1_while_C_8 : begin
        fsm_output = 11'b10010010010;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_9;
      end
      COMP_LOOP_12_modExp_1_while_C_9 : begin
        fsm_output = 11'b10010010011;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_10;
      end
      COMP_LOOP_12_modExp_1_while_C_10 : begin
        fsm_output = 11'b10010010100;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_11;
      end
      COMP_LOOP_12_modExp_1_while_C_11 : begin
        fsm_output = 11'b10010010101;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_12;
      end
      COMP_LOOP_12_modExp_1_while_C_12 : begin
        fsm_output = 11'b10010010110;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_13;
      end
      COMP_LOOP_12_modExp_1_while_C_13 : begin
        fsm_output = 11'b10010010111;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_14;
      end
      COMP_LOOP_12_modExp_1_while_C_14 : begin
        fsm_output = 11'b10010011000;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_15;
      end
      COMP_LOOP_12_modExp_1_while_C_15 : begin
        fsm_output = 11'b10010011001;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_16;
      end
      COMP_LOOP_12_modExp_1_while_C_16 : begin
        fsm_output = 11'b10010011010;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_17;
      end
      COMP_LOOP_12_modExp_1_while_C_17 : begin
        fsm_output = 11'b10010011011;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_18;
      end
      COMP_LOOP_12_modExp_1_while_C_18 : begin
        fsm_output = 11'b10010011100;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_19;
      end
      COMP_LOOP_12_modExp_1_while_C_19 : begin
        fsm_output = 11'b10010011101;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_20;
      end
      COMP_LOOP_12_modExp_1_while_C_20 : begin
        fsm_output = 11'b10010011110;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_21;
      end
      COMP_LOOP_12_modExp_1_while_C_21 : begin
        fsm_output = 11'b10010011111;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_22;
      end
      COMP_LOOP_12_modExp_1_while_C_22 : begin
        fsm_output = 11'b10010100000;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_23;
      end
      COMP_LOOP_12_modExp_1_while_C_23 : begin
        fsm_output = 11'b10010100001;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_24;
      end
      COMP_LOOP_12_modExp_1_while_C_24 : begin
        fsm_output = 11'b10010100010;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_25;
      end
      COMP_LOOP_12_modExp_1_while_C_25 : begin
        fsm_output = 11'b10010100011;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_26;
      end
      COMP_LOOP_12_modExp_1_while_C_26 : begin
        fsm_output = 11'b10010100100;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_27;
      end
      COMP_LOOP_12_modExp_1_while_C_27 : begin
        fsm_output = 11'b10010100101;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_28;
      end
      COMP_LOOP_12_modExp_1_while_C_28 : begin
        fsm_output = 11'b10010100110;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_29;
      end
      COMP_LOOP_12_modExp_1_while_C_29 : begin
        fsm_output = 11'b10010100111;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_30;
      end
      COMP_LOOP_12_modExp_1_while_C_30 : begin
        fsm_output = 11'b10010101000;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_31;
      end
      COMP_LOOP_12_modExp_1_while_C_31 : begin
        fsm_output = 11'b10010101001;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_32;
      end
      COMP_LOOP_12_modExp_1_while_C_32 : begin
        fsm_output = 11'b10010101010;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_33;
      end
      COMP_LOOP_12_modExp_1_while_C_33 : begin
        fsm_output = 11'b10010101011;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_34;
      end
      COMP_LOOP_12_modExp_1_while_C_34 : begin
        fsm_output = 11'b10010101100;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_35;
      end
      COMP_LOOP_12_modExp_1_while_C_35 : begin
        fsm_output = 11'b10010101101;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_36;
      end
      COMP_LOOP_12_modExp_1_while_C_36 : begin
        fsm_output = 11'b10010101110;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_37;
      end
      COMP_LOOP_12_modExp_1_while_C_37 : begin
        fsm_output = 11'b10010101111;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_38;
      end
      COMP_LOOP_12_modExp_1_while_C_38 : begin
        fsm_output = 11'b10010110000;
        if ( COMP_LOOP_12_modExp_1_while_C_38_tr0 ) begin
          state_var_NS = COMP_LOOP_C_684;
        end
        else begin
          state_var_NS = COMP_LOOP_12_modExp_1_while_C_0;
        end
      end
      COMP_LOOP_C_684 : begin
        fsm_output = 11'b10010110001;
        state_var_NS = COMP_LOOP_C_685;
      end
      COMP_LOOP_C_685 : begin
        fsm_output = 11'b10010110010;
        state_var_NS = COMP_LOOP_C_686;
      end
      COMP_LOOP_C_686 : begin
        fsm_output = 11'b10010110011;
        state_var_NS = COMP_LOOP_C_687;
      end
      COMP_LOOP_C_687 : begin
        fsm_output = 11'b10010110100;
        state_var_NS = COMP_LOOP_C_688;
      end
      COMP_LOOP_C_688 : begin
        fsm_output = 11'b10010110101;
        state_var_NS = COMP_LOOP_C_689;
      end
      COMP_LOOP_C_689 : begin
        fsm_output = 11'b10010110110;
        state_var_NS = COMP_LOOP_C_690;
      end
      COMP_LOOP_C_690 : begin
        fsm_output = 11'b10010110111;
        state_var_NS = COMP_LOOP_C_691;
      end
      COMP_LOOP_C_691 : begin
        fsm_output = 11'b10010111000;
        state_var_NS = COMP_LOOP_C_692;
      end
      COMP_LOOP_C_692 : begin
        fsm_output = 11'b10010111001;
        state_var_NS = COMP_LOOP_C_693;
      end
      COMP_LOOP_C_693 : begin
        fsm_output = 11'b10010111010;
        state_var_NS = COMP_LOOP_C_694;
      end
      COMP_LOOP_C_694 : begin
        fsm_output = 11'b10010111011;
        state_var_NS = COMP_LOOP_C_695;
      end
      COMP_LOOP_C_695 : begin
        fsm_output = 11'b10010111100;
        state_var_NS = COMP_LOOP_C_696;
      end
      COMP_LOOP_C_696 : begin
        fsm_output = 11'b10010111101;
        state_var_NS = COMP_LOOP_C_697;
      end
      COMP_LOOP_C_697 : begin
        fsm_output = 11'b10010111110;
        state_var_NS = COMP_LOOP_C_698;
      end
      COMP_LOOP_C_698 : begin
        fsm_output = 11'b10010111111;
        state_var_NS = COMP_LOOP_C_699;
      end
      COMP_LOOP_C_699 : begin
        fsm_output = 11'b10011000000;
        state_var_NS = COMP_LOOP_C_700;
      end
      COMP_LOOP_C_700 : begin
        fsm_output = 11'b10011000001;
        state_var_NS = COMP_LOOP_C_701;
      end
      COMP_LOOP_C_701 : begin
        fsm_output = 11'b10011000010;
        state_var_NS = COMP_LOOP_C_702;
      end
      COMP_LOOP_C_702 : begin
        fsm_output = 11'b10011000011;
        state_var_NS = COMP_LOOP_C_703;
      end
      COMP_LOOP_C_703 : begin
        fsm_output = 11'b10011000100;
        state_var_NS = COMP_LOOP_C_704;
      end
      COMP_LOOP_C_704 : begin
        fsm_output = 11'b10011000101;
        state_var_NS = COMP_LOOP_C_705;
      end
      COMP_LOOP_C_705 : begin
        fsm_output = 11'b10011000110;
        state_var_NS = COMP_LOOP_C_706;
      end
      COMP_LOOP_C_706 : begin
        fsm_output = 11'b10011000111;
        state_var_NS = COMP_LOOP_C_707;
      end
      COMP_LOOP_C_707 : begin
        fsm_output = 11'b10011001000;
        state_var_NS = COMP_LOOP_C_708;
      end
      COMP_LOOP_C_708 : begin
        fsm_output = 11'b10011001001;
        state_var_NS = COMP_LOOP_C_709;
      end
      COMP_LOOP_C_709 : begin
        fsm_output = 11'b10011001010;
        state_var_NS = COMP_LOOP_C_710;
      end
      COMP_LOOP_C_710 : begin
        fsm_output = 11'b10011001011;
        state_var_NS = COMP_LOOP_C_711;
      end
      COMP_LOOP_C_711 : begin
        fsm_output = 11'b10011001100;
        state_var_NS = COMP_LOOP_C_712;
      end
      COMP_LOOP_C_712 : begin
        fsm_output = 11'b10011001101;
        state_var_NS = COMP_LOOP_C_713;
      end
      COMP_LOOP_C_713 : begin
        fsm_output = 11'b10011001110;
        state_var_NS = COMP_LOOP_C_714;
      end
      COMP_LOOP_C_714 : begin
        fsm_output = 11'b10011001111;
        state_var_NS = COMP_LOOP_C_715;
      end
      COMP_LOOP_C_715 : begin
        fsm_output = 11'b10011010000;
        state_var_NS = COMP_LOOP_C_716;
      end
      COMP_LOOP_C_716 : begin
        fsm_output = 11'b10011010001;
        state_var_NS = COMP_LOOP_C_717;
      end
      COMP_LOOP_C_717 : begin
        fsm_output = 11'b10011010010;
        state_var_NS = COMP_LOOP_C_718;
      end
      COMP_LOOP_C_718 : begin
        fsm_output = 11'b10011010011;
        state_var_NS = COMP_LOOP_C_719;
      end
      COMP_LOOP_C_719 : begin
        fsm_output = 11'b10011010100;
        state_var_NS = COMP_LOOP_C_720;
      end
      COMP_LOOP_C_720 : begin
        fsm_output = 11'b10011010101;
        state_var_NS = COMP_LOOP_C_721;
      end
      COMP_LOOP_C_721 : begin
        fsm_output = 11'b10011010110;
        state_var_NS = COMP_LOOP_C_722;
      end
      COMP_LOOP_C_722 : begin
        fsm_output = 11'b10011010111;
        state_var_NS = COMP_LOOP_C_723;
      end
      COMP_LOOP_C_723 : begin
        fsm_output = 11'b10011011000;
        state_var_NS = COMP_LOOP_C_724;
      end
      COMP_LOOP_C_724 : begin
        fsm_output = 11'b10011011001;
        state_var_NS = COMP_LOOP_C_725;
      end
      COMP_LOOP_C_725 : begin
        fsm_output = 11'b10011011010;
        state_var_NS = COMP_LOOP_C_726;
      end
      COMP_LOOP_C_726 : begin
        fsm_output = 11'b10011011011;
        state_var_NS = COMP_LOOP_C_727;
      end
      COMP_LOOP_C_727 : begin
        fsm_output = 11'b10011011100;
        state_var_NS = COMP_LOOP_C_728;
      end
      COMP_LOOP_C_728 : begin
        fsm_output = 11'b10011011101;
        state_var_NS = COMP_LOOP_C_729;
      end
      COMP_LOOP_C_729 : begin
        fsm_output = 11'b10011011110;
        state_var_NS = COMP_LOOP_C_730;
      end
      COMP_LOOP_C_730 : begin
        fsm_output = 11'b10011011111;
        state_var_NS = COMP_LOOP_C_731;
      end
      COMP_LOOP_C_731 : begin
        fsm_output = 11'b10011100000;
        state_var_NS = COMP_LOOP_C_732;
      end
      COMP_LOOP_C_732 : begin
        fsm_output = 11'b10011100001;
        state_var_NS = COMP_LOOP_C_733;
      end
      COMP_LOOP_C_733 : begin
        fsm_output = 11'b10011100010;
        state_var_NS = COMP_LOOP_C_734;
      end
      COMP_LOOP_C_734 : begin
        fsm_output = 11'b10011100011;
        state_var_NS = COMP_LOOP_C_735;
      end
      COMP_LOOP_C_735 : begin
        fsm_output = 11'b10011100100;
        state_var_NS = COMP_LOOP_C_736;
      end
      COMP_LOOP_C_736 : begin
        fsm_output = 11'b10011100101;
        state_var_NS = COMP_LOOP_C_737;
      end
      COMP_LOOP_C_737 : begin
        fsm_output = 11'b10011100110;
        state_var_NS = COMP_LOOP_C_738;
      end
      COMP_LOOP_C_738 : begin
        fsm_output = 11'b10011100111;
        state_var_NS = COMP_LOOP_C_739;
      end
      COMP_LOOP_C_739 : begin
        fsm_output = 11'b10011101000;
        state_var_NS = COMP_LOOP_C_740;
      end
      COMP_LOOP_C_740 : begin
        fsm_output = 11'b10011101001;
        state_var_NS = COMP_LOOP_C_741;
      end
      COMP_LOOP_C_741 : begin
        fsm_output = 11'b10011101010;
        state_var_NS = COMP_LOOP_C_742;
      end
      COMP_LOOP_C_742 : begin
        fsm_output = 11'b10011101011;
        state_var_NS = COMP_LOOP_C_743;
      end
      COMP_LOOP_C_743 : begin
        fsm_output = 11'b10011101100;
        state_var_NS = COMP_LOOP_C_744;
      end
      COMP_LOOP_C_744 : begin
        fsm_output = 11'b10011101101;
        if ( COMP_LOOP_C_744_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_745;
        end
      end
      COMP_LOOP_C_745 : begin
        fsm_output = 11'b10011101110;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_0;
      end
      COMP_LOOP_13_modExp_1_while_C_0 : begin
        fsm_output = 11'b10011101111;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_1;
      end
      COMP_LOOP_13_modExp_1_while_C_1 : begin
        fsm_output = 11'b10011110000;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_2;
      end
      COMP_LOOP_13_modExp_1_while_C_2 : begin
        fsm_output = 11'b10011110001;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_3;
      end
      COMP_LOOP_13_modExp_1_while_C_3 : begin
        fsm_output = 11'b10011110010;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_4;
      end
      COMP_LOOP_13_modExp_1_while_C_4 : begin
        fsm_output = 11'b10011110011;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_5;
      end
      COMP_LOOP_13_modExp_1_while_C_5 : begin
        fsm_output = 11'b10011110100;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_6;
      end
      COMP_LOOP_13_modExp_1_while_C_6 : begin
        fsm_output = 11'b10011110101;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_7;
      end
      COMP_LOOP_13_modExp_1_while_C_7 : begin
        fsm_output = 11'b10011110110;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_8;
      end
      COMP_LOOP_13_modExp_1_while_C_8 : begin
        fsm_output = 11'b10011110111;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_9;
      end
      COMP_LOOP_13_modExp_1_while_C_9 : begin
        fsm_output = 11'b10011111000;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_10;
      end
      COMP_LOOP_13_modExp_1_while_C_10 : begin
        fsm_output = 11'b10011111001;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_11;
      end
      COMP_LOOP_13_modExp_1_while_C_11 : begin
        fsm_output = 11'b10011111010;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_12;
      end
      COMP_LOOP_13_modExp_1_while_C_12 : begin
        fsm_output = 11'b10011111011;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_13;
      end
      COMP_LOOP_13_modExp_1_while_C_13 : begin
        fsm_output = 11'b10011111100;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_14;
      end
      COMP_LOOP_13_modExp_1_while_C_14 : begin
        fsm_output = 11'b10011111101;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_15;
      end
      COMP_LOOP_13_modExp_1_while_C_15 : begin
        fsm_output = 11'b10011111110;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_16;
      end
      COMP_LOOP_13_modExp_1_while_C_16 : begin
        fsm_output = 11'b10011111111;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_17;
      end
      COMP_LOOP_13_modExp_1_while_C_17 : begin
        fsm_output = 11'b10100000000;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_18;
      end
      COMP_LOOP_13_modExp_1_while_C_18 : begin
        fsm_output = 11'b10100000001;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_19;
      end
      COMP_LOOP_13_modExp_1_while_C_19 : begin
        fsm_output = 11'b10100000010;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_20;
      end
      COMP_LOOP_13_modExp_1_while_C_20 : begin
        fsm_output = 11'b10100000011;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_21;
      end
      COMP_LOOP_13_modExp_1_while_C_21 : begin
        fsm_output = 11'b10100000100;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_22;
      end
      COMP_LOOP_13_modExp_1_while_C_22 : begin
        fsm_output = 11'b10100000101;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_23;
      end
      COMP_LOOP_13_modExp_1_while_C_23 : begin
        fsm_output = 11'b10100000110;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_24;
      end
      COMP_LOOP_13_modExp_1_while_C_24 : begin
        fsm_output = 11'b10100000111;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_25;
      end
      COMP_LOOP_13_modExp_1_while_C_25 : begin
        fsm_output = 11'b10100001000;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_26;
      end
      COMP_LOOP_13_modExp_1_while_C_26 : begin
        fsm_output = 11'b10100001001;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_27;
      end
      COMP_LOOP_13_modExp_1_while_C_27 : begin
        fsm_output = 11'b10100001010;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_28;
      end
      COMP_LOOP_13_modExp_1_while_C_28 : begin
        fsm_output = 11'b10100001011;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_29;
      end
      COMP_LOOP_13_modExp_1_while_C_29 : begin
        fsm_output = 11'b10100001100;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_30;
      end
      COMP_LOOP_13_modExp_1_while_C_30 : begin
        fsm_output = 11'b10100001101;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_31;
      end
      COMP_LOOP_13_modExp_1_while_C_31 : begin
        fsm_output = 11'b10100001110;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_32;
      end
      COMP_LOOP_13_modExp_1_while_C_32 : begin
        fsm_output = 11'b10100001111;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_33;
      end
      COMP_LOOP_13_modExp_1_while_C_33 : begin
        fsm_output = 11'b10100010000;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_34;
      end
      COMP_LOOP_13_modExp_1_while_C_34 : begin
        fsm_output = 11'b10100010001;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_35;
      end
      COMP_LOOP_13_modExp_1_while_C_35 : begin
        fsm_output = 11'b10100010010;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_36;
      end
      COMP_LOOP_13_modExp_1_while_C_36 : begin
        fsm_output = 11'b10100010011;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_37;
      end
      COMP_LOOP_13_modExp_1_while_C_37 : begin
        fsm_output = 11'b10100010100;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_38;
      end
      COMP_LOOP_13_modExp_1_while_C_38 : begin
        fsm_output = 11'b10100010101;
        if ( COMP_LOOP_13_modExp_1_while_C_38_tr0 ) begin
          state_var_NS = COMP_LOOP_C_746;
        end
        else begin
          state_var_NS = COMP_LOOP_13_modExp_1_while_C_0;
        end
      end
      COMP_LOOP_C_746 : begin
        fsm_output = 11'b10100010110;
        state_var_NS = COMP_LOOP_C_747;
      end
      COMP_LOOP_C_747 : begin
        fsm_output = 11'b10100010111;
        state_var_NS = COMP_LOOP_C_748;
      end
      COMP_LOOP_C_748 : begin
        fsm_output = 11'b10100011000;
        state_var_NS = COMP_LOOP_C_749;
      end
      COMP_LOOP_C_749 : begin
        fsm_output = 11'b10100011001;
        state_var_NS = COMP_LOOP_C_750;
      end
      COMP_LOOP_C_750 : begin
        fsm_output = 11'b10100011010;
        state_var_NS = COMP_LOOP_C_751;
      end
      COMP_LOOP_C_751 : begin
        fsm_output = 11'b10100011011;
        state_var_NS = COMP_LOOP_C_752;
      end
      COMP_LOOP_C_752 : begin
        fsm_output = 11'b10100011100;
        state_var_NS = COMP_LOOP_C_753;
      end
      COMP_LOOP_C_753 : begin
        fsm_output = 11'b10100011101;
        state_var_NS = COMP_LOOP_C_754;
      end
      COMP_LOOP_C_754 : begin
        fsm_output = 11'b10100011110;
        state_var_NS = COMP_LOOP_C_755;
      end
      COMP_LOOP_C_755 : begin
        fsm_output = 11'b10100011111;
        state_var_NS = COMP_LOOP_C_756;
      end
      COMP_LOOP_C_756 : begin
        fsm_output = 11'b10100100000;
        state_var_NS = COMP_LOOP_C_757;
      end
      COMP_LOOP_C_757 : begin
        fsm_output = 11'b10100100001;
        state_var_NS = COMP_LOOP_C_758;
      end
      COMP_LOOP_C_758 : begin
        fsm_output = 11'b10100100010;
        state_var_NS = COMP_LOOP_C_759;
      end
      COMP_LOOP_C_759 : begin
        fsm_output = 11'b10100100011;
        state_var_NS = COMP_LOOP_C_760;
      end
      COMP_LOOP_C_760 : begin
        fsm_output = 11'b10100100100;
        state_var_NS = COMP_LOOP_C_761;
      end
      COMP_LOOP_C_761 : begin
        fsm_output = 11'b10100100101;
        state_var_NS = COMP_LOOP_C_762;
      end
      COMP_LOOP_C_762 : begin
        fsm_output = 11'b10100100110;
        state_var_NS = COMP_LOOP_C_763;
      end
      COMP_LOOP_C_763 : begin
        fsm_output = 11'b10100100111;
        state_var_NS = COMP_LOOP_C_764;
      end
      COMP_LOOP_C_764 : begin
        fsm_output = 11'b10100101000;
        state_var_NS = COMP_LOOP_C_765;
      end
      COMP_LOOP_C_765 : begin
        fsm_output = 11'b10100101001;
        state_var_NS = COMP_LOOP_C_766;
      end
      COMP_LOOP_C_766 : begin
        fsm_output = 11'b10100101010;
        state_var_NS = COMP_LOOP_C_767;
      end
      COMP_LOOP_C_767 : begin
        fsm_output = 11'b10100101011;
        state_var_NS = COMP_LOOP_C_768;
      end
      COMP_LOOP_C_768 : begin
        fsm_output = 11'b10100101100;
        state_var_NS = COMP_LOOP_C_769;
      end
      COMP_LOOP_C_769 : begin
        fsm_output = 11'b10100101101;
        state_var_NS = COMP_LOOP_C_770;
      end
      COMP_LOOP_C_770 : begin
        fsm_output = 11'b10100101110;
        state_var_NS = COMP_LOOP_C_771;
      end
      COMP_LOOP_C_771 : begin
        fsm_output = 11'b10100101111;
        state_var_NS = COMP_LOOP_C_772;
      end
      COMP_LOOP_C_772 : begin
        fsm_output = 11'b10100110000;
        state_var_NS = COMP_LOOP_C_773;
      end
      COMP_LOOP_C_773 : begin
        fsm_output = 11'b10100110001;
        state_var_NS = COMP_LOOP_C_774;
      end
      COMP_LOOP_C_774 : begin
        fsm_output = 11'b10100110010;
        state_var_NS = COMP_LOOP_C_775;
      end
      COMP_LOOP_C_775 : begin
        fsm_output = 11'b10100110011;
        state_var_NS = COMP_LOOP_C_776;
      end
      COMP_LOOP_C_776 : begin
        fsm_output = 11'b10100110100;
        state_var_NS = COMP_LOOP_C_777;
      end
      COMP_LOOP_C_777 : begin
        fsm_output = 11'b10100110101;
        state_var_NS = COMP_LOOP_C_778;
      end
      COMP_LOOP_C_778 : begin
        fsm_output = 11'b10100110110;
        state_var_NS = COMP_LOOP_C_779;
      end
      COMP_LOOP_C_779 : begin
        fsm_output = 11'b10100110111;
        state_var_NS = COMP_LOOP_C_780;
      end
      COMP_LOOP_C_780 : begin
        fsm_output = 11'b10100111000;
        state_var_NS = COMP_LOOP_C_781;
      end
      COMP_LOOP_C_781 : begin
        fsm_output = 11'b10100111001;
        state_var_NS = COMP_LOOP_C_782;
      end
      COMP_LOOP_C_782 : begin
        fsm_output = 11'b10100111010;
        state_var_NS = COMP_LOOP_C_783;
      end
      COMP_LOOP_C_783 : begin
        fsm_output = 11'b10100111011;
        state_var_NS = COMP_LOOP_C_784;
      end
      COMP_LOOP_C_784 : begin
        fsm_output = 11'b10100111100;
        state_var_NS = COMP_LOOP_C_785;
      end
      COMP_LOOP_C_785 : begin
        fsm_output = 11'b10100111101;
        state_var_NS = COMP_LOOP_C_786;
      end
      COMP_LOOP_C_786 : begin
        fsm_output = 11'b10100111110;
        state_var_NS = COMP_LOOP_C_787;
      end
      COMP_LOOP_C_787 : begin
        fsm_output = 11'b10100111111;
        state_var_NS = COMP_LOOP_C_788;
      end
      COMP_LOOP_C_788 : begin
        fsm_output = 11'b10101000000;
        state_var_NS = COMP_LOOP_C_789;
      end
      COMP_LOOP_C_789 : begin
        fsm_output = 11'b10101000001;
        state_var_NS = COMP_LOOP_C_790;
      end
      COMP_LOOP_C_790 : begin
        fsm_output = 11'b10101000010;
        state_var_NS = COMP_LOOP_C_791;
      end
      COMP_LOOP_C_791 : begin
        fsm_output = 11'b10101000011;
        state_var_NS = COMP_LOOP_C_792;
      end
      COMP_LOOP_C_792 : begin
        fsm_output = 11'b10101000100;
        state_var_NS = COMP_LOOP_C_793;
      end
      COMP_LOOP_C_793 : begin
        fsm_output = 11'b10101000101;
        state_var_NS = COMP_LOOP_C_794;
      end
      COMP_LOOP_C_794 : begin
        fsm_output = 11'b10101000110;
        state_var_NS = COMP_LOOP_C_795;
      end
      COMP_LOOP_C_795 : begin
        fsm_output = 11'b10101000111;
        state_var_NS = COMP_LOOP_C_796;
      end
      COMP_LOOP_C_796 : begin
        fsm_output = 11'b10101001000;
        state_var_NS = COMP_LOOP_C_797;
      end
      COMP_LOOP_C_797 : begin
        fsm_output = 11'b10101001001;
        state_var_NS = COMP_LOOP_C_798;
      end
      COMP_LOOP_C_798 : begin
        fsm_output = 11'b10101001010;
        state_var_NS = COMP_LOOP_C_799;
      end
      COMP_LOOP_C_799 : begin
        fsm_output = 11'b10101001011;
        state_var_NS = COMP_LOOP_C_800;
      end
      COMP_LOOP_C_800 : begin
        fsm_output = 11'b10101001100;
        state_var_NS = COMP_LOOP_C_801;
      end
      COMP_LOOP_C_801 : begin
        fsm_output = 11'b10101001101;
        state_var_NS = COMP_LOOP_C_802;
      end
      COMP_LOOP_C_802 : begin
        fsm_output = 11'b10101001110;
        state_var_NS = COMP_LOOP_C_803;
      end
      COMP_LOOP_C_803 : begin
        fsm_output = 11'b10101001111;
        state_var_NS = COMP_LOOP_C_804;
      end
      COMP_LOOP_C_804 : begin
        fsm_output = 11'b10101010000;
        state_var_NS = COMP_LOOP_C_805;
      end
      COMP_LOOP_C_805 : begin
        fsm_output = 11'b10101010001;
        state_var_NS = COMP_LOOP_C_806;
      end
      COMP_LOOP_C_806 : begin
        fsm_output = 11'b10101010010;
        if ( COMP_LOOP_C_806_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_807;
        end
      end
      COMP_LOOP_C_807 : begin
        fsm_output = 11'b10101010011;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_0;
      end
      COMP_LOOP_14_modExp_1_while_C_0 : begin
        fsm_output = 11'b10101010100;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_1;
      end
      COMP_LOOP_14_modExp_1_while_C_1 : begin
        fsm_output = 11'b10101010101;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_2;
      end
      COMP_LOOP_14_modExp_1_while_C_2 : begin
        fsm_output = 11'b10101010110;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_3;
      end
      COMP_LOOP_14_modExp_1_while_C_3 : begin
        fsm_output = 11'b10101010111;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_4;
      end
      COMP_LOOP_14_modExp_1_while_C_4 : begin
        fsm_output = 11'b10101011000;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_5;
      end
      COMP_LOOP_14_modExp_1_while_C_5 : begin
        fsm_output = 11'b10101011001;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_6;
      end
      COMP_LOOP_14_modExp_1_while_C_6 : begin
        fsm_output = 11'b10101011010;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_7;
      end
      COMP_LOOP_14_modExp_1_while_C_7 : begin
        fsm_output = 11'b10101011011;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_8;
      end
      COMP_LOOP_14_modExp_1_while_C_8 : begin
        fsm_output = 11'b10101011100;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_9;
      end
      COMP_LOOP_14_modExp_1_while_C_9 : begin
        fsm_output = 11'b10101011101;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_10;
      end
      COMP_LOOP_14_modExp_1_while_C_10 : begin
        fsm_output = 11'b10101011110;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_11;
      end
      COMP_LOOP_14_modExp_1_while_C_11 : begin
        fsm_output = 11'b10101011111;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_12;
      end
      COMP_LOOP_14_modExp_1_while_C_12 : begin
        fsm_output = 11'b10101100000;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_13;
      end
      COMP_LOOP_14_modExp_1_while_C_13 : begin
        fsm_output = 11'b10101100001;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_14;
      end
      COMP_LOOP_14_modExp_1_while_C_14 : begin
        fsm_output = 11'b10101100010;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_15;
      end
      COMP_LOOP_14_modExp_1_while_C_15 : begin
        fsm_output = 11'b10101100011;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_16;
      end
      COMP_LOOP_14_modExp_1_while_C_16 : begin
        fsm_output = 11'b10101100100;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_17;
      end
      COMP_LOOP_14_modExp_1_while_C_17 : begin
        fsm_output = 11'b10101100101;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_18;
      end
      COMP_LOOP_14_modExp_1_while_C_18 : begin
        fsm_output = 11'b10101100110;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_19;
      end
      COMP_LOOP_14_modExp_1_while_C_19 : begin
        fsm_output = 11'b10101100111;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_20;
      end
      COMP_LOOP_14_modExp_1_while_C_20 : begin
        fsm_output = 11'b10101101000;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_21;
      end
      COMP_LOOP_14_modExp_1_while_C_21 : begin
        fsm_output = 11'b10101101001;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_22;
      end
      COMP_LOOP_14_modExp_1_while_C_22 : begin
        fsm_output = 11'b10101101010;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_23;
      end
      COMP_LOOP_14_modExp_1_while_C_23 : begin
        fsm_output = 11'b10101101011;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_24;
      end
      COMP_LOOP_14_modExp_1_while_C_24 : begin
        fsm_output = 11'b10101101100;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_25;
      end
      COMP_LOOP_14_modExp_1_while_C_25 : begin
        fsm_output = 11'b10101101101;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_26;
      end
      COMP_LOOP_14_modExp_1_while_C_26 : begin
        fsm_output = 11'b10101101110;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_27;
      end
      COMP_LOOP_14_modExp_1_while_C_27 : begin
        fsm_output = 11'b10101101111;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_28;
      end
      COMP_LOOP_14_modExp_1_while_C_28 : begin
        fsm_output = 11'b10101110000;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_29;
      end
      COMP_LOOP_14_modExp_1_while_C_29 : begin
        fsm_output = 11'b10101110001;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_30;
      end
      COMP_LOOP_14_modExp_1_while_C_30 : begin
        fsm_output = 11'b10101110010;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_31;
      end
      COMP_LOOP_14_modExp_1_while_C_31 : begin
        fsm_output = 11'b10101110011;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_32;
      end
      COMP_LOOP_14_modExp_1_while_C_32 : begin
        fsm_output = 11'b10101110100;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_33;
      end
      COMP_LOOP_14_modExp_1_while_C_33 : begin
        fsm_output = 11'b10101110101;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_34;
      end
      COMP_LOOP_14_modExp_1_while_C_34 : begin
        fsm_output = 11'b10101110110;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_35;
      end
      COMP_LOOP_14_modExp_1_while_C_35 : begin
        fsm_output = 11'b10101110111;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_36;
      end
      COMP_LOOP_14_modExp_1_while_C_36 : begin
        fsm_output = 11'b10101111000;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_37;
      end
      COMP_LOOP_14_modExp_1_while_C_37 : begin
        fsm_output = 11'b10101111001;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_38;
      end
      COMP_LOOP_14_modExp_1_while_C_38 : begin
        fsm_output = 11'b10101111010;
        if ( COMP_LOOP_14_modExp_1_while_C_38_tr0 ) begin
          state_var_NS = COMP_LOOP_C_808;
        end
        else begin
          state_var_NS = COMP_LOOP_14_modExp_1_while_C_0;
        end
      end
      COMP_LOOP_C_808 : begin
        fsm_output = 11'b10101111011;
        state_var_NS = COMP_LOOP_C_809;
      end
      COMP_LOOP_C_809 : begin
        fsm_output = 11'b10101111100;
        state_var_NS = COMP_LOOP_C_810;
      end
      COMP_LOOP_C_810 : begin
        fsm_output = 11'b10101111101;
        state_var_NS = COMP_LOOP_C_811;
      end
      COMP_LOOP_C_811 : begin
        fsm_output = 11'b10101111110;
        state_var_NS = COMP_LOOP_C_812;
      end
      COMP_LOOP_C_812 : begin
        fsm_output = 11'b10101111111;
        state_var_NS = COMP_LOOP_C_813;
      end
      COMP_LOOP_C_813 : begin
        fsm_output = 11'b10110000000;
        state_var_NS = COMP_LOOP_C_814;
      end
      COMP_LOOP_C_814 : begin
        fsm_output = 11'b10110000001;
        state_var_NS = COMP_LOOP_C_815;
      end
      COMP_LOOP_C_815 : begin
        fsm_output = 11'b10110000010;
        state_var_NS = COMP_LOOP_C_816;
      end
      COMP_LOOP_C_816 : begin
        fsm_output = 11'b10110000011;
        state_var_NS = COMP_LOOP_C_817;
      end
      COMP_LOOP_C_817 : begin
        fsm_output = 11'b10110000100;
        state_var_NS = COMP_LOOP_C_818;
      end
      COMP_LOOP_C_818 : begin
        fsm_output = 11'b10110000101;
        state_var_NS = COMP_LOOP_C_819;
      end
      COMP_LOOP_C_819 : begin
        fsm_output = 11'b10110000110;
        state_var_NS = COMP_LOOP_C_820;
      end
      COMP_LOOP_C_820 : begin
        fsm_output = 11'b10110000111;
        state_var_NS = COMP_LOOP_C_821;
      end
      COMP_LOOP_C_821 : begin
        fsm_output = 11'b10110001000;
        state_var_NS = COMP_LOOP_C_822;
      end
      COMP_LOOP_C_822 : begin
        fsm_output = 11'b10110001001;
        state_var_NS = COMP_LOOP_C_823;
      end
      COMP_LOOP_C_823 : begin
        fsm_output = 11'b10110001010;
        state_var_NS = COMP_LOOP_C_824;
      end
      COMP_LOOP_C_824 : begin
        fsm_output = 11'b10110001011;
        state_var_NS = COMP_LOOP_C_825;
      end
      COMP_LOOP_C_825 : begin
        fsm_output = 11'b10110001100;
        state_var_NS = COMP_LOOP_C_826;
      end
      COMP_LOOP_C_826 : begin
        fsm_output = 11'b10110001101;
        state_var_NS = COMP_LOOP_C_827;
      end
      COMP_LOOP_C_827 : begin
        fsm_output = 11'b10110001110;
        state_var_NS = COMP_LOOP_C_828;
      end
      COMP_LOOP_C_828 : begin
        fsm_output = 11'b10110001111;
        state_var_NS = COMP_LOOP_C_829;
      end
      COMP_LOOP_C_829 : begin
        fsm_output = 11'b10110010000;
        state_var_NS = COMP_LOOP_C_830;
      end
      COMP_LOOP_C_830 : begin
        fsm_output = 11'b10110010001;
        state_var_NS = COMP_LOOP_C_831;
      end
      COMP_LOOP_C_831 : begin
        fsm_output = 11'b10110010010;
        state_var_NS = COMP_LOOP_C_832;
      end
      COMP_LOOP_C_832 : begin
        fsm_output = 11'b10110010011;
        state_var_NS = COMP_LOOP_C_833;
      end
      COMP_LOOP_C_833 : begin
        fsm_output = 11'b10110010100;
        state_var_NS = COMP_LOOP_C_834;
      end
      COMP_LOOP_C_834 : begin
        fsm_output = 11'b10110010101;
        state_var_NS = COMP_LOOP_C_835;
      end
      COMP_LOOP_C_835 : begin
        fsm_output = 11'b10110010110;
        state_var_NS = COMP_LOOP_C_836;
      end
      COMP_LOOP_C_836 : begin
        fsm_output = 11'b10110010111;
        state_var_NS = COMP_LOOP_C_837;
      end
      COMP_LOOP_C_837 : begin
        fsm_output = 11'b10110011000;
        state_var_NS = COMP_LOOP_C_838;
      end
      COMP_LOOP_C_838 : begin
        fsm_output = 11'b10110011001;
        state_var_NS = COMP_LOOP_C_839;
      end
      COMP_LOOP_C_839 : begin
        fsm_output = 11'b10110011010;
        state_var_NS = COMP_LOOP_C_840;
      end
      COMP_LOOP_C_840 : begin
        fsm_output = 11'b10110011011;
        state_var_NS = COMP_LOOP_C_841;
      end
      COMP_LOOP_C_841 : begin
        fsm_output = 11'b10110011100;
        state_var_NS = COMP_LOOP_C_842;
      end
      COMP_LOOP_C_842 : begin
        fsm_output = 11'b10110011101;
        state_var_NS = COMP_LOOP_C_843;
      end
      COMP_LOOP_C_843 : begin
        fsm_output = 11'b10110011110;
        state_var_NS = COMP_LOOP_C_844;
      end
      COMP_LOOP_C_844 : begin
        fsm_output = 11'b10110011111;
        state_var_NS = COMP_LOOP_C_845;
      end
      COMP_LOOP_C_845 : begin
        fsm_output = 11'b10110100000;
        state_var_NS = COMP_LOOP_C_846;
      end
      COMP_LOOP_C_846 : begin
        fsm_output = 11'b10110100001;
        state_var_NS = COMP_LOOP_C_847;
      end
      COMP_LOOP_C_847 : begin
        fsm_output = 11'b10110100010;
        state_var_NS = COMP_LOOP_C_848;
      end
      COMP_LOOP_C_848 : begin
        fsm_output = 11'b10110100011;
        state_var_NS = COMP_LOOP_C_849;
      end
      COMP_LOOP_C_849 : begin
        fsm_output = 11'b10110100100;
        state_var_NS = COMP_LOOP_C_850;
      end
      COMP_LOOP_C_850 : begin
        fsm_output = 11'b10110100101;
        state_var_NS = COMP_LOOP_C_851;
      end
      COMP_LOOP_C_851 : begin
        fsm_output = 11'b10110100110;
        state_var_NS = COMP_LOOP_C_852;
      end
      COMP_LOOP_C_852 : begin
        fsm_output = 11'b10110100111;
        state_var_NS = COMP_LOOP_C_853;
      end
      COMP_LOOP_C_853 : begin
        fsm_output = 11'b10110101000;
        state_var_NS = COMP_LOOP_C_854;
      end
      COMP_LOOP_C_854 : begin
        fsm_output = 11'b10110101001;
        state_var_NS = COMP_LOOP_C_855;
      end
      COMP_LOOP_C_855 : begin
        fsm_output = 11'b10110101010;
        state_var_NS = COMP_LOOP_C_856;
      end
      COMP_LOOP_C_856 : begin
        fsm_output = 11'b10110101011;
        state_var_NS = COMP_LOOP_C_857;
      end
      COMP_LOOP_C_857 : begin
        fsm_output = 11'b10110101100;
        state_var_NS = COMP_LOOP_C_858;
      end
      COMP_LOOP_C_858 : begin
        fsm_output = 11'b10110101101;
        state_var_NS = COMP_LOOP_C_859;
      end
      COMP_LOOP_C_859 : begin
        fsm_output = 11'b10110101110;
        state_var_NS = COMP_LOOP_C_860;
      end
      COMP_LOOP_C_860 : begin
        fsm_output = 11'b10110101111;
        state_var_NS = COMP_LOOP_C_861;
      end
      COMP_LOOP_C_861 : begin
        fsm_output = 11'b10110110000;
        state_var_NS = COMP_LOOP_C_862;
      end
      COMP_LOOP_C_862 : begin
        fsm_output = 11'b10110110001;
        state_var_NS = COMP_LOOP_C_863;
      end
      COMP_LOOP_C_863 : begin
        fsm_output = 11'b10110110010;
        state_var_NS = COMP_LOOP_C_864;
      end
      COMP_LOOP_C_864 : begin
        fsm_output = 11'b10110110011;
        state_var_NS = COMP_LOOP_C_865;
      end
      COMP_LOOP_C_865 : begin
        fsm_output = 11'b10110110100;
        state_var_NS = COMP_LOOP_C_866;
      end
      COMP_LOOP_C_866 : begin
        fsm_output = 11'b10110110101;
        state_var_NS = COMP_LOOP_C_867;
      end
      COMP_LOOP_C_867 : begin
        fsm_output = 11'b10110110110;
        state_var_NS = COMP_LOOP_C_868;
      end
      COMP_LOOP_C_868 : begin
        fsm_output = 11'b10110110111;
        if ( COMP_LOOP_C_868_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_869;
        end
      end
      COMP_LOOP_C_869 : begin
        fsm_output = 11'b10110111000;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_0;
      end
      COMP_LOOP_15_modExp_1_while_C_0 : begin
        fsm_output = 11'b10110111001;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_1;
      end
      COMP_LOOP_15_modExp_1_while_C_1 : begin
        fsm_output = 11'b10110111010;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_2;
      end
      COMP_LOOP_15_modExp_1_while_C_2 : begin
        fsm_output = 11'b10110111011;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_3;
      end
      COMP_LOOP_15_modExp_1_while_C_3 : begin
        fsm_output = 11'b10110111100;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_4;
      end
      COMP_LOOP_15_modExp_1_while_C_4 : begin
        fsm_output = 11'b10110111101;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_5;
      end
      COMP_LOOP_15_modExp_1_while_C_5 : begin
        fsm_output = 11'b10110111110;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_6;
      end
      COMP_LOOP_15_modExp_1_while_C_6 : begin
        fsm_output = 11'b10110111111;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_7;
      end
      COMP_LOOP_15_modExp_1_while_C_7 : begin
        fsm_output = 11'b10111000000;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_8;
      end
      COMP_LOOP_15_modExp_1_while_C_8 : begin
        fsm_output = 11'b10111000001;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_9;
      end
      COMP_LOOP_15_modExp_1_while_C_9 : begin
        fsm_output = 11'b10111000010;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_10;
      end
      COMP_LOOP_15_modExp_1_while_C_10 : begin
        fsm_output = 11'b10111000011;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_11;
      end
      COMP_LOOP_15_modExp_1_while_C_11 : begin
        fsm_output = 11'b10111000100;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_12;
      end
      COMP_LOOP_15_modExp_1_while_C_12 : begin
        fsm_output = 11'b10111000101;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_13;
      end
      COMP_LOOP_15_modExp_1_while_C_13 : begin
        fsm_output = 11'b10111000110;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_14;
      end
      COMP_LOOP_15_modExp_1_while_C_14 : begin
        fsm_output = 11'b10111000111;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_15;
      end
      COMP_LOOP_15_modExp_1_while_C_15 : begin
        fsm_output = 11'b10111001000;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_16;
      end
      COMP_LOOP_15_modExp_1_while_C_16 : begin
        fsm_output = 11'b10111001001;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_17;
      end
      COMP_LOOP_15_modExp_1_while_C_17 : begin
        fsm_output = 11'b10111001010;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_18;
      end
      COMP_LOOP_15_modExp_1_while_C_18 : begin
        fsm_output = 11'b10111001011;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_19;
      end
      COMP_LOOP_15_modExp_1_while_C_19 : begin
        fsm_output = 11'b10111001100;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_20;
      end
      COMP_LOOP_15_modExp_1_while_C_20 : begin
        fsm_output = 11'b10111001101;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_21;
      end
      COMP_LOOP_15_modExp_1_while_C_21 : begin
        fsm_output = 11'b10111001110;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_22;
      end
      COMP_LOOP_15_modExp_1_while_C_22 : begin
        fsm_output = 11'b10111001111;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_23;
      end
      COMP_LOOP_15_modExp_1_while_C_23 : begin
        fsm_output = 11'b10111010000;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_24;
      end
      COMP_LOOP_15_modExp_1_while_C_24 : begin
        fsm_output = 11'b10111010001;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_25;
      end
      COMP_LOOP_15_modExp_1_while_C_25 : begin
        fsm_output = 11'b10111010010;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_26;
      end
      COMP_LOOP_15_modExp_1_while_C_26 : begin
        fsm_output = 11'b10111010011;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_27;
      end
      COMP_LOOP_15_modExp_1_while_C_27 : begin
        fsm_output = 11'b10111010100;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_28;
      end
      COMP_LOOP_15_modExp_1_while_C_28 : begin
        fsm_output = 11'b10111010101;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_29;
      end
      COMP_LOOP_15_modExp_1_while_C_29 : begin
        fsm_output = 11'b10111010110;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_30;
      end
      COMP_LOOP_15_modExp_1_while_C_30 : begin
        fsm_output = 11'b10111010111;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_31;
      end
      COMP_LOOP_15_modExp_1_while_C_31 : begin
        fsm_output = 11'b10111011000;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_32;
      end
      COMP_LOOP_15_modExp_1_while_C_32 : begin
        fsm_output = 11'b10111011001;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_33;
      end
      COMP_LOOP_15_modExp_1_while_C_33 : begin
        fsm_output = 11'b10111011010;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_34;
      end
      COMP_LOOP_15_modExp_1_while_C_34 : begin
        fsm_output = 11'b10111011011;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_35;
      end
      COMP_LOOP_15_modExp_1_while_C_35 : begin
        fsm_output = 11'b10111011100;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_36;
      end
      COMP_LOOP_15_modExp_1_while_C_36 : begin
        fsm_output = 11'b10111011101;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_37;
      end
      COMP_LOOP_15_modExp_1_while_C_37 : begin
        fsm_output = 11'b10111011110;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_38;
      end
      COMP_LOOP_15_modExp_1_while_C_38 : begin
        fsm_output = 11'b10111011111;
        if ( COMP_LOOP_15_modExp_1_while_C_38_tr0 ) begin
          state_var_NS = COMP_LOOP_C_870;
        end
        else begin
          state_var_NS = COMP_LOOP_15_modExp_1_while_C_0;
        end
      end
      COMP_LOOP_C_870 : begin
        fsm_output = 11'b10111100000;
        state_var_NS = COMP_LOOP_C_871;
      end
      COMP_LOOP_C_871 : begin
        fsm_output = 11'b10111100001;
        state_var_NS = COMP_LOOP_C_872;
      end
      COMP_LOOP_C_872 : begin
        fsm_output = 11'b10111100010;
        state_var_NS = COMP_LOOP_C_873;
      end
      COMP_LOOP_C_873 : begin
        fsm_output = 11'b10111100011;
        state_var_NS = COMP_LOOP_C_874;
      end
      COMP_LOOP_C_874 : begin
        fsm_output = 11'b10111100100;
        state_var_NS = COMP_LOOP_C_875;
      end
      COMP_LOOP_C_875 : begin
        fsm_output = 11'b10111100101;
        state_var_NS = COMP_LOOP_C_876;
      end
      COMP_LOOP_C_876 : begin
        fsm_output = 11'b10111100110;
        state_var_NS = COMP_LOOP_C_877;
      end
      COMP_LOOP_C_877 : begin
        fsm_output = 11'b10111100111;
        state_var_NS = COMP_LOOP_C_878;
      end
      COMP_LOOP_C_878 : begin
        fsm_output = 11'b10111101000;
        state_var_NS = COMP_LOOP_C_879;
      end
      COMP_LOOP_C_879 : begin
        fsm_output = 11'b10111101001;
        state_var_NS = COMP_LOOP_C_880;
      end
      COMP_LOOP_C_880 : begin
        fsm_output = 11'b10111101010;
        state_var_NS = COMP_LOOP_C_881;
      end
      COMP_LOOP_C_881 : begin
        fsm_output = 11'b10111101011;
        state_var_NS = COMP_LOOP_C_882;
      end
      COMP_LOOP_C_882 : begin
        fsm_output = 11'b10111101100;
        state_var_NS = COMP_LOOP_C_883;
      end
      COMP_LOOP_C_883 : begin
        fsm_output = 11'b10111101101;
        state_var_NS = COMP_LOOP_C_884;
      end
      COMP_LOOP_C_884 : begin
        fsm_output = 11'b10111101110;
        state_var_NS = COMP_LOOP_C_885;
      end
      COMP_LOOP_C_885 : begin
        fsm_output = 11'b10111101111;
        state_var_NS = COMP_LOOP_C_886;
      end
      COMP_LOOP_C_886 : begin
        fsm_output = 11'b10111110000;
        state_var_NS = COMP_LOOP_C_887;
      end
      COMP_LOOP_C_887 : begin
        fsm_output = 11'b10111110001;
        state_var_NS = COMP_LOOP_C_888;
      end
      COMP_LOOP_C_888 : begin
        fsm_output = 11'b10111110010;
        state_var_NS = COMP_LOOP_C_889;
      end
      COMP_LOOP_C_889 : begin
        fsm_output = 11'b10111110011;
        state_var_NS = COMP_LOOP_C_890;
      end
      COMP_LOOP_C_890 : begin
        fsm_output = 11'b10111110100;
        state_var_NS = COMP_LOOP_C_891;
      end
      COMP_LOOP_C_891 : begin
        fsm_output = 11'b10111110101;
        state_var_NS = COMP_LOOP_C_892;
      end
      COMP_LOOP_C_892 : begin
        fsm_output = 11'b10111110110;
        state_var_NS = COMP_LOOP_C_893;
      end
      COMP_LOOP_C_893 : begin
        fsm_output = 11'b10111110111;
        state_var_NS = COMP_LOOP_C_894;
      end
      COMP_LOOP_C_894 : begin
        fsm_output = 11'b10111111000;
        state_var_NS = COMP_LOOP_C_895;
      end
      COMP_LOOP_C_895 : begin
        fsm_output = 11'b10111111001;
        state_var_NS = COMP_LOOP_C_896;
      end
      COMP_LOOP_C_896 : begin
        fsm_output = 11'b10111111010;
        state_var_NS = COMP_LOOP_C_897;
      end
      COMP_LOOP_C_897 : begin
        fsm_output = 11'b10111111011;
        state_var_NS = COMP_LOOP_C_898;
      end
      COMP_LOOP_C_898 : begin
        fsm_output = 11'b10111111100;
        state_var_NS = COMP_LOOP_C_899;
      end
      COMP_LOOP_C_899 : begin
        fsm_output = 11'b10111111101;
        state_var_NS = COMP_LOOP_C_900;
      end
      COMP_LOOP_C_900 : begin
        fsm_output = 11'b10111111110;
        state_var_NS = COMP_LOOP_C_901;
      end
      COMP_LOOP_C_901 : begin
        fsm_output = 11'b10111111111;
        state_var_NS = COMP_LOOP_C_902;
      end
      COMP_LOOP_C_902 : begin
        fsm_output = 11'b11000000000;
        state_var_NS = COMP_LOOP_C_903;
      end
      COMP_LOOP_C_903 : begin
        fsm_output = 11'b11000000001;
        state_var_NS = COMP_LOOP_C_904;
      end
      COMP_LOOP_C_904 : begin
        fsm_output = 11'b11000000010;
        state_var_NS = COMP_LOOP_C_905;
      end
      COMP_LOOP_C_905 : begin
        fsm_output = 11'b11000000011;
        state_var_NS = COMP_LOOP_C_906;
      end
      COMP_LOOP_C_906 : begin
        fsm_output = 11'b11000000100;
        state_var_NS = COMP_LOOP_C_907;
      end
      COMP_LOOP_C_907 : begin
        fsm_output = 11'b11000000101;
        state_var_NS = COMP_LOOP_C_908;
      end
      COMP_LOOP_C_908 : begin
        fsm_output = 11'b11000000110;
        state_var_NS = COMP_LOOP_C_909;
      end
      COMP_LOOP_C_909 : begin
        fsm_output = 11'b11000000111;
        state_var_NS = COMP_LOOP_C_910;
      end
      COMP_LOOP_C_910 : begin
        fsm_output = 11'b11000001000;
        state_var_NS = COMP_LOOP_C_911;
      end
      COMP_LOOP_C_911 : begin
        fsm_output = 11'b11000001001;
        state_var_NS = COMP_LOOP_C_912;
      end
      COMP_LOOP_C_912 : begin
        fsm_output = 11'b11000001010;
        state_var_NS = COMP_LOOP_C_913;
      end
      COMP_LOOP_C_913 : begin
        fsm_output = 11'b11000001011;
        state_var_NS = COMP_LOOP_C_914;
      end
      COMP_LOOP_C_914 : begin
        fsm_output = 11'b11000001100;
        state_var_NS = COMP_LOOP_C_915;
      end
      COMP_LOOP_C_915 : begin
        fsm_output = 11'b11000001101;
        state_var_NS = COMP_LOOP_C_916;
      end
      COMP_LOOP_C_916 : begin
        fsm_output = 11'b11000001110;
        state_var_NS = COMP_LOOP_C_917;
      end
      COMP_LOOP_C_917 : begin
        fsm_output = 11'b11000001111;
        state_var_NS = COMP_LOOP_C_918;
      end
      COMP_LOOP_C_918 : begin
        fsm_output = 11'b11000010000;
        state_var_NS = COMP_LOOP_C_919;
      end
      COMP_LOOP_C_919 : begin
        fsm_output = 11'b11000010001;
        state_var_NS = COMP_LOOP_C_920;
      end
      COMP_LOOP_C_920 : begin
        fsm_output = 11'b11000010010;
        state_var_NS = COMP_LOOP_C_921;
      end
      COMP_LOOP_C_921 : begin
        fsm_output = 11'b11000010011;
        state_var_NS = COMP_LOOP_C_922;
      end
      COMP_LOOP_C_922 : begin
        fsm_output = 11'b11000010100;
        state_var_NS = COMP_LOOP_C_923;
      end
      COMP_LOOP_C_923 : begin
        fsm_output = 11'b11000010101;
        state_var_NS = COMP_LOOP_C_924;
      end
      COMP_LOOP_C_924 : begin
        fsm_output = 11'b11000010110;
        state_var_NS = COMP_LOOP_C_925;
      end
      COMP_LOOP_C_925 : begin
        fsm_output = 11'b11000010111;
        state_var_NS = COMP_LOOP_C_926;
      end
      COMP_LOOP_C_926 : begin
        fsm_output = 11'b11000011000;
        state_var_NS = COMP_LOOP_C_927;
      end
      COMP_LOOP_C_927 : begin
        fsm_output = 11'b11000011001;
        state_var_NS = COMP_LOOP_C_928;
      end
      COMP_LOOP_C_928 : begin
        fsm_output = 11'b11000011010;
        state_var_NS = COMP_LOOP_C_929;
      end
      COMP_LOOP_C_929 : begin
        fsm_output = 11'b11000011011;
        state_var_NS = COMP_LOOP_C_930;
      end
      COMP_LOOP_C_930 : begin
        fsm_output = 11'b11000011100;
        if ( COMP_LOOP_C_930_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_931;
        end
      end
      COMP_LOOP_C_931 : begin
        fsm_output = 11'b11000011101;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_0;
      end
      COMP_LOOP_16_modExp_1_while_C_0 : begin
        fsm_output = 11'b11000011110;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_1;
      end
      COMP_LOOP_16_modExp_1_while_C_1 : begin
        fsm_output = 11'b11000011111;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_2;
      end
      COMP_LOOP_16_modExp_1_while_C_2 : begin
        fsm_output = 11'b11000100000;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_3;
      end
      COMP_LOOP_16_modExp_1_while_C_3 : begin
        fsm_output = 11'b11000100001;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_4;
      end
      COMP_LOOP_16_modExp_1_while_C_4 : begin
        fsm_output = 11'b11000100010;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_5;
      end
      COMP_LOOP_16_modExp_1_while_C_5 : begin
        fsm_output = 11'b11000100011;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_6;
      end
      COMP_LOOP_16_modExp_1_while_C_6 : begin
        fsm_output = 11'b11000100100;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_7;
      end
      COMP_LOOP_16_modExp_1_while_C_7 : begin
        fsm_output = 11'b11000100101;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_8;
      end
      COMP_LOOP_16_modExp_1_while_C_8 : begin
        fsm_output = 11'b11000100110;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_9;
      end
      COMP_LOOP_16_modExp_1_while_C_9 : begin
        fsm_output = 11'b11000100111;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_10;
      end
      COMP_LOOP_16_modExp_1_while_C_10 : begin
        fsm_output = 11'b11000101000;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_11;
      end
      COMP_LOOP_16_modExp_1_while_C_11 : begin
        fsm_output = 11'b11000101001;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_12;
      end
      COMP_LOOP_16_modExp_1_while_C_12 : begin
        fsm_output = 11'b11000101010;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_13;
      end
      COMP_LOOP_16_modExp_1_while_C_13 : begin
        fsm_output = 11'b11000101011;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_14;
      end
      COMP_LOOP_16_modExp_1_while_C_14 : begin
        fsm_output = 11'b11000101100;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_15;
      end
      COMP_LOOP_16_modExp_1_while_C_15 : begin
        fsm_output = 11'b11000101101;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_16;
      end
      COMP_LOOP_16_modExp_1_while_C_16 : begin
        fsm_output = 11'b11000101110;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_17;
      end
      COMP_LOOP_16_modExp_1_while_C_17 : begin
        fsm_output = 11'b11000101111;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_18;
      end
      COMP_LOOP_16_modExp_1_while_C_18 : begin
        fsm_output = 11'b11000110000;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_19;
      end
      COMP_LOOP_16_modExp_1_while_C_19 : begin
        fsm_output = 11'b11000110001;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_20;
      end
      COMP_LOOP_16_modExp_1_while_C_20 : begin
        fsm_output = 11'b11000110010;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_21;
      end
      COMP_LOOP_16_modExp_1_while_C_21 : begin
        fsm_output = 11'b11000110011;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_22;
      end
      COMP_LOOP_16_modExp_1_while_C_22 : begin
        fsm_output = 11'b11000110100;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_23;
      end
      COMP_LOOP_16_modExp_1_while_C_23 : begin
        fsm_output = 11'b11000110101;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_24;
      end
      COMP_LOOP_16_modExp_1_while_C_24 : begin
        fsm_output = 11'b11000110110;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_25;
      end
      COMP_LOOP_16_modExp_1_while_C_25 : begin
        fsm_output = 11'b11000110111;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_26;
      end
      COMP_LOOP_16_modExp_1_while_C_26 : begin
        fsm_output = 11'b11000111000;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_27;
      end
      COMP_LOOP_16_modExp_1_while_C_27 : begin
        fsm_output = 11'b11000111001;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_28;
      end
      COMP_LOOP_16_modExp_1_while_C_28 : begin
        fsm_output = 11'b11000111010;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_29;
      end
      COMP_LOOP_16_modExp_1_while_C_29 : begin
        fsm_output = 11'b11000111011;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_30;
      end
      COMP_LOOP_16_modExp_1_while_C_30 : begin
        fsm_output = 11'b11000111100;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_31;
      end
      COMP_LOOP_16_modExp_1_while_C_31 : begin
        fsm_output = 11'b11000111101;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_32;
      end
      COMP_LOOP_16_modExp_1_while_C_32 : begin
        fsm_output = 11'b11000111110;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_33;
      end
      COMP_LOOP_16_modExp_1_while_C_33 : begin
        fsm_output = 11'b11000111111;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_34;
      end
      COMP_LOOP_16_modExp_1_while_C_34 : begin
        fsm_output = 11'b11001000000;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_35;
      end
      COMP_LOOP_16_modExp_1_while_C_35 : begin
        fsm_output = 11'b11001000001;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_36;
      end
      COMP_LOOP_16_modExp_1_while_C_36 : begin
        fsm_output = 11'b11001000010;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_37;
      end
      COMP_LOOP_16_modExp_1_while_C_37 : begin
        fsm_output = 11'b11001000011;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_38;
      end
      COMP_LOOP_16_modExp_1_while_C_38 : begin
        fsm_output = 11'b11001000100;
        if ( COMP_LOOP_16_modExp_1_while_C_38_tr0 ) begin
          state_var_NS = COMP_LOOP_C_932;
        end
        else begin
          state_var_NS = COMP_LOOP_16_modExp_1_while_C_0;
        end
      end
      COMP_LOOP_C_932 : begin
        fsm_output = 11'b11001000101;
        state_var_NS = COMP_LOOP_C_933;
      end
      COMP_LOOP_C_933 : begin
        fsm_output = 11'b11001000110;
        state_var_NS = COMP_LOOP_C_934;
      end
      COMP_LOOP_C_934 : begin
        fsm_output = 11'b11001000111;
        state_var_NS = COMP_LOOP_C_935;
      end
      COMP_LOOP_C_935 : begin
        fsm_output = 11'b11001001000;
        state_var_NS = COMP_LOOP_C_936;
      end
      COMP_LOOP_C_936 : begin
        fsm_output = 11'b11001001001;
        state_var_NS = COMP_LOOP_C_937;
      end
      COMP_LOOP_C_937 : begin
        fsm_output = 11'b11001001010;
        state_var_NS = COMP_LOOP_C_938;
      end
      COMP_LOOP_C_938 : begin
        fsm_output = 11'b11001001011;
        state_var_NS = COMP_LOOP_C_939;
      end
      COMP_LOOP_C_939 : begin
        fsm_output = 11'b11001001100;
        state_var_NS = COMP_LOOP_C_940;
      end
      COMP_LOOP_C_940 : begin
        fsm_output = 11'b11001001101;
        state_var_NS = COMP_LOOP_C_941;
      end
      COMP_LOOP_C_941 : begin
        fsm_output = 11'b11001001110;
        state_var_NS = COMP_LOOP_C_942;
      end
      COMP_LOOP_C_942 : begin
        fsm_output = 11'b11001001111;
        state_var_NS = COMP_LOOP_C_943;
      end
      COMP_LOOP_C_943 : begin
        fsm_output = 11'b11001010000;
        state_var_NS = COMP_LOOP_C_944;
      end
      COMP_LOOP_C_944 : begin
        fsm_output = 11'b11001010001;
        state_var_NS = COMP_LOOP_C_945;
      end
      COMP_LOOP_C_945 : begin
        fsm_output = 11'b11001010010;
        state_var_NS = COMP_LOOP_C_946;
      end
      COMP_LOOP_C_946 : begin
        fsm_output = 11'b11001010011;
        state_var_NS = COMP_LOOP_C_947;
      end
      COMP_LOOP_C_947 : begin
        fsm_output = 11'b11001010100;
        state_var_NS = COMP_LOOP_C_948;
      end
      COMP_LOOP_C_948 : begin
        fsm_output = 11'b11001010101;
        state_var_NS = COMP_LOOP_C_949;
      end
      COMP_LOOP_C_949 : begin
        fsm_output = 11'b11001010110;
        state_var_NS = COMP_LOOP_C_950;
      end
      COMP_LOOP_C_950 : begin
        fsm_output = 11'b11001010111;
        state_var_NS = COMP_LOOP_C_951;
      end
      COMP_LOOP_C_951 : begin
        fsm_output = 11'b11001011000;
        state_var_NS = COMP_LOOP_C_952;
      end
      COMP_LOOP_C_952 : begin
        fsm_output = 11'b11001011001;
        state_var_NS = COMP_LOOP_C_953;
      end
      COMP_LOOP_C_953 : begin
        fsm_output = 11'b11001011010;
        state_var_NS = COMP_LOOP_C_954;
      end
      COMP_LOOP_C_954 : begin
        fsm_output = 11'b11001011011;
        state_var_NS = COMP_LOOP_C_955;
      end
      COMP_LOOP_C_955 : begin
        fsm_output = 11'b11001011100;
        state_var_NS = COMP_LOOP_C_956;
      end
      COMP_LOOP_C_956 : begin
        fsm_output = 11'b11001011101;
        state_var_NS = COMP_LOOP_C_957;
      end
      COMP_LOOP_C_957 : begin
        fsm_output = 11'b11001011110;
        state_var_NS = COMP_LOOP_C_958;
      end
      COMP_LOOP_C_958 : begin
        fsm_output = 11'b11001011111;
        state_var_NS = COMP_LOOP_C_959;
      end
      COMP_LOOP_C_959 : begin
        fsm_output = 11'b11001100000;
        state_var_NS = COMP_LOOP_C_960;
      end
      COMP_LOOP_C_960 : begin
        fsm_output = 11'b11001100001;
        state_var_NS = COMP_LOOP_C_961;
      end
      COMP_LOOP_C_961 : begin
        fsm_output = 11'b11001100010;
        state_var_NS = COMP_LOOP_C_962;
      end
      COMP_LOOP_C_962 : begin
        fsm_output = 11'b11001100011;
        state_var_NS = COMP_LOOP_C_963;
      end
      COMP_LOOP_C_963 : begin
        fsm_output = 11'b11001100100;
        state_var_NS = COMP_LOOP_C_964;
      end
      COMP_LOOP_C_964 : begin
        fsm_output = 11'b11001100101;
        state_var_NS = COMP_LOOP_C_965;
      end
      COMP_LOOP_C_965 : begin
        fsm_output = 11'b11001100110;
        state_var_NS = COMP_LOOP_C_966;
      end
      COMP_LOOP_C_966 : begin
        fsm_output = 11'b11001100111;
        state_var_NS = COMP_LOOP_C_967;
      end
      COMP_LOOP_C_967 : begin
        fsm_output = 11'b11001101000;
        state_var_NS = COMP_LOOP_C_968;
      end
      COMP_LOOP_C_968 : begin
        fsm_output = 11'b11001101001;
        state_var_NS = COMP_LOOP_C_969;
      end
      COMP_LOOP_C_969 : begin
        fsm_output = 11'b11001101010;
        state_var_NS = COMP_LOOP_C_970;
      end
      COMP_LOOP_C_970 : begin
        fsm_output = 11'b11001101011;
        state_var_NS = COMP_LOOP_C_971;
      end
      COMP_LOOP_C_971 : begin
        fsm_output = 11'b11001101100;
        state_var_NS = COMP_LOOP_C_972;
      end
      COMP_LOOP_C_972 : begin
        fsm_output = 11'b11001101101;
        state_var_NS = COMP_LOOP_C_973;
      end
      COMP_LOOP_C_973 : begin
        fsm_output = 11'b11001101110;
        state_var_NS = COMP_LOOP_C_974;
      end
      COMP_LOOP_C_974 : begin
        fsm_output = 11'b11001101111;
        state_var_NS = COMP_LOOP_C_975;
      end
      COMP_LOOP_C_975 : begin
        fsm_output = 11'b11001110000;
        state_var_NS = COMP_LOOP_C_976;
      end
      COMP_LOOP_C_976 : begin
        fsm_output = 11'b11001110001;
        state_var_NS = COMP_LOOP_C_977;
      end
      COMP_LOOP_C_977 : begin
        fsm_output = 11'b11001110010;
        state_var_NS = COMP_LOOP_C_978;
      end
      COMP_LOOP_C_978 : begin
        fsm_output = 11'b11001110011;
        state_var_NS = COMP_LOOP_C_979;
      end
      COMP_LOOP_C_979 : begin
        fsm_output = 11'b11001110100;
        state_var_NS = COMP_LOOP_C_980;
      end
      COMP_LOOP_C_980 : begin
        fsm_output = 11'b11001110101;
        state_var_NS = COMP_LOOP_C_981;
      end
      COMP_LOOP_C_981 : begin
        fsm_output = 11'b11001110110;
        state_var_NS = COMP_LOOP_C_982;
      end
      COMP_LOOP_C_982 : begin
        fsm_output = 11'b11001110111;
        state_var_NS = COMP_LOOP_C_983;
      end
      COMP_LOOP_C_983 : begin
        fsm_output = 11'b11001111000;
        state_var_NS = COMP_LOOP_C_984;
      end
      COMP_LOOP_C_984 : begin
        fsm_output = 11'b11001111001;
        state_var_NS = COMP_LOOP_C_985;
      end
      COMP_LOOP_C_985 : begin
        fsm_output = 11'b11001111010;
        state_var_NS = COMP_LOOP_C_986;
      end
      COMP_LOOP_C_986 : begin
        fsm_output = 11'b11001111011;
        state_var_NS = COMP_LOOP_C_987;
      end
      COMP_LOOP_C_987 : begin
        fsm_output = 11'b11001111100;
        state_var_NS = COMP_LOOP_C_988;
      end
      COMP_LOOP_C_988 : begin
        fsm_output = 11'b11001111101;
        state_var_NS = COMP_LOOP_C_989;
      end
      COMP_LOOP_C_989 : begin
        fsm_output = 11'b11001111110;
        state_var_NS = COMP_LOOP_C_990;
      end
      COMP_LOOP_C_990 : begin
        fsm_output = 11'b11001111111;
        state_var_NS = COMP_LOOP_C_991;
      end
      COMP_LOOP_C_991 : begin
        fsm_output = 11'b11010000000;
        state_var_NS = COMP_LOOP_C_992;
      end
      COMP_LOOP_C_992 : begin
        fsm_output = 11'b11010000001;
        if ( COMP_LOOP_C_992_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_0;
        end
      end
      VEC_LOOP_C_0 : begin
        fsm_output = 11'b11010000010;
        if ( VEC_LOOP_C_0_tr0 ) begin
          state_var_NS = STAGE_LOOP_C_9;
        end
        else begin
          state_var_NS = COMP_LOOP_C_0;
        end
      end
      STAGE_LOOP_C_9 : begin
        fsm_output = 11'b11010000011;
        if ( STAGE_LOOP_C_9_tr0 ) begin
          state_var_NS = main_C_1;
        end
        else begin
          state_var_NS = STAGE_LOOP_C_0;
        end
      end
      main_C_1 : begin
        fsm_output = 11'b11010000100;
        state_var_NS = main_C_0;
      end
      // main_C_0
      default : begin
        fsm_output = 11'b00000000000;
        state_var_NS = STAGE_LOOP_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( rst ) begin
      state_var <= main_C_0;
    end
    else begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_core
// ------------------------------------------------------------------


module inPlaceNTT_DIT_core (
  clk, rst, vec_rsc_triosy_0_0_lz, vec_rsc_triosy_0_1_lz, vec_rsc_triosy_0_2_lz,
      vec_rsc_triosy_0_3_lz, vec_rsc_triosy_0_4_lz, vec_rsc_triosy_0_5_lz, vec_rsc_triosy_0_6_lz,
      vec_rsc_triosy_0_7_lz, vec_rsc_triosy_0_8_lz, vec_rsc_triosy_0_9_lz, vec_rsc_triosy_0_10_lz,
      vec_rsc_triosy_0_11_lz, vec_rsc_triosy_0_12_lz, vec_rsc_triosy_0_13_lz, vec_rsc_triosy_0_14_lz,
      vec_rsc_triosy_0_15_lz, p_rsc_dat, p_rsc_triosy_lz, r_rsc_dat, r_rsc_triosy_lz,
      vec_rsc_0_0_i_qa_d, vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d, vec_rsc_0_1_i_qa_d,
      vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d, vec_rsc_0_2_i_qa_d, vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_3_i_qa_d, vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d, vec_rsc_0_4_i_qa_d,
      vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d, vec_rsc_0_5_i_qa_d, vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_6_i_qa_d, vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d, vec_rsc_0_7_i_qa_d,
      vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d, vec_rsc_0_8_i_qa_d, vec_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_9_i_qa_d, vec_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d, vec_rsc_0_10_i_qa_d,
      vec_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d, vec_rsc_0_11_i_qa_d, vec_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_12_i_qa_d, vec_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d, vec_rsc_0_13_i_qa_d,
      vec_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d, vec_rsc_0_14_i_qa_d, vec_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_15_i_qa_d, vec_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d, vec_rsc_0_0_i_adra_d_pff,
      vec_rsc_0_0_i_da_d_pff, vec_rsc_0_0_i_wea_d_pff, vec_rsc_0_1_i_wea_d_pff, vec_rsc_0_2_i_wea_d_pff,
      vec_rsc_0_3_i_wea_d_pff, vec_rsc_0_4_i_wea_d_pff, vec_rsc_0_5_i_wea_d_pff,
      vec_rsc_0_6_i_wea_d_pff, vec_rsc_0_7_i_wea_d_pff, vec_rsc_0_8_i_wea_d_pff,
      vec_rsc_0_9_i_wea_d_pff, vec_rsc_0_10_i_wea_d_pff, vec_rsc_0_11_i_wea_d_pff,
      vec_rsc_0_12_i_wea_d_pff, vec_rsc_0_13_i_wea_d_pff, vec_rsc_0_14_i_wea_d_pff,
      vec_rsc_0_15_i_wea_d_pff
);
  input clk;
  input rst;
  output vec_rsc_triosy_0_0_lz;
  output vec_rsc_triosy_0_1_lz;
  output vec_rsc_triosy_0_2_lz;
  output vec_rsc_triosy_0_3_lz;
  output vec_rsc_triosy_0_4_lz;
  output vec_rsc_triosy_0_5_lz;
  output vec_rsc_triosy_0_6_lz;
  output vec_rsc_triosy_0_7_lz;
  output vec_rsc_triosy_0_8_lz;
  output vec_rsc_triosy_0_9_lz;
  output vec_rsc_triosy_0_10_lz;
  output vec_rsc_triosy_0_11_lz;
  output vec_rsc_triosy_0_12_lz;
  output vec_rsc_triosy_0_13_lz;
  output vec_rsc_triosy_0_14_lz;
  output vec_rsc_triosy_0_15_lz;
  input [63:0] p_rsc_dat;
  output p_rsc_triosy_lz;
  input [63:0] r_rsc_dat;
  output r_rsc_triosy_lz;
  input [63:0] vec_rsc_0_0_i_qa_d;
  output vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_1_i_qa_d;
  output vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_2_i_qa_d;
  output vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_3_i_qa_d;
  output vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_4_i_qa_d;
  output vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_5_i_qa_d;
  output vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_6_i_qa_d;
  output vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_7_i_qa_d;
  output vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_8_i_qa_d;
  output vec_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_9_i_qa_d;
  output vec_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_10_i_qa_d;
  output vec_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_11_i_qa_d;
  output vec_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_12_i_qa_d;
  output vec_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_13_i_qa_d;
  output vec_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_14_i_qa_d;
  output vec_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_15_i_qa_d;
  output vec_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] vec_rsc_0_0_i_adra_d_pff;
  output [63:0] vec_rsc_0_0_i_da_d_pff;
  output vec_rsc_0_0_i_wea_d_pff;
  output vec_rsc_0_1_i_wea_d_pff;
  output vec_rsc_0_2_i_wea_d_pff;
  output vec_rsc_0_3_i_wea_d_pff;
  output vec_rsc_0_4_i_wea_d_pff;
  output vec_rsc_0_5_i_wea_d_pff;
  output vec_rsc_0_6_i_wea_d_pff;
  output vec_rsc_0_7_i_wea_d_pff;
  output vec_rsc_0_8_i_wea_d_pff;
  output vec_rsc_0_9_i_wea_d_pff;
  output vec_rsc_0_10_i_wea_d_pff;
  output vec_rsc_0_11_i_wea_d_pff;
  output vec_rsc_0_12_i_wea_d_pff;
  output vec_rsc_0_13_i_wea_d_pff;
  output vec_rsc_0_14_i_wea_d_pff;
  output vec_rsc_0_15_i_wea_d_pff;


  // Interconnect Declarations
  wire [63:0] p_rsci_idat;
  wire [63:0] r_rsci_idat;
  reg [63:0] modulo_result_rem_cmp_a;
  reg [63:0] modulo_result_rem_cmp_b;
  wire [63:0] modulo_result_rem_cmp_z;
  reg [64:0] operator_66_true_div_cmp_a;
  wire [64:0] operator_66_true_div_cmp_z;
  reg [9:0] operator_66_true_div_cmp_b_9_0;
  wire [10:0] fsm_output;
  wire or_tmp_3;
  wire or_tmp_4;
  wire or_tmp_8;
  wire or_tmp_9;
  wire or_tmp_14;
  wire nor_tmp_6;
  wire or_tmp_21;
  wire nor_tmp_9;
  wire not_tmp_34;
  wire not_tmp_45;
  wire or_tmp_110;
  wire not_tmp_51;
  wire or_tmp_118;
  wire or_tmp_141;
  wire mux_tmp_207;
  wire mux_tmp_226;
  wire or_tmp_150;
  wire or_tmp_178;
  wire or_tmp_179;
  wire or_tmp_180;
  wire or_tmp_181;
  wire mux_tmp_373;
  wire or_tmp_182;
  wire mux_tmp_374;
  wire mux_tmp_375;
  wire or_tmp_183;
  wire mux_tmp_378;
  wire mux_tmp_379;
  wire mux_tmp_380;
  wire mux_tmp_381;
  wire nor_tmp_46;
  wire nand_tmp_12;
  wire nand_tmp_13;
  wire or_tmp_187;
  wire mux_tmp_399;
  wire or_tmp_188;
  wire or_tmp_189;
  wire or_tmp_191;
  wire nand_tmp_14;
  wire or_tmp_195;
  wire mux_tmp_412;
  wire mux_tmp_413;
  wire and_dcpl;
  wire and_dcpl_1;
  wire and_dcpl_2;
  wire or_tmp_237;
  wire nor_tmp_116;
  wire mux_tmp_741;
  wire or_tmp_434;
  wire mux_tmp_893;
  wire mux_tmp_917;
  wire and_dcpl_21;
  wire and_dcpl_22;
  wire and_dcpl_26;
  wire and_dcpl_30;
  wire and_dcpl_31;
  wire and_dcpl_32;
  wire and_dcpl_40;
  wire and_dcpl_46;
  wire and_dcpl_50;
  wire not_tmp_219;
  wire and_dcpl_96;
  wire and_dcpl_97;
  wire and_dcpl_98;
  wire and_dcpl_99;
  wire and_dcpl_100;
  wire and_dcpl_101;
  wire and_dcpl_102;
  wire and_dcpl_103;
  wire and_dcpl_106;
  wire and_dcpl_107;
  wire and_dcpl_108;
  wire and_dcpl_109;
  wire and_dcpl_110;
  wire and_dcpl_111;
  wire and_dcpl_116;
  wire and_dcpl_117;
  wire and_dcpl_118;
  wire and_dcpl_119;
  wire and_dcpl_121;
  wire and_dcpl_122;
  wire and_dcpl_123;
  wire and_dcpl_124;
  wire and_dcpl_125;
  wire and_dcpl_126;
  wire and_dcpl_127;
  wire and_dcpl_128;
  wire and_dcpl_129;
  wire or_tmp_453;
  wire not_tmp_240;
  wire and_dcpl_139;
  wire and_dcpl_140;
  wire and_dcpl_141;
  wire and_dcpl_145;
  wire and_dcpl_146;
  wire and_dcpl_147;
  wire and_dcpl_148;
  wire and_dcpl_154;
  wire and_dcpl_156;
  wire and_dcpl_158;
  wire and_dcpl_162;
  wire and_dcpl_164;
  wire and_dcpl_165;
  wire nor_tmp_217;
  wire mux_tmp_1049;
  wire and_dcpl_172;
  wire and_dcpl_173;
  wire and_dcpl_175;
  wire and_dcpl_182;
  wire and_dcpl_191;
  wire and_dcpl_192;
  wire and_dcpl_198;
  wire and_dcpl_204;
  wire and_dcpl_206;
  wire and_dcpl_215;
  wire and_dcpl_217;
  wire and_dcpl_223;
  wire and_dcpl_225;
  wire and_dcpl_232;
  wire and_dcpl_239;
  wire and_dcpl_240;
  wire and_dcpl_242;
  wire and_dcpl_243;
  wire and_dcpl_245;
  wire and_dcpl_247;
  wire and_dcpl_255;
  wire or_tmp_515;
  wire or_tmp_518;
  wire mux_tmp_1062;
  wire mux_tmp_1067;
  wire mux_tmp_1068;
  wire not_tmp_260;
  wire or_tmp_626;
  wire or_tmp_630;
  wire mux_tmp_1139;
  wire mux_tmp_1150;
  wire mux_tmp_1152;
  wire or_tmp_728;
  wire or_tmp_731;
  wire mux_tmp_1206;
  wire mux_tmp_1211;
  wire mux_tmp_1212;
  wire or_tmp_839;
  wire or_tmp_843;
  wire mux_tmp_1283;
  wire mux_tmp_1294;
  wire mux_tmp_1296;
  wire or_tmp_941;
  wire or_tmp_944;
  wire mux_tmp_1350;
  wire mux_tmp_1355;
  wire mux_tmp_1356;
  wire or_tmp_1052;
  wire or_tmp_1056;
  wire mux_tmp_1427;
  wire mux_tmp_1438;
  wire mux_tmp_1440;
  wire or_tmp_1154;
  wire or_tmp_1157;
  wire mux_tmp_1494;
  wire mux_tmp_1499;
  wire mux_tmp_1500;
  wire or_tmp_1265;
  wire or_tmp_1269;
  wire mux_tmp_1571;
  wire mux_tmp_1582;
  wire mux_tmp_1584;
  wire or_tmp_1367;
  wire or_tmp_1370;
  wire mux_tmp_1638;
  wire mux_tmp_1643;
  wire mux_tmp_1644;
  wire or_tmp_1478;
  wire or_tmp_1482;
  wire mux_tmp_1715;
  wire mux_tmp_1726;
  wire mux_tmp_1728;
  wire or_tmp_1580;
  wire or_tmp_1583;
  wire mux_tmp_1782;
  wire mux_tmp_1787;
  wire mux_tmp_1788;
  wire or_tmp_1691;
  wire or_tmp_1695;
  wire mux_tmp_1859;
  wire mux_tmp_1870;
  wire mux_tmp_1872;
  wire or_tmp_1797;
  wire not_tmp_378;
  wire mux_tmp_1927;
  wire nand_tmp_74;
  wire or_tmp_1811;
  wire or_tmp_1812;
  wire not_tmp_381;
  wire or_tmp_1821;
  wire or_tmp_1907;
  wire or_tmp_1911;
  wire mux_tmp_2004;
  wire mux_tmp_2015;
  wire mux_tmp_2017;
  wire or_tmp_2009;
  wire or_tmp_2012;
  wire mux_tmp_2071;
  wire mux_tmp_2076;
  wire mux_tmp_2077;
  wire or_tmp_2120;
  wire or_tmp_2124;
  wire mux_tmp_2148;
  wire mux_tmp_2159;
  wire mux_tmp_2161;
  wire and_dcpl_260;
  wire or_tmp_2220;
  wire or_tmp_2223;
  wire or_tmp_2225;
  wire or_tmp_2230;
  wire or_tmp_2233;
  wire mux_tmp_2218;
  wire mux_tmp_2220;
  wire mux_tmp_2223;
  wire or_tmp_2237;
  wire or_tmp_2238;
  wire mux_tmp_2239;
  wire nand_tmp_92;
  wire nor_tmp_286;
  wire or_tmp_2246;
  wire or_tmp_2248;
  wire not_tmp_426;
  wire nor_tmp_288;
  wire and_tmp_10;
  wire mux_tmp_2250;
  wire mux_tmp_2251;
  wire mux_tmp_2254;
  wire or_tmp_2253;
  wire or_tmp_2255;
  wire mux_tmp_2265;
  wire nor_tmp_291;
  wire or_tmp_2257;
  wire nor_tmp_295;
  wire mux_tmp_2285;
  wire mux_tmp_2290;
  wire or_tmp_2260;
  wire or_tmp_2263;
  wire nand_tmp_93;
  wire or_tmp_2266;
  wire mux_tmp_2309;
  wire or_tmp_2267;
  wire or_tmp_2269;
  wire nand_tmp_95;
  wire or_tmp_2271;
  wire nand_tmp_96;
  wire or_tmp_2275;
  wire or_tmp_2276;
  wire or_tmp_2277;
  wire mux_tmp_2327;
  wire or_tmp_2280;
  wire or_tmp_2281;
  wire or_tmp_2282;
  wire or_tmp_2289;
  wire not_tmp_463;
  wire mux_tmp_2349;
  wire and_tmp_16;
  wire or_tmp_2293;
  wire mux_tmp_2362;
  wire nor_tmp_300;
  wire or_tmp_2327;
  wire or_tmp_2329;
  wire or_tmp_2331;
  wire or_tmp_2333;
  wire or_tmp_2334;
  wire mux_tmp_2400;
  wire mux_tmp_2401;
  wire mux_tmp_2402;
  wire or_tmp_2335;
  wire mux_tmp_2406;
  wire or_tmp_2338;
  wire nand_tmp_105;
  wire mux_tmp_2423;
  wire nor_tmp_307;
  wire mux_tmp_2425;
  wire mux_tmp_2426;
  wire or_tmp_2342;
  wire or_tmp_2343;
  wire mux_tmp_2436;
  wire nand_tmp_107;
  wire nand_tmp_108;
  wire mux_tmp_2466;
  wire not_tmp_519;
  wire and_dcpl_264;
  wire and_dcpl_266;
  wire and_dcpl_268;
  wire and_dcpl_273;
  wire mux_tmp_2502;
  wire not_tmp_529;
  wire nor_tmp_330;
  wire mux_tmp_2508;
  wire or_tmp_2416;
  wire or_tmp_2419;
  wire mux_tmp_2519;
  wire mux_tmp_2523;
  wire mux_tmp_2525;
  wire nor_tmp_338;
  wire or_tmp_2429;
  wire nor_tmp_342;
  wire mux_tmp_2549;
  wire mux_tmp_2650;
  wire and_dcpl_279;
  wire and_dcpl_281;
  wire mux_tmp_2687;
  wire or_tmp_2474;
  wire mux_tmp_2696;
  wire mux_tmp_2698;
  wire mux_tmp_2701;
  wire or_tmp_2479;
  wire nand_tmp_119;
  wire or_tmp_2483;
  wire and_dcpl_283;
  wire and_dcpl_305;
  wire not_tmp_596;
  wire or_tmp_2516;
  wire mux_tmp_2758;
  wire mux_tmp_2788;
  wire mux_tmp_2790;
  wire mux_tmp_2796;
  wire mux_tmp_2800;
  wire mux_tmp_2813;
  wire or_tmp_2594;
  wire not_tmp_634;
  wire or_tmp_2631;
  wire not_tmp_646;
  wire or_tmp_2649;
  wire nand_tmp_136;
  wire mux_tmp_2905;
  wire nand_tmp_137;
  wire mux_tmp_2907;
  wire or_tmp_2652;
  wire or_tmp_2653;
  wire mux_tmp_2911;
  wire mux_tmp_2912;
  wire mux_tmp_2913;
  wire mux_tmp_2919;
  wire mux_tmp_2921;
  wire mux_tmp_2930;
  wire or_tmp_2659;
  wire or_tmp_2663;
  wire nand_tmp_140;
  wire or_tmp_2707;
  wire and_dcpl_332;
  wire nand_tmp_148;
  wire not_tmp_708;
  wire nor_tmp_445;
  wire mux_tmp_3219;
  wire mux_tmp_3236;
  wire or_tmp_2849;
  wire mux_tmp_3244;
  wire nor_tmp_456;
  wire mux_tmp_3256;
  wire not_tmp_728;
  wire or_tmp_2864;
  wire mux_tmp_3269;
  wire nor_tmp_461;
  wire mux_tmp_3280;
  wire mux_tmp_3281;
  wire nand_tmp_157;
  wire mux_tmp_3323;
  wire not_tmp_762;
  wire mux_tmp_3386;
  wire not_tmp_776;
  wire mux_tmp_3418;
  wire mux_tmp_3422;
  wire mux_tmp_3426;
  wire mux_tmp_3430;
  wire mux_tmp_3436;
  wire nand_tmp_167;
  wire mux_tmp_3449;
  wire mux_tmp_3450;
  wire mux_tmp_3452;
  wire mux_tmp_3456;
  wire mux_tmp_3458;
  wire mux_tmp_3459;
  wire mux_tmp_3467;
  wire mux_tmp_3468;
  wire mux_tmp_3471;
  wire and_tmp_36;
  wire or_tmp_3025;
  wire or_tmp_3107;
  reg COMP_LOOP_COMP_LOOP_and_137_itm;
  reg COMP_LOOP_COMP_LOOP_and_10_itm;
  reg COMP_LOOP_nor_11_itm;
  wire [11:0] COMP_LOOP_acc_1_cse_6_sva_1;
  wire [12:0] nl_COMP_LOOP_acc_1_cse_6_sva_1;
  reg [11:0] VEC_LOOP_j_sva_11_0;
  reg [4:0] COMP_LOOP_k_9_4_sva_4_0;
  reg COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm;
  reg COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  wire [5:0] COMP_LOOP_k_9_4_sva_2;
  wire [6:0] nl_COMP_LOOP_k_9_4_sva_2;
  reg [11:0] COMP_LOOP_acc_10_cse_12_1_1_sva;
  reg [11:0] COMP_LOOP_acc_1_cse_2_sva;
  reg [9:0] COMP_LOOP_acc_19_psp_sva;
  reg [9:0] COMP_LOOP_acc_13_psp_sva;
  reg [11:0] COMP_LOOP_acc_1_cse_10_sva;
  wire [12:0] nl_COMP_LOOP_acc_1_cse_10_sva;
  reg [11:0] COMP_LOOP_acc_1_cse_14_sva;
  wire [12:0] nl_COMP_LOOP_acc_1_cse_14_sva;
  reg [8:0] COMP_LOOP_acc_16_psp_sva;
  reg [11:0] COMP_LOOP_acc_1_cse_6_sva;
  reg [10:0] COMP_LOOP_acc_17_psp_sva;
  wire [11:0] nl_COMP_LOOP_acc_17_psp_sva;
  reg [11:0] COMP_LOOP_acc_1_cse_sva;
  wire [12:0] nl_COMP_LOOP_acc_1_cse_sva;
  reg [11:0] COMP_LOOP_acc_1_cse_8_sva;
  wire [12:0] nl_COMP_LOOP_acc_1_cse_8_sva;
  reg [10:0] COMP_LOOP_acc_11_psp_sva;
  wire [11:0] nl_COMP_LOOP_acc_11_psp_sva;
  reg [11:0] COMP_LOOP_acc_1_cse_4_sva;
  reg [11:0] COMP_LOOP_acc_1_cse_12_sva;
  wire [12:0] nl_COMP_LOOP_acc_1_cse_12_sva;
  reg [10:0] COMP_LOOP_acc_14_psp_sva;
  wire [11:0] nl_COMP_LOOP_acc_14_psp_sva;
  reg [10:0] COMP_LOOP_acc_20_psp_sva;
  wire [11:0] nl_COMP_LOOP_acc_20_psp_sva;
  reg [63:0] tmp_10_lpi_4_dfm;
  wire [11:0] COMP_LOOP_acc_1_cse_2_sva_1;
  wire [12:0] nl_COMP_LOOP_acc_1_cse_2_sva_1;
  wire mux_2770_m1c;
  wire and_305_m1c;
  wire and_307_m1c;
  wire and_309_m1c;
  wire and_312_m1c;
  wire and_315_m1c;
  wire and_317_m1c;
  wire and_320_m1c;
  wire and_322_m1c;
  wire and_324_m1c;
  wire and_327_m1c;
  wire and_329_m1c;
  wire and_331_m1c;
  wire and_334_m1c;
  wire and_336_m1c;
  wire and_339_m1c;
  wire and_300_m1c;
  wire nor_223_cse;
  reg reg_vec_rsc_triosy_0_15_obj_ld_cse;
  wire and_574_cse;
  wire or_2348_cse;
  wire and_573_cse;
  wire nand_375_cse;
  wire or_495_cse;
  wire nand_376_cse;
  wire nor_412_cse;
  wire and_563_cse;
  wire or_2385_cse;
  wire or_2894_cse;
  wire and_517_cse;
  wire and_528_cse;
  wire and_565_cse;
  wire and_456_cse;
  wire and_458_cse;
  wire or_3328_cse;
  wire or_2520_cse;
  wire nor_1203_cse;
  wire or_2935_cse;
  wire nand_398_cse;
  wire or_2679_cse;
  wire nor_381_cse;
  wire nor_670_cse;
  wire nand_237_cse;
  wire [63:0] modulo_result_mux_1_cse;
  wire nor_544_cse;
  wire or_212_cse;
  wire nor_422_cse;
  wire and_472_cse;
  wire and_491_cse;
  wire and_816_cse;
  wire mux_726_cse;
  wire nor_601_cse;
  wire nor_610_cse;
  wire or_622_cse;
  wire or_617_cse;
  wire mux_1088_cse;
  wire or_609_cse;
  wire or_607_cse;
  wire nand_25_cse;
  wire or_601_cse;
  wire mux_1073_cse;
  wire or_2898_cse;
  wire or_15_cse;
  wire nor_784_cse;
  wire or_2824_cse;
  wire or_529_cse;
  wire nand_226_cse;
  wire or_2826_cse;
  wire or_2839_cse;
  wire nor_1276_cse;
  wire nor_1279_cse;
  wire and_459_cse;
  wire and_440_cse;
  wire nand_402_cse;
  wire and_815_cse;
  wire nor_539_cse;
  wire mux_71_cse;
  wire and_464_cse;
  wire or_525_cse;
  wire nand_240_cse;
  wire mux_3498_cse;
  wire or_154_cse;
  wire or_2951_cse;
  wire nor_1316_cse;
  wire and_450_cse;
  wire nor_515_cse;
  wire mux_2746_cse;
  wire or_3002_cse;
  wire or_163_cse;
  wire or_3308_cse;
  wire or_3279_cse;
  wire or_621_cse;
  wire or_596_cse;
  wire and_359_cse;
  wire mux_3394_cse;
  wire mux_3385_cse;
  wire or_2729_cse;
  wire and_754_cse;
  wire mux_28_cse;
  wire or_2902_cse;
  wire or_36_cse;
  wire or_2819_cse;
  wire mux_3_cse;
  wire mux_7_cse;
  wire mux_9_cse;
  wire mux_3143_cse;
  wire mux_2463_cse;
  wire mux_3603_cse;
  wire nor_545_cse;
  wire or_3018_cse;
  wire or_3016_cse;
  wire mux_3392_cse;
  wire and_540_cse;
  wire mux_3388_cse;
  wire mux_384_cse;
  wire mux_382_cse;
  wire mux_3557_cse;
  wire mux_3575_cse;
  wire mux_3555_cse;
  wire mux_3551_cse;
  wire [7:0] COMP_LOOP_acc_psp_sva_1;
  wire [8:0] nl_COMP_LOOP_acc_psp_sva_1;
  reg [7:0] COMP_LOOP_acc_psp_sva;
  wire mux_2433_itm;
  wire mux_2435_itm;
  wire mux_2475_itm;
  wire mux_3369_itm;
  wire and_dcpl_348;
  wire and_dcpl_350;
  wire and_dcpl_351;
  wire and_dcpl_353;
  wire and_dcpl_354;
  wire and_dcpl_356;
  wire and_dcpl_358;
  wire and_dcpl_359;
  wire and_dcpl_361;
  wire and_dcpl_365;
  wire and_dcpl_368;
  wire and_dcpl_373;
  wire and_dcpl_374;
  wire and_dcpl_375;
  wire and_dcpl_376;
  wire and_dcpl_378;
  wire and_dcpl_380;
  wire and_dcpl_384;
  wire and_dcpl_386;
  wire and_dcpl_391;
  wire and_dcpl_392;
  wire and_dcpl_394;
  wire and_dcpl_397;
  wire and_dcpl_401;
  wire and_dcpl_404;
  wire and_dcpl_406;
  wire and_dcpl_408;
  wire and_dcpl_411;
  wire and_dcpl_415;
  wire [9:0] z_out;
  wire and_dcpl_430;
  wire and_dcpl_433;
  wire and_dcpl_441;
  wire [9:0] z_out_1;
  wire [10:0] nl_z_out_1;
  wire [9:0] z_out_2;
  wire [10:0] nl_z_out_2;
  wire and_dcpl_480;
  wire and_dcpl_502;
  wire and_dcpl_503;
  wire and_dcpl_511;
  wire [9:0] z_out_3;
  wire [10:0] nl_z_out_3;
  wire and_dcpl_517;
  wire [9:0] z_out_4;
  wire [10:0] nl_z_out_4;
  wire and_dcpl_555;
  wire not_tmp_930;
  wire mux_tmp;
  wire not_tmp_933;
  wire and_dcpl_564;
  wire [63:0] z_out_5;
  wire [64:0] nl_z_out_5;
  wire and_dcpl_568;
  wire and_dcpl_574;
  wire or_tmp_3188;
  wire or_tmp_3189;
  wire mux_tmp_3724;
  wire or_tmp_3191;
  wire or_tmp_3193;
  wire mux_tmp_3725;
  wire or_tmp_3195;
  wire or_tmp_3196;
  wire mux_tmp_3728;
  wire or_tmp_3200;
  wire or_tmp_3202;
  wire or_tmp_3203;
  wire mux_tmp_3733;
  wire or_tmp_3204;
  wire or_tmp_3205;
  wire mux_tmp_3735;
  wire mux_tmp_3737;
  wire or_tmp_3211;
  wire mux_tmp_3742;
  wire or_tmp_3212;
  wire mux_tmp_3743;
  wire or_tmp_3213;
  wire or_tmp_3218;
  wire mux_tmp_3751;
  wire mux_tmp_3753;
  wire mux_tmp_3762;
  wire mux_tmp_3771;
  wire and_dcpl_579;
  wire and_dcpl_588;
  wire [64:0] z_out_6;
  wire [65:0] nl_z_out_6;
  wire and_dcpl_591;
  wire and_dcpl_592;
  wire and_dcpl_598;
  wire and_dcpl_614;
  wire and_dcpl_615;
  wire and_dcpl_618;
  wire and_dcpl_622;
  wire and_dcpl_623;
  wire and_dcpl_624;
  wire and_dcpl_628;
  wire and_dcpl_641;
  wire and_dcpl_642;
  wire and_dcpl_646;
  wire and_dcpl_651;
  wire and_dcpl_654;
  wire and_dcpl_657;
  wire and_dcpl_659;
  wire and_dcpl_663;
  wire and_dcpl_666;
  wire and_dcpl_669;
  wire and_dcpl_672;
  wire and_dcpl_676;
  wire and_dcpl_678;
  wire [64:0] z_out_7;
  wire [65:0] nl_z_out_7;
  wire and_dcpl_688;
  wire and_dcpl_698;
  wire not_tmp_980;
  wire and_dcpl_707;
  wire and_dcpl_717;
  wire and_dcpl_727;
  wire and_dcpl_734;
  wire and_dcpl_741;
  wire [6:0] z_out_9;
  wire [63:0] z_out_10;
  wire signed [128:0] nl_z_out_10;
  reg [63:0] p_sva;
  reg [63:0] r_sva;
  reg [3:0] STAGE_LOOP_i_3_0_sva;
  reg [9:0] STAGE_LOOP_lshift_psp_sva;
  reg [63:0] modExp_result_sva;
  reg modExp_exp_1_7_1_sva;
  reg modExp_exp_1_6_1_sva;
  reg modExp_exp_1_5_1_sva;
  reg modExp_exp_1_4_1_sva;
  reg [63:0] COMP_LOOP_10_mul_mut;
  reg COMP_LOOP_COMP_LOOP_nor_itm;
  reg COMP_LOOP_COMP_LOOP_and_2_itm;
  reg COMP_LOOP_COMP_LOOP_and_4_itm;
  reg COMP_LOOP_COMP_LOOP_and_5_itm;
  reg COMP_LOOP_COMP_LOOP_and_6_itm;
  reg COMP_LOOP_COMP_LOOP_and_8_itm;
  reg COMP_LOOP_COMP_LOOP_and_9_itm;
  reg COMP_LOOP_COMP_LOOP_and_11_itm;
  reg COMP_LOOP_COMP_LOOP_and_12_itm;
  reg COMP_LOOP_COMP_LOOP_and_13_itm;
  reg COMP_LOOP_COMP_LOOP_and_14_itm;
  reg COMP_LOOP_COMP_LOOP_nor_1_itm;
  reg COMP_LOOP_nor_12_itm;
  reg COMP_LOOP_COMP_LOOP_and_62_itm;
  reg COMP_LOOP_COMP_LOOP_and_64_itm;
  reg COMP_LOOP_COMP_LOOP_and_68_itm;
  reg COMP_LOOP_COMP_LOOP_and_139_itm;
  reg COMP_LOOP_COMP_LOOP_and_140_itm;
  reg COMP_LOOP_COMP_LOOP_and_141_itm;
  reg COMP_LOOP_COMP_LOOP_and_143_itm;
  reg COMP_LOOP_COMP_LOOP_and_144_itm;
  reg COMP_LOOP_COMP_LOOP_and_145_itm;
  reg COMP_LOOP_COMP_LOOP_and_146_itm;
  reg COMP_LOOP_COMP_LOOP_and_147_itm;
  reg COMP_LOOP_COMP_LOOP_and_148_itm;
  reg COMP_LOOP_COMP_LOOP_and_149_itm;
  reg COMP_LOOP_nor_134_itm;
  reg COMP_LOOP_nor_137_itm;
  reg COMP_LOOP_COMP_LOOP_and_305_itm;
  reg [63:0] COMP_LOOP_10_acc_8_itm;
  wire STAGE_LOOP_i_3_0_sva_mx0c1;
  wire [3:0] STAGE_LOOP_i_3_0_sva_2;
  wire [4:0] nl_STAGE_LOOP_i_3_0_sva_2;
  wire [63:0] COMP_LOOP_1_modExp_1_while_if_mul_mut_1;
  wire signed [127:0] nl_COMP_LOOP_1_modExp_1_while_if_mul_mut_1;
  wire [9:0] STAGE_LOOP_lshift_psp_sva_mx0w0;
  wire VEC_LOOP_j_sva_11_0_mx0c1;
  wire modExp_result_sva_mx0c0;
  wire [62:0] operator_64_false_slc_modExp_exp_63_1_3;
  wire modExp_while_and_3;
  wire modExp_while_and_5;
  wire and_345_m1c;
  wire modExp_result_and_rgt;
  wire modExp_result_and_1_rgt;
  wire COMP_LOOP_or_32_cse;
  wire nor_1148_cse;
  wire or_642_cse;
  wire nor_1123_cse;
  wire or_748_cse;
  wire nor_1098_cse;
  wire or_855_cse;
  wire nor_1073_cse;
  wire or_961_cse;
  wire nor_1048_cse;
  wire or_1068_cse;
  wire nor_1023_cse;
  wire or_1174_cse;
  wire nor_998_cse;
  wire or_1281_cse;
  wire nor_975_cse;
  wire or_1387_cse;
  wire nor_950_cse;
  wire or_1494_cse;
  wire nor_925_cse;
  wire or_1600_cse;
  wire nor_900_cse;
  wire or_1707_cse;
  wire nor_877_cse;
  wire or_1813_cse;
  wire nor_850_cse;
  wire or_1923_cse;
  wire nor_827_cse;
  wire or_2029_cse;
  wire nor_804_cse;
  wire or_2136_cse;
  wire and_591_cse;
  wire nand_278_cse;
  wire nand_257_cse;
  wire nor_738_cse;
  wire COMP_LOOP_or_55_ssc;
  wire COMP_LOOP_or_56_ssc;
  wire COMP_LOOP_or_57_ssc;
  wire COMP_LOOP_or_58_ssc;
  wire and_850_cse;
  wire and_857_cse;
  wire and_869_cse;
  wire and_875_cse;
  wire and_886_cse;
  wire or_tmp;
  wire nor_tmp;
  wire mux_tmp_3818;
  wire not_tmp_1007;
  wire mux_tmp_3819;
  wire mux_tmp_3822;
  wire or_tmp_3291;
  wire or_tmp_3293;
  wire nor_tmp_535;
  wire nor_tmp_536;
  wire mux_tmp_3828;
  wire mux_tmp_3834;
  wire nor_tmp_539;
  wire nor_tmp_540;
  wire or_tmp_3303;
  wire or_tmp_3304;
  wire mux_tmp_3846;
  wire mux_tmp_3853;
  wire not_tmp_1021;
  wire mux_tmp_3861;
  wire mux_tmp_3878;
  wire or_tmp_3320;
  wire not_tmp_1034;
  wire or_tmp_3327;
  wire mux_tmp_3898;
  wire or_tmp_3332;
  wire nand_tmp;
  wire mux_tmp_3902;
  wire mux_tmp_3906;
  wire or_tmp_3343;
  wire mux_tmp_3915;
  wire or_tmp_3369;
  wire [64:0] operator_64_false_mux1h_2_rgt;
  reg operator_64_false_acc_mut_64;
  reg [63:0] operator_64_false_acc_mut_63_0;
  wire and_1262_cse;
  wire nor_1450_cse;
  wire or_2747_cse;
  wire nand_201_cse;
  wire or_2415_cse;
  wire or_3280_cse;
  wire mux_3724_itm;
  wire mux_3788_itm;
  wire COMP_LOOP_or_60_itm;
  wire COMP_LOOP_or_24_itm;
  wire COMP_LOOP_or_67_itm;
  wire COMP_LOOP_nor_680_itm;
  wire STAGE_LOOP_acc_itm_2_1;
  wire COMP_LOOP_COMP_LOOP_or_6_cse;
  wire COMP_LOOP_COMP_LOOP_or_9_cse;
  wire [1:0] z_out_8_8_7;

  wire[0:0] mux_1092_nl;
  wire[0:0] nand_360_nl;
  wire[0:0] or_619_nl;
  wire[0:0] modulo_result_or_nl;
  wire[0:0] mux_2303_nl;
  wire[0:0] mux_2302_nl;
  wire[0:0] mux_2301_nl;
  wire[0:0] mux_2300_nl;
  wire[0:0] mux_2299_nl;
  wire[0:0] mux_2298_nl;
  wire[0:0] mux_2297_nl;
  wire[0:0] mux_2296_nl;
  wire[0:0] mux_2295_nl;
  wire[0:0] mux_2294_nl;
  wire[0:0] mux_2293_nl;
  wire[0:0] mux_2292_nl;
  wire[0:0] mux_2291_nl;
  wire[0:0] nand_264_nl;
  wire[0:0] mux_2288_nl;
  wire[0:0] mux_2287_nl;
  wire[0:0] mux_2286_nl;
  wire[0:0] mux_2284_nl;
  wire[0:0] mux_2283_nl;
  wire[0:0] mux_2282_nl;
  wire[0:0] mux_2281_nl;
  wire[0:0] mux_2280_nl;
  wire[0:0] mux_2278_nl;
  wire[0:0] mux_2277_nl;
  wire[0:0] nand_265_nl;
  wire[0:0] mux_2276_nl;
  wire[0:0] mux_2275_nl;
  wire[0:0] mux_2274_nl;
  wire[0:0] mux_2273_nl;
  wire[0:0] mux_2272_nl;
  wire[0:0] mux_2271_nl;
  wire[0:0] mux_2270_nl;
  wire[0:0] mux_2269_nl;
  wire[0:0] mux_2268_nl;
  wire[0:0] mux_2267_nl;
  wire[0:0] mux_2266_nl;
  wire[0:0] mux_2264_nl;
  wire[0:0] mux_2263_nl;
  wire[0:0] mux_2262_nl;
  wire[0:0] nor_778_nl;
  wire[0:0] mux_2261_nl;
  wire[0:0] mux_2260_nl;
  wire[0:0] mux_2259_nl;
  wire[0:0] mux_2258_nl;
  wire[0:0] mux_2257_nl;
  wire[0:0] mux_2256_nl;
  wire[0:0] nor_779_nl;
  wire[0:0] mux_2255_nl;
  wire[0:0] mux_2253_nl;
  wire[0:0] mux_2252_nl;
  wire[0:0] mux_2249_nl;
  wire[0:0] mux_2248_nl;
  wire[0:0] mux_2247_nl;
  wire[0:0] mux_2246_nl;
  wire[0:0] or_2306_nl;
  wire[0:0] mux_2245_nl;
  wire[0:0] mux_2244_nl;
  wire[0:0] mux_2243_nl;
  wire[0:0] mux_2242_nl;
  wire[0:0] mux_2241_nl;
  wire[0:0] mux_2238_nl;
  wire[0:0] mux_2237_nl;
  wire[0:0] mux_2236_nl;
  wire[0:0] mux_2235_nl;
  wire[0:0] or_2300_nl;
  wire[0:0] nand_91_nl;
  wire[0:0] mux_2234_nl;
  wire[0:0] or_2297_nl;
  wire[0:0] mux_2233_nl;
  wire[0:0] mux_2232_nl;
  wire[0:0] or_2293_nl;
  wire[0:0] mux_2231_nl;
  wire[0:0] mux_2230_nl;
  wire[0:0] mux_2229_nl;
  wire[0:0] mux_2228_nl;
  wire[0:0] mux_2227_nl;
  wire[0:0] mux_2226_nl;
  wire[0:0] mux_2225_nl;
  wire[0:0] mux_2224_nl;
  wire[0:0] mux_2222_nl;
  wire[0:0] mux_2221_nl;
  wire[0:0] mux_2219_nl;
  wire[0:0] or_2288_nl;
  wire[0:0] mux_2217_nl;
  wire[0:0] mux_2216_nl;
  wire[0:0] mux_2215_nl;
  wire[0:0] or_2285_nl;
  wire[0:0] or_2283_nl;
  wire[0:0] mux_2214_nl;
  wire[0:0] mux_2213_nl;
  wire[0:0] mux_2212_nl;
  wire[0:0] or_2279_nl;
  wire[0:0] mux_2211_nl;
  wire[0:0] nand_90_nl;
  wire[0:0] mux_2378_nl;
  wire[0:0] mux_2377_nl;
  wire[0:0] mux_2376_nl;
  wire[0:0] mux_2375_nl;
  wire[0:0] mux_2374_nl;
  wire[0:0] mux_2373_nl;
  wire[0:0] or_2355_nl;
  wire[0:0] mux_2372_nl;
  wire[0:0] mux_2371_nl;
  wire[0:0] mux_2370_nl;
  wire[0:0] mux_2369_nl;
  wire[0:0] or_2354_nl;
  wire[0:0] mux_2368_nl;
  wire[0:0] or_2351_nl;
  wire[0:0] mux_2367_nl;
  wire[0:0] mux_2366_nl;
  wire[0:0] mux_2365_nl;
  wire[0:0] mux_2364_nl;
  wire[0:0] mux_2363_nl;
  wire[0:0] nand_100_nl;
  wire[0:0] mux_2361_nl;
  wire[0:0] mux_2360_nl;
  wire[0:0] nand_99_nl;
  wire[0:0] mux_2359_nl;
  wire[0:0] nand_98_nl;
  wire[0:0] mux_2358_nl;
  wire[0:0] mux_2357_nl;
  wire[0:0] mux_2356_nl;
  wire[0:0] mux_2355_nl;
  wire[0:0] mux_2354_nl;
  wire[0:0] mux_2353_nl;
  wire[0:0] mux_2352_nl;
  wire[0:0] mux_2351_nl;
  wire[0:0] mux_2350_nl;
  wire[0:0] mux_2348_nl;
  wire[0:0] nand_261_nl;
  wire[0:0] mux_2347_nl;
  wire[0:0] and_275_nl;
  wire[0:0] mux_2346_nl;
  wire[0:0] mux_2345_nl;
  wire[0:0] mux_2344_nl;
  wire[0:0] mux_2343_nl;
  wire[0:0] or_2343_nl;
  wire[0:0] mux_2342_nl;
  wire[0:0] or_2342_nl;
  wire[0:0] mux_2341_nl;
  wire[0:0] mux_2340_nl;
  wire[0:0] nand_262_nl;
  wire[0:0] mux_2339_nl;
  wire[0:0] or_2341_nl;
  wire[0:0] mux_2338_nl;
  wire[0:0] mux_2337_nl;
  wire[0:0] mux_2336_nl;
  wire[0:0] mux_2335_nl;
  wire[0:0] mux_2334_nl;
  wire[0:0] mux_2333_nl;
  wire[0:0] mux_2332_nl;
  wire[0:0] mux_2331_nl;
  wire[0:0] mux_2330_nl;
  wire[0:0] mux_2329_nl;
  wire[0:0] mux_2328_nl;
  wire[0:0] mux_2326_nl;
  wire[0:0] mux_2325_nl;
  wire[0:0] mux_2324_nl;
  wire[0:0] mux_2323_nl;
  wire[0:0] nand_97_nl;
  wire[0:0] mux_2322_nl;
  wire[0:0] mux_2321_nl;
  wire[0:0] mux_2320_nl;
  wire[0:0] mux_2319_nl;
  wire[0:0] mux_2318_nl;
  wire[0:0] mux_2317_nl;
  wire[0:0] mux_2316_nl;
  wire[0:0] mux_2315_nl;
  wire[0:0] mux_2314_nl;
  wire[0:0] or_2330_nl;
  wire[0:0] or_2329_nl;
  wire[0:0] mux_2313_nl;
  wire[0:0] mux_2312_nl;
  wire[0:0] mux_2311_nl;
  wire[0:0] mux_2308_nl;
  wire[0:0] nand_94_nl;
  wire[0:0] mux_2307_nl;
  wire[0:0] mux_2306_nl;
  wire[0:0] mux_2305_nl;
  wire[0:0] or_2321_nl;
  wire[0:0] mux_2304_nl;
  wire[0:0] or_2319_nl;
  wire[0:0] mux_2394_nl;
  wire[0:0] mux_2393_nl;
  wire[0:0] mux_2392_nl;
  wire[0:0] mux_2391_nl;
  wire[0:0] nor_758_nl;
  wire[0:0] nor_759_nl;
  wire[0:0] and_568_nl;
  wire[0:0] mux_2390_nl;
  wire[0:0] nor_760_nl;
  wire[0:0] nor_761_nl;
  wire[0:0] mux_2389_nl;
  wire[0:0] mux_2388_nl;
  wire[0:0] nor_762_nl;
  wire[0:0] nor_763_nl;
  wire[0:0] nor_764_nl;
  wire[0:0] mux_2387_nl;
  wire[0:0] or_2372_nl;
  wire[0:0] or_2370_nl;
  wire[0:0] mux_2386_nl;
  wire[0:0] and_569_nl;
  wire[0:0] mux_2385_nl;
  wire[0:0] and_570_nl;
  wire[0:0] mux_2384_nl;
  wire[0:0] nor_765_nl;
  wire[0:0] nor_766_nl;
  wire[0:0] nor_767_nl;
  wire[0:0] mux_2383_nl;
  wire[0:0] or_2365_nl;
  wire[0:0] or_2364_nl;
  wire[0:0] mux_2382_nl;
  wire[0:0] mux_2381_nl;
  wire[0:0] nor_768_nl;
  wire[0:0] mux_2380_nl;
  wire[0:0] mux_2379_nl;
  wire[0:0] nor_769_nl;
  wire[0:0] nor_770_nl;
  wire[0:0] nor_771_nl;
  wire[0:0] nor_772_nl;
  wire[0:0] mux_2461_nl;
  wire[0:0] mux_2460_nl;
  wire[0:0] mux_2459_nl;
  wire[0:0] mux_2458_nl;
  wire[0:0] mux_2457_nl;
  wire[0:0] mux_2456_nl;
  wire[0:0] nand_109_nl;
  wire[0:0] mux_2455_nl;
  wire[0:0] mux_2454_nl;
  wire[0:0] mux_2453_nl;
  wire[0:0] mux_2452_nl;
  wire[0:0] mux_2451_nl;
  wire[0:0] mux_2450_nl;
  wire[0:0] mux_2449_nl;
  wire[0:0] mux_2448_nl;
  wire[0:0] mux_2447_nl;
  wire[0:0] mux_2446_nl;
  wire[0:0] mux_2445_nl;
  wire[0:0] mux_2444_nl;
  wire[0:0] mux_2443_nl;
  wire[0:0] mux_2442_nl;
  wire[0:0] mux_2441_nl;
  wire[0:0] mux_2440_nl;
  wire[0:0] mux_2439_nl;
  wire[0:0] mux_2438_nl;
  wire[0:0] mux_2437_nl;
  wire[0:0] mux_2434_nl;
  wire[0:0] mux_2432_nl;
  wire[0:0] mux_2431_nl;
  wire[0:0] mux_2430_nl;
  wire[0:0] mux_2429_nl;
  wire[0:0] mux_2428_nl;
  wire[0:0] mux_2424_nl;
  wire[0:0] nand_106_nl;
  wire[0:0] mux_2421_nl;
  wire[0:0] mux_2420_nl;
  wire[0:0] mux_2419_nl;
  wire[0:0] mux_2418_nl;
  wire[0:0] mux_2417_nl;
  wire[0:0] mux_2416_nl;
  wire[0:0] or_2397_nl;
  wire[0:0] mux_2415_nl;
  wire[0:0] mux_2414_nl;
  wire[0:0] mux_2413_nl;
  wire[0:0] mux_2412_nl;
  wire[0:0] mux_2411_nl;
  wire[0:0] mux_2410_nl;
  wire[0:0] mux_2409_nl;
  wire[0:0] mux_2408_nl;
  wire[0:0] mux_2407_nl;
  wire[0:0] mux_2405_nl;
  wire[0:0] mux_2404_nl;
  wire[0:0] mux_2403_nl;
  wire[0:0] mux_2399_nl;
  wire[0:0] mux_2398_nl;
  wire[0:0] mux_2397_nl;
  wire[0:0] mux_2396_nl;
  wire[0:0] nand_104_nl;
  wire[0:0] mux_2395_nl;
  wire[0:0] or_2381_nl;
  wire[0:0] mux_2495_nl;
  wire[0:0] mux_2494_nl;
  wire[0:0] mux_2493_nl;
  wire[0:0] or_3297_nl;
  wire[0:0] nand_250_nl;
  wire[0:0] or_2778_nl;
  wire[63:0] modExp_while_if_mux1h_nl;
  wire[0:0] and_353_nl;
  wire[0:0] mux_3149_nl;
  wire[0:0] mux_3148_nl;
  wire[0:0] mux_3147_nl;
  wire[0:0] mux_3146_nl;
  wire[0:0] and_466_nl;
  wire[0:0] mux_3145_nl;
  wire[0:0] nor_637_nl;
  wire[0:0] nor_638_nl;
  wire[0:0] nor_639_nl;
  wire[0:0] and_467_nl;
  wire[0:0] and_468_nl;
  wire[0:0] mux_3144_nl;
  wire[0:0] nor_640_nl;
  wire[0:0] nor_641_nl;
  wire[0:0] mux_3142_nl;
  wire[0:0] mux_3141_nl;
  wire[0:0] mux_3140_nl;
  wire[0:0] nor_642_nl;
  wire[0:0] and_469_nl;
  wire[0:0] nor_643_nl;
  wire[0:0] mux_3139_nl;
  wire[0:0] mux_3138_nl;
  wire[0:0] or_2773_nl;
  wire[0:0] or_2772_nl;
  wire[0:0] or_2771_nl;
  wire[0:0] mux_3137_nl;
  wire[0:0] or_2770_nl;
  wire[0:0] and_470_nl;
  wire[0:0] mux_3136_nl;
  wire[0:0] nor_644_nl;
  wire[0:0] mux_3135_nl;
  wire[0:0] nor_645_nl;
  wire[0:0] modExp_while_if_and_nl;
  wire[0:0] modExp_while_if_and_1_nl;
  wire[0:0] and_284_nl;
  wire[0:0] mux_2566_nl;
  wire[0:0] mux_2565_nl;
  wire[0:0] mux_2564_nl;
  wire[0:0] mux_2563_nl;
  wire[0:0] mux_2562_nl;
  wire[0:0] mux_2561_nl;
  wire[0:0] mux_2560_nl;
  wire[0:0] mux_2559_nl;
  wire[0:0] mux_2558_nl;
  wire[0:0] and_532_nl;
  wire[0:0] and_533_nl;
  wire[0:0] mux_2557_nl;
  wire[0:0] or_2494_nl;
  wire[0:0] mux_2556_nl;
  wire[0:0] mux_2555_nl;
  wire[0:0] mux_2554_nl;
  wire[0:0] mux_2553_nl;
  wire[0:0] and_535_nl;
  wire[0:0] or_2491_nl;
  wire[0:0] mux_2552_nl;
  wire[0:0] mux_2551_nl;
  wire[0:0] mux_2550_nl;
  wire[0:0] mux_2548_nl;
  wire[0:0] nor_731_nl;
  wire[0:0] mux_2547_nl;
  wire[0:0] mux_2546_nl;
  wire[0:0] mux_2545_nl;
  wire[0:0] mux_2544_nl;
  wire[0:0] mux_2543_nl;
  wire[0:0] mux_2542_nl;
  wire[0:0] mux_2541_nl;
  wire[0:0] or_2484_nl;
  wire[0:0] mux_2540_nl;
  wire[0:0] mux_2539_nl;
  wire[0:0] mux_2538_nl;
  wire[0:0] or_2483_nl;
  wire[0:0] mux_2537_nl;
  wire[0:0] mux_2536_nl;
  wire[0:0] mux_2535_nl;
  wire[0:0] nor_732_nl;
  wire[0:0] mux_2534_nl;
  wire[0:0] or_2480_nl;
  wire[0:0] mux_2533_nl;
  wire[0:0] mux_2532_nl;
  wire[0:0] mux_2531_nl;
  wire[0:0] mux_2530_nl;
  wire[0:0] mux_2529_nl;
  wire[0:0] mux_2528_nl;
  wire[0:0] mux_2527_nl;
  wire[0:0] mux_2526_nl;
  wire[0:0] mux_2524_nl;
  wire[0:0] mux_2522_nl;
  wire[0:0] mux_2521_nl;
  wire[0:0] nor_733_nl;
  wire[0:0] mux_2520_nl;
  wire[0:0] mux_2518_nl;
  wire[0:0] mux_2517_nl;
  wire[0:0] mux_2516_nl;
  wire[0:0] mux_2515_nl;
  wire[0:0] or_2475_nl;
  wire[0:0] mux_2514_nl;
  wire[0:0] mux_2513_nl;
  wire[0:0] or_2472_nl;
  wire[0:0] mux_2512_nl;
  wire[0:0] mux_2511_nl;
  wire[0:0] mux_2510_nl;
  wire[0:0] mux_2509_nl;
  wire[0:0] mux_2507_nl;
  wire[0:0] or_2466_nl;
  wire[0:0] mux_2506_nl;
  wire[0:0] mux_2505_nl;
  wire[0:0] mux_2504_nl;
  wire[0:0] mux_2503_nl;
  wire[0:0] or_2460_nl;
  wire[0:0] mux_2500_nl;
  wire[0:0] and_544_nl;
  wire[0:0] mux_2499_nl;
  wire[0:0] mux_2498_nl;
  wire[0:0] nand_247_nl;
  wire[0:0] mux_2497_nl;
  wire[0:0] nand_248_nl;
  wire[0:0] or_2454_nl;
  wire[0:0] mux_3896_nl;
  wire[0:0] mux_3895_nl;
  wire[0:0] mux_3894_nl;
  wire[0:0] mux_3893_nl;
  wire[0:0] mux_3892_nl;
  wire[0:0] mux_3891_nl;
  wire[0:0] mux_3890_nl;
  wire[0:0] nor_1453_nl;
  wire[0:0] mux_3889_nl;
  wire[0:0] mux_3888_nl;
  wire[0:0] mux_3887_nl;
  wire[0:0] and_1258_nl;
  wire[0:0] mux_3886_nl;
  wire[0:0] or_3508_nl;
  wire[0:0] mux_3885_nl;
  wire[0:0] mux_3884_nl;
  wire[0:0] and_1259_nl;
  wire[0:0] mux_3883_nl;
  wire[0:0] mux_3882_nl;
  wire[0:0] mux_3881_nl;
  wire[0:0] and_1260_nl;
  wire[0:0] mux_3880_nl;
  wire[0:0] or_3506_nl;
  wire[0:0] mux_3878_nl;
  wire[0:0] mux_3877_nl;
  wire[0:0] mux_3876_nl;
  wire[0:0] mux_3875_nl;
  wire[0:0] or_3505_nl;
  wire[0:0] mux_3874_nl;
  wire[0:0] or_3504_nl;
  wire[0:0] mux_3873_nl;
  wire[0:0] and_1256_nl;
  wire[0:0] mux_3872_nl;
  wire[0:0] or_3502_nl;
  wire[0:0] mux_3871_nl;
  wire[0:0] mux_3870_nl;
  wire[0:0] mux_3869_nl;
  wire[0:0] mux_3868_nl;
  wire[0:0] mux_3867_nl;
  wire[0:0] mux_3866_nl;
  wire[0:0] mux_3865_nl;
  wire[0:0] mux_3864_nl;
  wire[0:0] mux_3863_nl;
  wire[0:0] mux_3861_nl;
  wire[0:0] or_3500_nl;
  wire[0:0] mux_3860_nl;
  wire[0:0] mux_3859_nl;
  wire[0:0] mux_3858_nl;
  wire[0:0] mux_3857_nl;
  wire[0:0] mux_3856_nl;
  wire[0:0] and_1255_nl;
  wire[0:0] mux_3855_nl;
  wire[0:0] mux_3853_nl;
  wire[0:0] mux_3852_nl;
  wire[0:0] mux_3851_nl;
  wire[0:0] nor_1456_nl;
  wire[0:0] mux_3850_nl;
  wire[0:0] mux_3849_nl;
  wire[0:0] mux_3848_nl;
  wire[0:0] and_1264_nl;
  wire[0:0] mux_3846_nl;
  wire[0:0] mux_3845_nl;
  wire[0:0] mux_3844_nl;
  wire[0:0] mux_3843_nl;
  wire[0:0] mux_3842_nl;
  wire[0:0] or_3493_nl;
  wire[0:0] mux_3841_nl;
  wire[0:0] nor_1457_nl;
  wire[0:0] mux_3840_nl;
  wire[0:0] or_3490_nl;
  wire[0:0] mux_3839_nl;
  wire[0:0] mux_3838_nl;
  wire[0:0] mux_3837_nl;
  wire[0:0] mux_3836_nl;
  wire[0:0] mux_3834_nl;
  wire[0:0] mux_3833_nl;
  wire[0:0] nor_1458_nl;
  wire[0:0] mux_3832_nl;
  wire[0:0] mux_3831_nl;
  wire[0:0] mux_3830_nl;
  wire[0:0] mux_3828_nl;
  wire[0:0] mux_3827_nl;
  wire[0:0] mux_3826_nl;
  wire[0:0] nor_1459_nl;
  wire[0:0] mux_3825_nl;
  wire[0:0] mux_3824_nl;
  wire[0:0] mux_3822_nl;
  wire[0:0] or_3480_nl;
  wire[0:0] mux_3821_nl;
  wire[0:0] mux_3949_nl;
  wire[0:0] mux_3948_nl;
  wire[0:0] mux_3947_nl;
  wire[0:0] mux_3946_nl;
  wire[0:0] mux_3945_nl;
  wire[0:0] or_3579_nl;
  wire[0:0] mux_3944_nl;
  wire[0:0] nand_463_nl;
  wire[0:0] mux_3943_nl;
  wire[0:0] mux_3942_nl;
  wire[0:0] or_3577_nl;
  wire[0:0] mux_3941_nl;
  wire[0:0] mux_3940_nl;
  wire[0:0] mux_3939_nl;
  wire[0:0] nand_462_nl;
  wire[0:0] mux_3938_nl;
  wire[0:0] nor_1448_nl;
  wire[0:0] nor_1449_nl;
  wire[0:0] or_3574_nl;
  wire[0:0] or_3572_nl;
  wire[0:0] mux_3937_nl;
  wire[0:0] mux_3936_nl;
  wire[0:0] mux_3935_nl;
  wire[0:0] or_3568_nl;
  wire[0:0] mux_3934_nl;
  wire[0:0] or_3567_nl;
  wire[0:0] or_3565_nl;
  wire[0:0] mux_3933_nl;
  wire[0:0] mux_3932_nl;
  wire[0:0] nand_461_nl;
  wire[0:0] mux_3931_nl;
  wire[0:0] or_3559_nl;
  wire[0:0] mux_3930_nl;
  wire[0:0] nand_465_nl;
  wire[0:0] mux_3929_nl;
  wire[0:0] or_3556_nl;
  wire[0:0] mux_3928_nl;
  wire[0:0] mux_3927_nl;
  wire[0:0] mux_3926_nl;
  wire[0:0] mux_3925_nl;
  wire[0:0] mux_3924_nl;
  wire[0:0] mux_3923_nl;
  wire[0:0] mux_3922_nl;
  wire[0:0] or_3554_nl;
  wire[0:0] nand_471_nl;
  wire[0:0] mux_3921_nl;
  wire[0:0] or_3551_nl;
  wire[0:0] or_3550_nl;
  wire[0:0] mux_3920_nl;
  wire[0:0] mux_3919_nl;
  wire[0:0] nand_460_nl;
  wire[0:0] mux_3918_nl;
  wire[0:0] mux_3917_nl;
  wire[0:0] or_3548_nl;
  wire[0:0] or_3547_nl;
  wire[0:0] mux_3915_nl;
  wire[0:0] or_3546_nl;
  wire[0:0] mux_3914_nl;
  wire[0:0] or_3544_nl;
  wire[0:0] mux_3913_nl;
  wire[0:0] mux_3912_nl;
  wire[0:0] or_3542_nl;
  wire[0:0] or_3540_nl;
  wire[0:0] nand_459_nl;
  wire[0:0] mux_3911_nl;
  wire[0:0] or_3536_nl;
  wire[0:0] mux_3910_nl;
  wire[0:0] or_3534_nl;
  wire[0:0] mux_3909_nl;
  wire[0:0] or_3533_nl;
  wire[0:0] or_3532_nl;
  wire[0:0] mux_3908_nl;
  wire[0:0] or_3527_nl;
  wire[0:0] mux_3905_nl;
  wire[0:0] mux_3904_nl;
  wire[0:0] or_3589_nl;
  wire[0:0] mux_3901_nl;
  wire[0:0] mux_3900_nl;
  wire[0:0] or_3521_nl;
  wire[0:0] mux_3897_nl;
  wire[0:0] or_3514_nl;
  wire[0:0] or_3477_nl;
  wire[0:0] mux_2649_nl;
  wire[0:0] mux_2648_nl;
  wire[0:0] or_2515_nl;
  wire[0:0] or_2514_nl;
  wire[0:0] or_2513_nl;
  wire[0:0] mux_3952_nl;
  wire[0:0] or_3587_nl;
  wire[0:0] mux_3951_nl;
  wire[0:0] or_3585_nl;
  wire[0:0] mux_3950_nl;
  wire[0:0] or_3584_nl;
  wire[0:0] or_3583_nl;
  wire[0:0] or_3581_nl;
  wire[0:0] or_3588_nl;
  wire[0:0] mux_2675_nl;
  wire[0:0] mux_2674_nl;
  wire[0:0] mux_2673_nl;
  wire[0:0] mux_2672_nl;
  wire[0:0] mux_2671_nl;
  wire[0:0] mux_2670_nl;
  wire[0:0] nor_725_nl;
  wire[0:0] mux_2669_nl;
  wire[0:0] mux_2668_nl;
  wire[0:0] mux_2667_nl;
  wire[0:0] nand_244_nl;
  wire[0:0] or_4_nl;
  wire[0:0] COMP_LOOP_or_8_nl;
  wire[0:0] COMP_LOOP_or_9_nl;
  wire[0:0] COMP_LOOP_or_10_nl;
  wire[0:0] COMP_LOOP_or_11_nl;
  wire[0:0] COMP_LOOP_or_12_nl;
  wire[0:0] COMP_LOOP_or_13_nl;
  wire[0:0] COMP_LOOP_or_14_nl;
  wire[0:0] COMP_LOOP_or_15_nl;
  wire[0:0] COMP_LOOP_or_16_nl;
  wire[0:0] COMP_LOOP_or_17_nl;
  wire[0:0] COMP_LOOP_or_18_nl;
  wire[0:0] COMP_LOOP_or_19_nl;
  wire[0:0] COMP_LOOP_or_20_nl;
  wire[0:0] COMP_LOOP_or_21_nl;
  wire[0:0] COMP_LOOP_or_22_nl;
  wire[0:0] COMP_LOOP_or_23_nl;
  wire[0:0] mux_2740_nl;
  wire[0:0] mux_2739_nl;
  wire[0:0] mux_2738_nl;
  wire[0:0] mux_2737_nl;
  wire[0:0] mux_2736_nl;
  wire[0:0] nor_716_nl;
  wire[0:0] mux_2735_nl;
  wire[0:0] mux_2734_nl;
  wire[0:0] mux_2733_nl;
  wire[0:0] mux_2732_nl;
  wire[0:0] or_3268_nl;
  wire[0:0] mux_2731_nl;
  wire[0:0] mux_2730_nl;
  wire[0:0] mux_2729_nl;
  wire[0:0] mux_2728_nl;
  wire[0:0] mux_2727_nl;
  wire[0:0] mux_55_nl;
  wire[0:0] mux_2725_nl;
  wire[0:0] mux_2724_nl;
  wire[0:0] mux_2723_nl;
  wire[0:0] mux_2722_nl;
  wire[0:0] mux_50_nl;
  wire[0:0] mux_2720_nl;
  wire[0:0] mux_2719_nl;
  wire[0:0] mux_2718_nl;
  wire[0:0] mux_2717_nl;
  wire[0:0] mux_2716_nl;
  wire[0:0] mux_2715_nl;
  wire[0:0] mux_2714_nl;
  wire[0:0] mux_2713_nl;
  wire[0:0] mux_2712_nl;
  wire[0:0] nand_118_nl;
  wire[0:0] mux_2711_nl;
  wire[0:0] or_3269_nl;
  wire[0:0] mux_2710_nl;
  wire[0:0] mux_2709_nl;
  wire[0:0] mux_2708_nl;
  wire[0:0] or_2540_nl;
  wire[0:0] mux_2707_nl;
  wire[0:0] mux_2706_nl;
  wire[0:0] mux_2705_nl;
  wire[0:0] mux_2704_nl;
  wire[0:0] mux_2703_nl;
  wire[0:0] mux_2702_nl;
  wire[0:0] mux_29_nl;
  wire[0:0] mux_2699_nl;
  wire[0:0] mux_2697_nl;
  wire[0:0] mux_22_nl;
  wire[0:0] or_25_nl;
  wire[0:0] or_24_nl;
  wire[0:0] mux_2694_nl;
  wire[0:0] mux_2693_nl;
  wire[0:0] mux_2692_nl;
  wire[0:0] mux_2691_nl;
  wire[0:0] nand_116_nl;
  wire[0:0] mux_17_nl;
  wire[0:0] mux_2689_nl;
  wire[0:0] mux_2688_nl;
  wire[0:0] mux_13_nl;
  wire[0:0] or_18_nl;
  wire[0:0] mux_2685_nl;
  wire[0:0] mux_11_nl;
  wire[0:0] mux_10_nl;
  wire[0:0] mux_8_nl;
  wire[0:0] mux_2679_nl;
  wire[0:0] mux_2678_nl;
  wire[0:0] mux_2677_nl;
  wire[0:0] mux_2769_nl;
  wire[0:0] nor_694_nl;
  wire[0:0] mux_2768_nl;
  wire[0:0] or_2591_nl;
  wire[0:0] or_2589_nl;
  wire[0:0] mux_2767_nl;
  wire[0:0] or_2588_nl;
  wire[0:0] and_513_nl;
  wire[0:0] mux_2766_nl;
  wire[0:0] nor_695_nl;
  wire[0:0] nor_696_nl;
  wire[0:0] mux_2764_nl;
  wire[0:0] and_514_nl;
  wire[0:0] mux_2763_nl;
  wire[0:0] nor_697_nl;
  wire[0:0] nor_698_nl;
  wire[0:0] mux_2762_nl;
  wire[0:0] or_2581_nl;
  wire[0:0] or_2579_nl;
  wire[0:0] mux_2761_nl;
  wire[0:0] mux_2760_nl;
  wire[0:0] mux_2759_nl;
  wire[0:0] and_515_nl;
  wire[0:0] nor_699_nl;
  wire[0:0] nor_700_nl;
  wire[0:0] nor_701_nl;
  wire[0:0] nor_1302_nl;
  wire[0:0] and_801_nl;
  wire[0:0] mux_2742_nl;
  wire[0:0] nor_715_nl;
  wire[0:0] and_340_nl;
  wire[0:0] COMP_LOOP_or_30_nl;
  wire[0:0] COMP_LOOP_or_31_nl;
  wire[0:0] COMP_LOOP_and_277_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_932_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_934_nl;
  wire[0:0] COMP_LOOP_and_1_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_936_nl;
  wire[0:0] COMP_LOOP_and_2_nl;
  wire[0:0] COMP_LOOP_and_3_nl;
  wire[0:0] COMP_LOOP_and_4_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_930_nl;
  wire[0:0] COMP_LOOP_and_5_nl;
  wire[0:0] COMP_LOOP_and_6_nl;
  wire[0:0] COMP_LOOP_and_7_nl;
  wire[0:0] COMP_LOOP_and_8_nl;
  wire[0:0] COMP_LOOP_and_9_nl;
  wire[0:0] COMP_LOOP_and_10_nl;
  wire[0:0] COMP_LOOP_and_11_nl;
  wire[0:0] mux_114_nl;
  wire[0:0] mux_113_nl;
  wire[0:0] mux_112_nl;
  wire[0:0] nor_1265_nl;
  wire[0:0] nor_1266_nl;
  wire[0:0] mux_111_nl;
  wire[0:0] nor_1267_nl;
  wire[0:0] mux_110_nl;
  wire[0:0] or_113_nl;
  wire[0:0] nand_395_nl;
  wire[0:0] mux_109_nl;
  wire[0:0] nor_1268_nl;
  wire[0:0] mux_108_nl;
  wire[0:0] nor_1269_nl;
  wire[0:0] mux_107_nl;
  wire[0:0] or_109_nl;
  wire[0:0] or_108_nl;
  wire[0:0] nor_1270_nl;
  wire[0:0] mux_106_nl;
  wire[0:0] mux_105_nl;
  wire[0:0] mux_104_nl;
  wire[0:0] nor_1271_nl;
  wire[0:0] nor_1272_nl;
  wire[0:0] mux_103_nl;
  wire[0:0] and_794_nl;
  wire[0:0] mux_102_nl;
  wire[0:0] and_795_nl;
  wire[0:0] nor_1273_nl;
  wire[0:0] nor_1274_nl;
  wire[0:0] nor_1275_nl;
  wire[0:0] mux_101_nl;
  wire[0:0] or_98_nl;
  wire[0:0] or_96_nl;
  wire[0:0] mux_100_nl;
  wire[0:0] or_95_nl;
  wire[0:0] or_93_nl;
  wire[0:0] mux_2867_nl;
  wire[0:0] mux_2866_nl;
  wire[0:0] mux_2865_nl;
  wire[0:0] mux_2864_nl;
  wire[0:0] mux_2863_nl;
  wire[0:0] mux_2862_nl;
  wire[0:0] nor_1303_nl;
  wire[0:0] mux_2861_nl;
  wire[0:0] mux_2860_nl;
  wire[0:0] mux_2859_nl;
  wire[0:0] and_506_nl;
  wire[0:0] mux_2858_nl;
  wire[0:0] and_508_nl;
  wire[0:0] mux_2857_nl;
  wire[0:0] mux_2856_nl;
  wire[0:0] or_2643_nl;
  wire[0:0] mux_2855_nl;
  wire[0:0] mux_2854_nl;
  wire[0:0] mux_2853_nl;
  wire[0:0] mux_2852_nl;
  wire[0:0] mux_2851_nl;
  wire[0:0] mux_2850_nl;
  wire[0:0] mux_2849_nl;
  wire[0:0] and_346_nl;
  wire[0:0] mux_2848_nl;
  wire[0:0] mux_2847_nl;
  wire[0:0] mux_2846_nl;
  wire[0:0] mux_2845_nl;
  wire[0:0] mux_2844_nl;
  wire[0:0] mux_2843_nl;
  wire[0:0] mux_2842_nl;
  wire[0:0] mux_2841_nl;
  wire[0:0] mux_2840_nl;
  wire[0:0] mux_2839_nl;
  wire[0:0] or_2639_nl;
  wire[0:0] or_2638_nl;
  wire[0:0] mux_2838_nl;
  wire[0:0] mux_2837_nl;
  wire[0:0] or_2637_nl;
  wire[0:0] mux_2836_nl;
  wire[0:0] mux_2835_nl;
  wire[0:0] or_2636_nl;
  wire[0:0] mux_2834_nl;
  wire[0:0] mux_2833_nl;
  wire[0:0] mux_2832_nl;
  wire[0:0] or_3347_nl;
  wire[0:0] mux_2831_nl;
  wire[0:0] mux_2830_nl;
  wire[0:0] mux_2829_nl;
  wire[0:0] mux_2828_nl;
  wire[0:0] or_2632_nl;
  wire[0:0] mux_2827_nl;
  wire[0:0] mux_2826_nl;
  wire[0:0] mux_2825_nl;
  wire[0:0] mux_2824_nl;
  wire[0:0] mux_2823_nl;
  wire[0:0] mux_2822_nl;
  wire[0:0] mux_2821_nl;
  wire[0:0] mux_2820_nl;
  wire[0:0] mux_2819_nl;
  wire[0:0] mux_2818_nl;
  wire[0:0] nor_680_nl;
  wire[0:0] mux_2817_nl;
  wire[0:0] mux_2816_nl;
  wire[0:0] mux_2815_nl;
  wire[0:0] mux_2814_nl;
  wire[0:0] mux_2812_nl;
  wire[0:0] mux_2811_nl;
  wire[0:0] mux_2810_nl;
  wire[0:0] mux_2809_nl;
  wire[0:0] or_2629_nl;
  wire[0:0] mux_2808_nl;
  wire[0:0] nand_128_nl;
  wire[0:0] mux_2807_nl;
  wire[0:0] mux_2806_nl;
  wire[0:0] mux_2805_nl;
  wire[0:0] mux_2804_nl;
  wire[0:0] mux_2803_nl;
  wire[0:0] mux_2802_nl;
  wire[0:0] mux_2801_nl;
  wire[0:0] nand_127_nl;
  wire[0:0] or_2626_nl;
  wire[0:0] mux_2798_nl;
  wire[0:0] or_2625_nl;
  wire[0:0] or_2624_nl;
  wire[0:0] mux_2797_nl;
  wire[0:0] or_2622_nl;
  wire[0:0] mux_2795_nl;
  wire[0:0] mux_2794_nl;
  wire[0:0] or_2620_nl;
  wire[0:0] mux_2793_nl;
  wire[0:0] mux_2792_nl;
  wire[0:0] mux_2791_nl;
  wire[0:0] mux_2789_nl;
  wire[0:0] nand_126_nl;
  wire[0:0] mux_2787_nl;
  wire[0:0] mux_2786_nl;
  wire[0:0] or_199_nl;
  wire[0:0] COMP_LOOP_mux1h_428_nl;
  wire[0:0] COMP_LOOP_nor_11_nl;
  wire[0:0] COMP_LOOP_and_274_nl;
  wire[0:0] mux_2976_nl;
  wire[0:0] mux_2975_nl;
  wire[0:0] mux_2974_nl;
  wire[0:0] mux_2973_nl;
  wire[0:0] mux_2972_nl;
  wire[0:0] mux_2971_nl;
  wire[0:0] or_2728_nl;
  wire[0:0] mux_2970_nl;
  wire[0:0] mux_2969_nl;
  wire[0:0] mux_2968_nl;
  wire[0:0] mux_2967_nl;
  wire[0:0] mux_2966_nl;
  wire[0:0] mux_2965_nl;
  wire[0:0] mux_2964_nl;
  wire[0:0] mux_2963_nl;
  wire[0:0] mux_2962_nl;
  wire[0:0] mux_2961_nl;
  wire[0:0] mux_2960_nl;
  wire[0:0] mux_427_nl;
  wire[0:0] mux_426_nl;
  wire[0:0] mux_2957_nl;
  wire[0:0] mux_2956_nl;
  wire[0:0] mux_2955_nl;
  wire[0:0] mux_2954_nl;
  wire[0:0] mux_422_nl;
  wire[0:0] mux_421_nl;
  wire[0:0] mux_2951_nl;
  wire[0:0] mux_2950_nl;
  wire[0:0] mux_2949_nl;
  wire[0:0] mux_2948_nl;
  wire[0:0] mux_2947_nl;
  wire[0:0] mux_2946_nl;
  wire[0:0] mux_414_nl;
  wire[0:0] mux_2942_nl;
  wire[0:0] mux_2941_nl;
  wire[0:0] mux_2940_nl;
  wire[0:0] mux_2939_nl;
  wire[0:0] mux_2938_nl;
  wire[0:0] mux_2936_nl;
  wire[0:0] mux_2935_nl;
  wire[0:0] mux_2934_nl;
  wire[0:0] mux_2933_nl;
  wire[0:0] mux_2932_nl;
  wire[0:0] mux_2931_nl;
  wire[0:0] mux_2929_nl;
  wire[0:0] mux_2928_nl;
  wire[0:0] mux_2927_nl;
  wire[0:0] mux_2926_nl;
  wire[0:0] mux_2925_nl;
  wire[0:0] mux_2924_nl;
  wire[0:0] or_2718_nl;
  wire[0:0] mux_2923_nl;
  wire[0:0] mux_2922_nl;
  wire[0:0] mux_2918_nl;
  wire[0:0] mux_386_nl;
  wire[0:0] mux_2916_nl;
  wire[0:0] mux_2914_nl;
  wire[0:0] mux_2909_nl;
  wire[0:0] mux_2908_nl;
  wire[0:0] mux_2888_nl;
  wire[0:0] mux_2887_nl;
  wire[0:0] or_3351_nl;
  wire[0:0] nand_421_nl;
  wire[0:0] mux_2886_nl;
  wire[0:0] nor_667_nl;
  wire[0:0] mux_2885_nl;
  wire[0:0] or_2678_nl;
  wire[0:0] nor_668_nl;
  wire[0:0] mux_2884_nl;
  wire[0:0] or_3352_nl;
  wire[0:0] mux_2883_nl;
  wire[0:0] or_2674_nl;
  wire[0:0] or_2673_nl;
  wire[0:0] nand_422_nl;
  wire[0:0] mux_2882_nl;
  wire[0:0] nor_671_nl;
  wire[0:0] mux_2983_nl;
  wire[0:0] mux_2982_nl;
  wire[0:0] mux_2981_nl;
  wire[0:0] mux_2980_nl;
  wire[0:0] nor_646_nl;
  wire[0:0] nor_647_nl;
  wire[0:0] nor_648_nl;
  wire[0:0] nor_649_nl;
  wire[0:0] mux_2979_nl;
  wire[0:0] nor_650_nl;
  wire[0:0] and_490_nl;
  wire[0:0] mux_2978_nl;
  wire[0:0] mux_2977_nl;
  wire[0:0] nor_651_nl;
  wire[0:0] nor_652_nl;
  wire[0:0] nor_653_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_17_nl;
  wire[63:0] COMP_LOOP_1_acc_8_nl;
  wire[64:0] nl_COMP_LOOP_1_acc_8_nl;
  wire[0:0] mux_3181_nl;
  wire[0:0] mux_3180_nl;
  wire[0:0] nor_620_nl;
  wire[0:0] mux_3179_nl;
  wire[0:0] mux_3178_nl;
  wire[0:0] or_2838_nl;
  wire[0:0] mux_3177_nl;
  wire[0:0] nor_621_nl;
  wire[0:0] mux_3176_nl;
  wire[0:0] mux_3175_nl;
  wire[0:0] nor_622_nl;
  wire[0:0] nor_623_nl;
  wire[0:0] mux_3174_nl;
  wire[0:0] mux_3173_nl;
  wire[0:0] mux_3172_nl;
  wire[0:0] nor_624_nl;
  wire[0:0] nor_625_nl;
  wire[0:0] mux_3171_nl;
  wire[0:0] mux_3170_nl;
  wire[0:0] or_2828_nl;
  wire[0:0] or_2827_nl;
  wire[0:0] and_465_nl;
  wire[0:0] mux_3169_nl;
  wire[0:0] nor_626_nl;
  wire[0:0] mux_3167_nl;
  wire[0:0] or_2817_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_10_nl;
  wire[9:0] COMP_LOOP_1_acc_nl;
  wire[10:0] nl_COMP_LOOP_1_acc_nl;
  wire[0:0] nor_nl;
  wire[0:0] and_1253_nl;
  wire[0:0] mux_3217_nl;
  wire[0:0] mux_3216_nl;
  wire[0:0] or_3259_nl;
  wire[0:0] mux_3215_nl;
  wire[0:0] nor_617_nl;
  wire[0:0] or_2888_nl;
  wire[0:0] mux_3224_nl;
  wire[0:0] mux_3223_nl;
  wire[0:0] mux_3222_nl;
  wire[0:0] mux_3221_nl;
  wire[0:0] mux_3220_nl;
  wire[0:0] and_452_nl;
  wire[0:0] and_454_nl;
  wire[0:0] mux_3234_nl;
  wire[0:0] mux_3233_nl;
  wire[0:0] mux_3232_nl;
  wire[0:0] mux_3231_nl;
  wire[0:0] mux_3230_nl;
  wire[0:0] mux_3229_nl;
  wire[0:0] and_363_nl;
  wire[0:0] mux_3228_nl;
  wire[0:0] mux_3227_nl;
  wire[0:0] mux_3226_nl;
  wire[0:0] nor_729_nl;
  wire[0:0] mux_3225_nl;
  wire[0:0] mux_3242_nl;
  wire[0:0] mux_3241_nl;
  wire[0:0] mux_3240_nl;
  wire[0:0] mux_3239_nl;
  wire[0:0] mux_3238_nl;
  wire[0:0] or_2906_nl;
  wire[0:0] mux_3237_nl;
  wire[0:0] mux_3243_nl;
  wire[0:0] or_3252_nl;
  wire[0:0] nand_218_nl;
  wire[0:0] mux_3249_nl;
  wire[0:0] mux_3248_nl;
  wire[0:0] mux_3247_nl;
  wire[0:0] mux_3246_nl;
  wire[0:0] mux_3245_nl;
  wire[0:0] or_2915_nl;
  wire[0:0] or_2913_nl;
  wire[0:0] mux_3251_nl;
  wire[0:0] mux_3250_nl;
  wire[0:0] nor_1317_nl;
  wire[0:0] or_3346_nl;
  wire[0:0] mux_3255_nl;
  wire[0:0] mux_3254_nl;
  wire[0:0] mux_3253_nl;
  wire[0:0] nor_611_nl;
  wire[0:0] mux_3252_nl;
  wire[0:0] and_371_nl;
  wire[0:0] or_2922_nl;
  wire[0:0] mux_3263_nl;
  wire[0:0] mux_3262_nl;
  wire[0:0] mux_3261_nl;
  wire[0:0] mux_3260_nl;
  wire[0:0] mux_3259_nl;
  wire[0:0] mux_3258_nl;
  wire[0:0] mux_3257_nl;
  wire[0:0] mux_3267_nl;
  wire[0:0] mux_3266_nl;
  wire[0:0] mux_3265_nl;
  wire[0:0] or_2933_nl;
  wire[0:0] mux_3264_nl;
  wire[0:0] or_2930_nl;
  wire[0:0] mux_3276_nl;
  wire[0:0] mux_3275_nl;
  wire[0:0] mux_3274_nl;
  wire[0:0] mux_3273_nl;
  wire[0:0] mux_3272_nl;
  wire[0:0] mux_3271_nl;
  wire[0:0] mux_3270_nl;
  wire[0:0] and_439_nl;
  wire[0:0] mux_3288_nl;
  wire[0:0] mux_3287_nl;
  wire[0:0] mux_3286_nl;
  wire[0:0] mux_3285_nl;
  wire[0:0] and_434_nl;
  wire[0:0] mux_3284_nl;
  wire[0:0] mux_3283_nl;
  wire[0:0] mux_3282_nl;
  wire[0:0] mux_3292_nl;
  wire[0:0] mux_3291_nl;
  wire[0:0] nor_604_nl;
  wire[0:0] mux_3290_nl;
  wire[0:0] nor_605_nl;
  wire[0:0] and_431_nl;
  wire[0:0] and_433_nl;
  wire[0:0] mux_3297_nl;
  wire[0:0] nor_603_nl;
  wire[0:0] mux_3296_nl;
  wire[0:0] or_2947_nl;
  wire[0:0] and_375_nl;
  wire[0:0] mux_3295_nl;
  wire[0:0] and_374_nl;
  wire[0:0] mux_3294_nl;
  wire[0:0] and_430_nl;
  wire[0:0] or_2945_nl;
  wire[0:0] nor_1420_nl;
  wire[0:0] mux_3299_nl;
  wire[0:0] or_2950_nl;
  wire[0:0] and_1254_nl;
  wire[0:0] mux_3304_nl;
  wire[0:0] nor_1201_nl;
  wire[0:0] mux_3303_nl;
  wire[0:0] mux_3302_nl;
  wire[0:0] mux_3301_nl;
  wire[0:0] and_29_nl;
  wire[0:0] mux_3393_nl;
  wire[0:0] or_3014_nl;
  wire[0:0] mux_3384_nl;
  wire[0:0] or_3004_nl;
  wire[0:0] or_3001_nl;
  wire[0:0] nor_581_nl;
  wire[0:0] mux_3391_nl;
  wire[0:0] nor_582_nl;
  wire[0:0] mux_3390_nl;
  wire[0:0] and_414_nl;
  wire[0:0] mux_3389_nl;
  wire[0:0] nor_583_nl;
  wire[0:0] and_415_nl;
  wire[0:0] nor_584_nl;
  wire[0:0] mux_3387_nl;
  wire[0:0] and_416_nl;
  wire[0:0] nor_585_nl;
  wire[0:0] nor_586_nl;
  wire[0:0] COMP_LOOP_mux1h_464_nl;
  wire[0:0] mux_3396_nl;
  wire[0:0] mux_3395_nl;
  wire[0:0] nor_580_nl;
  wire[0:0] or_3241_nl;
  wire[0:0] nand_205_nl;
  wire[0:0] COMP_LOOP_mux1h_474_nl;
  wire[0:0] COMP_LOOP_nor_12_nl;
  wire[0:0] mux_3492_nl;
  wire[0:0] mux_3491_nl;
  wire[0:0] mux_3490_nl;
  wire[0:0] mux_3489_nl;
  wire[0:0] mux_3488_nl;
  wire[0:0] mux_3487_nl;
  wire[0:0] mux_3486_nl;
  wire[0:0] mux_3485_nl;
  wire[0:0] mux_3484_nl;
  wire[0:0] mux_3483_nl;
  wire[0:0] mux_3482_nl;
  wire[0:0] mux_3481_nl;
  wire[0:0] mux_3480_nl;
  wire[0:0] mux_3479_nl;
  wire[0:0] mux_3478_nl;
  wire[0:0] mux_3477_nl;
  wire[0:0] mux_3476_nl;
  wire[0:0] mux_3475_nl;
  wire[0:0] mux_3474_nl;
  wire[0:0] mux_3473_nl;
  wire[0:0] mux_3472_nl;
  wire[0:0] mux_3470_nl;
  wire[0:0] mux_3469_nl;
  wire[0:0] mux_3466_nl;
  wire[0:0] mux_3465_nl;
  wire[0:0] mux_3464_nl;
  wire[0:0] mux_3463_nl;
  wire[0:0] mux_3462_nl;
  wire[0:0] mux_3461_nl;
  wire[0:0] mux_3460_nl;
  wire[0:0] mux_3457_nl;
  wire[0:0] mux_3455_nl;
  wire[0:0] mux_3454_nl;
  wire[0:0] mux_3453_nl;
  wire[0:0] mux_3451_nl;
  wire[0:0] mux_3448_nl;
  wire[0:0] mux_3447_nl;
  wire[0:0] mux_3446_nl;
  wire[0:0] mux_3445_nl;
  wire[0:0] mux_3444_nl;
  wire[0:0] mux_3443_nl;
  wire[0:0] mux_3442_nl;
  wire[0:0] mux_3441_nl;
  wire[0:0] mux_3440_nl;
  wire[0:0] mux_3439_nl;
  wire[0:0] mux_3438_nl;
  wire[0:0] mux_3437_nl;
  wire[0:0] mux_3435_nl;
  wire[0:0] mux_3434_nl;
  wire[0:0] mux_3433_nl;
  wire[0:0] mux_3432_nl;
  wire[0:0] mux_3431_nl;
  wire[0:0] mux_3429_nl;
  wire[0:0] mux_3428_nl;
  wire[0:0] mux_3427_nl;
  wire[0:0] mux_3425_nl;
  wire[0:0] mux_3424_nl;
  wire[0:0] mux_3420_nl;
  wire[0:0] mux_3506_nl;
  wire[0:0] mux_3505_nl;
  wire[0:0] or_3090_nl;
  wire[0:0] mux_3502_nl;
  wire[0:0] or_3084_nl;
  wire[0:0] mux_3501_nl;
  wire[0:0] or_3083_nl;
  wire[0:0] mux_3500_nl;
  wire[0:0] mux_3499_nl;
  wire[0:0] or_3079_nl;
  wire[0:0] mux_3497_nl;
  wire[0:0] mux_3496_nl;
  wire[0:0] nand_168_nl;
  wire[0:0] or_3076_nl;
  wire[0:0] or_3071_nl;
  wire[0:0] mux_3417_nl;
  wire[0:0] nor_569_nl;
  wire[0:0] mux_3416_nl;
  wire[0:0] or_3055_nl;
  wire[0:0] mux_3415_nl;
  wire[0:0] or_3054_nl;
  wire[0:0] or_3053_nl;
  wire[0:0] mux_3414_nl;
  wire[0:0] or_3052_nl;
  wire[0:0] or_3051_nl;
  wire[0:0] and_409_nl;
  wire[0:0] mux_3413_nl;
  wire[0:0] and_410_nl;
  wire[0:0] mux_3412_nl;
  wire[0:0] nor_570_nl;
  wire[0:0] nor_571_nl;
  wire[0:0] nor_572_nl;
  wire[0:0] mux_3411_nl;
  wire[0:0] or_3044_nl;
  wire[0:0] nand_208_nl;
  wire[0:0] mux_3513_nl;
  wire[0:0] mux_3512_nl;
  wire[0:0] mux_3511_nl;
  wire[0:0] or_3348_nl;
  wire[0:0] or_3349_nl;
  wire[0:0] mux_3510_nl;
  wire[0:0] or_3099_nl;
  wire[0:0] or_3350_nl;
  wire[0:0] mux_3509_nl;
  wire[0:0] or_3097_nl;
  wire[0:0] or_3095_nl;
  wire[0:0] nand_420_nl;
  wire[0:0] mux_3508_nl;
  wire[0:0] nor_567_nl;
  wire[0:0] and_402_nl;
  wire[0:0] mux_3507_nl;
  wire[0:0] or_3091_nl;
  wire[0:0] mux_3556_nl;
  wire[0:0] mux_3574_nl;
  wire[0:0] mux_3573_nl;
  wire[0:0] mux_3572_nl;
  wire[0:0] or_3120_nl;
  wire[0:0] mux_3056_nl;
  wire[0:0] mux_3570_nl;
  wire[0:0] mux_3569_nl;
  wire[0:0] mux_433_nl;
  wire[0:0] or_3119_nl;
  wire[0:0] mux_3567_nl;
  wire[0:0] mux_3566_nl;
  wire[0:0] mux_438_nl;
  wire[0:0] mux_437_nl;
  wire[0:0] mux_431_nl;
  wire[0:0] mux_3554_nl;
  wire[0:0] mux_420_nl;
  wire[0:0] mux_419_nl;
  wire[0:0] mux_3550_nl;
  wire[0:0] mux_3549_nl;
  wire[0:0] mux_3548_nl;
  wire[0:0] mux_3547_nl;
  wire[0:0] mux_3546_nl;
  wire[0:0] mux_403_nl;
  wire[0:0] or_3115_nl;
  wire[0:0] mux_3544_nl;
  wire[0:0] mux_3543_nl;
  wire[0:0] mux_3542_nl;
  wire[0:0] mux_402_nl;
  wire[0:0] mux_401_nl;
  wire[0:0] mux_400_nl;
  wire[0:0] mux_3536_nl;
  wire[0:0] mux_3535_nl;
  wire[0:0] mux_3534_nl;
  wire[0:0] mux_3533_nl;
  wire[0:0] nand_173_nl;
  wire[0:0] mux_3532_nl;
  wire[0:0] mux_3529_nl;
  wire[0:0] mux_3528_nl;
  wire[0:0] mux_3527_nl;
  wire[0:0] mux_383_nl;
  wire[0:0] mux_377_nl;
  wire[0:0] mux_376_nl;
  wire[0:0] COMP_LOOP_mux1h_477_nl;
  wire[0:0] COMP_LOOP_nor_14_nl;
  wire[0:0] mux_3577_nl;
  wire[0:0] mux_3576_nl;
  wire[0:0] mux_3562_nl;
  wire[0:0] mux_3561_nl;
  wire[0:0] mux_3560_nl;
  wire[0:0] mux_3559_nl;
  wire[0:0] mux_3558_nl;
  wire[0:0] mux_3584_nl;
  wire[0:0] mux_3583_nl;
  wire[0:0] nand_452_nl;
  wire[0:0] mux_3582_nl;
  wire[0:0] nor_558_nl;
  wire[0:0] nor_559_nl;
  wire[0:0] or_3474_nl;
  wire[0:0] mux_3581_nl;
  wire[0:0] or_3475_nl;
  wire[0:0] mux_3580_nl;
  wire[0:0] mux_3579_nl;
  wire[0:0] or_3127_nl;
  wire[0:0] or_3126_nl;
  wire[0:0] or_3125_nl;
  wire[0:0] nand_453_nl;
  wire[0:0] mux_3578_nl;
  wire[0:0] nor_562_nl;
  wire[0:0] nor_563_nl;
  wire[0:0] mux_3591_nl;
  wire[0:0] and_391_nl;
  wire[0:0] mux_3590_nl;
  wire[0:0] nor_552_nl;
  wire[0:0] mux_3589_nl;
  wire[0:0] or_3145_nl;
  wire[0:0] and_392_nl;
  wire[0:0] mux_3588_nl;
  wire[0:0] nor_554_nl;
  wire[0:0] mux_3587_nl;
  wire[0:0] mux_3586_nl;
  wire[0:0] nor_555_nl;
  wire[0:0] nor_556_nl;
  wire[0:0] mux_3585_nl;
  wire[0:0] or_3136_nl;
  wire[0:0] or_3135_nl;
  wire[0:0] nor_557_nl;
  wire[0:0] nor_540_nl;
  wire[0:0] COMP_LOOP_mux1h_479_nl;
  wire[0:0] COMP_LOOP_nor_17_nl;
  wire[0:0] mux_3598_nl;
  wire[0:0] or_3342_nl;
  wire[0:0] mux_3597_nl;
  wire[0:0] mux_3596_nl;
  wire[0:0] or_3158_nl;
  wire[0:0] or_3156_nl;
  wire[0:0] or_3155_nl;
  wire[0:0] mux_3595_nl;
  wire[0:0] mux_3594_nl;
  wire[0:0] or_3343_nl;
  wire[0:0] nand_419_nl;
  wire[0:0] mux_3593_nl;
  wire[0:0] nor_548_nl;
  wire[0:0] and_820_nl;
  wire[0:0] mux_3592_nl;
  wire[0:0] or_3344_nl;
  wire[0:0] or_3345_nl;
  wire[0:0] mux_3605_nl;
  wire[0:0] nor_538_nl;
  wire[0:0] mux_3604_nl;
  wire[0:0] nand_181_nl;
  wire[0:0] nand_180_nl;
  wire[0:0] mux_3602_nl;
  wire[0:0] nor_541_nl;
  wire[0:0] nor_542_nl;
  wire[0:0] mux_3601_nl;
  wire[0:0] and_389_nl;
  wire[0:0] mux_3600_nl;
  wire[0:0] mux_3599_nl;
  wire[0:0] nor_543_nl;
  wire[0:0] COMP_LOOP_mux1h_480_nl;
  wire[0:0] mux_3673_nl;
  wire[0:0] mux_3672_nl;
  wire[0:0] mux_3671_nl;
  wire[0:0] mux_3670_nl;
  wire[0:0] mux_3669_nl;
  wire[0:0] mux_3668_nl;
  wire[0:0] mux_3667_nl;
  wire[0:0] mux_3666_nl;
  wire[0:0] mux_3665_nl;
  wire[0:0] nand_195_nl;
  wire[0:0] mux_3664_nl;
  wire[0:0] and_388_nl;
  wire[0:0] mux_3663_nl;
  wire[0:0] mux_3662_nl;
  wire[0:0] mux_3661_nl;
  wire[0:0] mux_3660_nl;
  wire[0:0] mux_3659_nl;
  wire[0:0] and_386_nl;
  wire[0:0] mux_3658_nl;
  wire[0:0] mux_3657_nl;
  wire[0:0] or_3182_nl;
  wire[0:0] and_385_nl;
  wire[0:0] mux_3656_nl;
  wire[0:0] mux_3655_nl;
  wire[0:0] mux_3654_nl;
  wire[0:0] mux_3653_nl;
  wire[0:0] mux_3652_nl;
  wire[0:0] mux_3651_nl;
  wire[0:0] mux_3650_nl;
  wire[0:0] nand_196_nl;
  wire[0:0] mux_3649_nl;
  wire[0:0] mux_3648_nl;
  wire[0:0] mux_3647_nl;
  wire[0:0] mux_3646_nl;
  wire[0:0] mux_3645_nl;
  wire[0:0] mux_3644_nl;
  wire[0:0] mux_3643_nl;
  wire[0:0] mux_3642_nl;
  wire[0:0] mux_3641_nl;
  wire[0:0] mux_3640_nl;
  wire[0:0] mux_3639_nl;
  wire[0:0] nor_536_nl;
  wire[0:0] mux_3638_nl;
  wire[0:0] nand_197_nl;
  wire[0:0] mux_3637_nl;
  wire[0:0] mux_3636_nl;
  wire[0:0] mux_3635_nl;
  wire[0:0] mux_3634_nl;
  wire[0:0] mux_3633_nl;
  wire[0:0] mux_3632_nl;
  wire[0:0] mux_3631_nl;
  wire[0:0] mux_3630_nl;
  wire[0:0] mux_3629_nl;
  wire[0:0] mux_3627_nl;
  wire[0:0] mux_3626_nl;
  wire[0:0] mux_3625_nl;
  wire[0:0] mux_3624_nl;
  wire[0:0] mux_3623_nl;
  wire[0:0] mux_2589_nl;
  wire[0:0] mux_3622_nl;
  wire[0:0] or_3179_nl;
  wire[0:0] mux_3621_nl;
  wire[0:0] mux_3620_nl;
  wire[0:0] mux_3619_nl;
  wire[0:0] mux_3618_nl;
  wire[0:0] mux_3617_nl;
  wire[0:0] or_3178_nl;
  wire[0:0] mux_3616_nl;
  wire[0:0] or_3176_nl;
  wire[0:0] mux_3615_nl;
  wire[0:0] mux_3614_nl;
  wire[0:0] mux_3612_nl;
  wire[0:0] mux_3611_nl;
  wire[0:0] mux_3610_nl;
  wire[0:0] mux_3609_nl;
  wire[0:0] mux_3608_nl;
  wire[0:0] mux_3607_nl;
  wire[0:0] mux_3606_nl;
  wire[0:0] COMP_LOOP_or_28_nl;
  wire[0:0] mux_371_nl;
  wire[0:0] mux_372_nl;
  wire[0:0] mux_406_nl;
  wire[0:0] mux_1027_nl;
  wire[0:0] or_3295_nl;
  wire[0:0] and_659_nl;
  wire[0:0] nor_1193_nl;
  wire[0:0] or_579_nl;
  wire[0:0] mux_1061_nl;
  wire[0:0] or_578_nl;
  wire[0:0] or_577_nl;
  wire[0:0] mux_1066_nl;
  wire[0:0] mux_1065_nl;
  wire[0:0] or_587_nl;
  wire[0:0] or_586_nl;
  wire[0:0] or_585_nl;
  wire[0:0] or_583_nl;
  wire[0:0] or_591_nl;
  wire[0:0] or_589_nl;
  wire[0:0] mux_1087_nl;
  wire[0:0] or_614_nl;
  wire[0:0] or_613_nl;
  wire[0:0] mux_1086_nl;
  wire[0:0] or_611_nl;
  wire[0:0] or_610_nl;
  wire[0:0] mux_1080_nl;
  wire[0:0] nor_1170_nl;
  wire[0:0] nor_1171_nl;
  wire[0:0] or_600_nl;
  wire[0:0] or_599_nl;
  wire[0:0] or_693_nl;
  wire[0:0] mux_1138_nl;
  wire[0:0] or_692_nl;
  wire[0:0] or_691_nl;
  wire[0:0] mux_1149_nl;
  wire[0:0] mux_1148_nl;
  wire[0:0] or_709_nl;
  wire[0:0] or_708_nl;
  wire[0:0] or_707_nl;
  wire[0:0] or_705_nl;
  wire[0:0] or_712_nl;
  wire[0:0] or_710_nl;
  wire[0:0] or_792_nl;
  wire[0:0] mux_1205_nl;
  wire[0:0] or_791_nl;
  wire[0:0] or_790_nl;
  wire[0:0] mux_1210_nl;
  wire[0:0] mux_1209_nl;
  wire[0:0] or_800_nl;
  wire[0:0] or_799_nl;
  wire[0:0] or_798_nl;
  wire[0:0] or_796_nl;
  wire[0:0] or_804_nl;
  wire[0:0] or_802_nl;
  wire[0:0] or_906_nl;
  wire[0:0] mux_1282_nl;
  wire[0:0] or_905_nl;
  wire[0:0] or_904_nl;
  wire[0:0] mux_1293_nl;
  wire[0:0] mux_1292_nl;
  wire[0:0] or_922_nl;
  wire[0:0] or_921_nl;
  wire[0:0] nand_433_nl;
  wire[0:0] or_918_nl;
  wire[0:0] or_925_nl;
  wire[0:0] or_923_nl;
  wire[0:0] or_1005_nl;
  wire[0:0] mux_1349_nl;
  wire[0:0] or_1004_nl;
  wire[0:0] or_1003_nl;
  wire[0:0] mux_1354_nl;
  wire[0:0] mux_1353_nl;
  wire[0:0] or_1013_nl;
  wire[0:0] or_1012_nl;
  wire[0:0] or_1011_nl;
  wire[0:0] or_1009_nl;
  wire[0:0] or_1017_nl;
  wire[0:0] or_1015_nl;
  wire[0:0] or_1119_nl;
  wire[0:0] mux_1426_nl;
  wire[0:0] or_1118_nl;
  wire[0:0] or_1117_nl;
  wire[0:0] mux_1437_nl;
  wire[0:0] mux_1436_nl;
  wire[0:0] or_1135_nl;
  wire[0:0] or_1134_nl;
  wire[0:0] nand_432_nl;
  wire[0:0] or_1131_nl;
  wire[0:0] or_1138_nl;
  wire[0:0] or_1136_nl;
  wire[0:0] or_1218_nl;
  wire[0:0] mux_1493_nl;
  wire[0:0] or_1217_nl;
  wire[0:0] or_1216_nl;
  wire[0:0] mux_1498_nl;
  wire[0:0] mux_1497_nl;
  wire[0:0] or_1226_nl;
  wire[0:0] or_1225_nl;
  wire[0:0] nand_431_nl;
  wire[0:0] or_1222_nl;
  wire[0:0] or_1230_nl;
  wire[0:0] or_1228_nl;
  wire[0:0] or_1332_nl;
  wire[0:0] mux_1570_nl;
  wire[0:0] or_1331_nl;
  wire[0:0] or_1330_nl;
  wire[0:0] mux_1581_nl;
  wire[0:0] mux_1580_nl;
  wire[0:0] or_1348_nl;
  wire[0:0] or_1347_nl;
  wire[0:0] nand_430_nl;
  wire[0:0] or_1344_nl;
  wire[0:0] nand_418_nl;
  wire[0:0] or_1349_nl;
  wire[0:0] or_1431_nl;
  wire[0:0] mux_1637_nl;
  wire[0:0] or_1430_nl;
  wire[0:0] or_1429_nl;
  wire[0:0] mux_1642_nl;
  wire[0:0] mux_1641_nl;
  wire[0:0] or_1439_nl;
  wire[0:0] or_1438_nl;
  wire[0:0] or_1437_nl;
  wire[0:0] or_1435_nl;
  wire[0:0] or_1443_nl;
  wire[0:0] or_1441_nl;
  wire[0:0] or_1545_nl;
  wire[0:0] mux_1714_nl;
  wire[0:0] or_1544_nl;
  wire[0:0] or_1543_nl;
  wire[0:0] mux_1725_nl;
  wire[0:0] mux_1724_nl;
  wire[0:0] or_1561_nl;
  wire[0:0] or_1560_nl;
  wire[0:0] nand_429_nl;
  wire[0:0] or_1557_nl;
  wire[0:0] or_1564_nl;
  wire[0:0] or_1562_nl;
  wire[0:0] or_1644_nl;
  wire[0:0] mux_1781_nl;
  wire[0:0] or_1643_nl;
  wire[0:0] or_1642_nl;
  wire[0:0] mux_1786_nl;
  wire[0:0] mux_1785_nl;
  wire[0:0] or_1652_nl;
  wire[0:0] or_1651_nl;
  wire[0:0] nand_428_nl;
  wire[0:0] or_1648_nl;
  wire[0:0] or_1656_nl;
  wire[0:0] or_1654_nl;
  wire[0:0] or_1758_nl;
  wire[0:0] mux_1858_nl;
  wire[0:0] or_1757_nl;
  wire[0:0] or_1756_nl;
  wire[0:0] mux_1869_nl;
  wire[0:0] mux_1868_nl;
  wire[0:0] or_1774_nl;
  wire[0:0] or_1773_nl;
  wire[0:0] nand_427_nl;
  wire[0:0] or_1770_nl;
  wire[0:0] nand_416_nl;
  wire[0:0] or_1775_nl;
  wire[0:0] mux_1922_nl;
  wire[0:0] or_1853_nl;
  wire[0:0] or_1852_nl;
  wire[0:0] nand_73_nl;
  wire[0:0] mux_1926_nl;
  wire[0:0] nor_874_nl;
  wire[0:0] nor_875_nl;
  wire[0:0] or_1857_nl;
  wire[0:0] mux_1925_nl;
  wire[0:0] or_1856_nl;
  wire[0:0] or_1855_nl;
  wire[0:0] mux_1929_nl;
  wire[0:0] nor_872_nl;
  wire[0:0] nor_873_nl;
  wire[0:0] or_1974_nl;
  wire[0:0] mux_2003_nl;
  wire[0:0] or_1973_nl;
  wire[0:0] or_1972_nl;
  wire[0:0] mux_2014_nl;
  wire[0:0] mux_2013_nl;
  wire[0:0] or_1990_nl;
  wire[0:0] or_1989_nl;
  wire[0:0] nand_426_nl;
  wire[0:0] or_1986_nl;
  wire[0:0] nand_414_nl;
  wire[0:0] or_1991_nl;
  wire[0:0] or_2073_nl;
  wire[0:0] mux_2070_nl;
  wire[0:0] or_2072_nl;
  wire[0:0] or_2071_nl;
  wire[0:0] mux_2075_nl;
  wire[0:0] mux_2074_nl;
  wire[0:0] or_2081_nl;
  wire[0:0] or_2080_nl;
  wire[0:0] nand_425_nl;
  wire[0:0] or_2077_nl;
  wire[0:0] nand_412_nl;
  wire[0:0] or_2083_nl;
  wire[0:0] or_2187_nl;
  wire[0:0] mux_2147_nl;
  wire[0:0] nand_291_nl;
  wire[0:0] or_2185_nl;
  wire[0:0] mux_2158_nl;
  wire[0:0] mux_2157_nl;
  wire[0:0] nand_288_nl;
  wire[0:0] nand_289_nl;
  wire[0:0] nand_424_nl;
  wire[0:0] or_2199_nl;
  wire[0:0] nand_410_nl;
  wire[0:0] or_2204_nl;
  wire[0:0] mux_2240_nl;
  wire[0:0] mux_2289_nl;
  wire[0:0] mux_2310_nl;
  wire[0:0] or_2393_nl;
  wire[0:0] mux_2427_nl;
  wire[0:0] or_2409_nl;
  wire[0:0] mux_2474_nl;
  wire[0:0] mux_2473_nl;
  wire[0:0] or_2425_nl;
  wire[0:0] mux_2472_nl;
  wire[0:0] or_2424_nl;
  wire[0:0] mux_2471_nl;
  wire[0:0] mux_2470_nl;
  wire[0:0] or_3285_nl;
  wire[0:0] mux_2469_nl;
  wire[0:0] or_2419_nl;
  wire[0:0] mux_2468_nl;
  wire[0:0] or_2417_nl;
  wire[0:0] mux_2467_nl;
  wire[0:0] nand_111_nl;
  wire[0:0] mux_2465_nl;
  wire[0:0] or_2412_nl;
  wire[0:0] mux_2464_nl;
  wire[0:0] nand_110_nl;
  wire[0:0] mux_2462_nl;
  wire[0:0] nor_756_nl;
  wire[0:0] nor_757_nl;
  wire[0:0] mux_2488_nl;
  wire[0:0] mux_2487_nl;
  wire[0:0] mux_2486_nl;
  wire[0:0] nor_743_nl;
  wire[0:0] nor_744_nl;
  wire[0:0] nor_745_nl;
  wire[0:0] mux_3706_nl;
  wire[0:0] or_3233_nl;
  wire[0:0] or_3232_nl;
  wire[0:0] mux_2484_nl;
  wire[0:0] nor_746_nl;
  wire[0:0] mux_2483_nl;
  wire[0:0] or_2441_nl;
  wire[0:0] or_2439_nl;
  wire[0:0] and_558_nl;
  wire[0:0] mux_89_nl;
  wire[0:0] nor_1285_nl;
  wire[0:0] nor_1286_nl;
  wire[0:0] mux_2481_nl;
  wire[0:0] mux_2480_nl;
  wire[0:0] mux_2479_nl;
  wire[0:0] mux_2478_nl;
  wire[0:0] nor_750_nl;
  wire[0:0] nor_1278_nl;
  wire[0:0] and_796_nl;
  wire[0:0] mux_94_nl;
  wire[0:0] mux_93_nl;
  wire[0:0] nor_1280_nl;
  wire[0:0] nor_1281_nl;
  wire[0:0] mux_2492_nl;
  wire[0:0] mux_2491_nl;
  wire[0:0] mux_2490_nl;
  wire[0:0] or_463_nl;
  wire[0:0] mux_2496_nl;
  wire[0:0] nor_741_nl;
  wire[0:0] nor_742_nl;
  wire[0:0] or_2468_nl;
  wire[0:0] or_2489_nl;
  wire[0:0] nand_117_nl;
  wire[0:0] nor_719_nl;
  wire[0:0] or_2556_nl;
  wire[0:0] or_2555_nl;
  wire[0:0] mux_2756_nl;
  wire[0:0] mux_2755_nl;
  wire[0:0] mux_2754_nl;
  wire[0:0] nor_702_nl;
  wire[0:0] mux_2753_nl;
  wire[0:0] nor_704_nl;
  wire[0:0] nor_705_nl;
  wire[0:0] mux_2752_nl;
  wire[0:0] nor_706_nl;
  wire[0:0] mux_2751_nl;
  wire[0:0] nor_707_nl;
  wire[0:0] mux_2750_nl;
  wire[0:0] nor_708_nl;
  wire[0:0] nor_1296_nl;
  wire[0:0] mux_2749_nl;
  wire[0:0] mux_2748_nl;
  wire[0:0] nor_710_nl;
  wire[0:0] mux_2747_nl;
  wire[0:0] nor_711_nl;
  wire[0:0] nor_712_nl;
  wire[0:0] nor_713_nl;
  wire[0:0] mux_2745_nl;
  wire[0:0] or_2553_nl;
  wire[0:0] mux_74_nl;
  wire[0:0] or_53_nl;
  wire[0:0] or_51_nl;
  wire[0:0] nand_120_nl;
  wire[0:0] or_2578_nl;
  wire[0:0] or_2621_nl;
  wire[0:0] mux_2799_nl;
  wire[0:0] mux_2871_nl;
  wire[0:0] or_207_nl;
  wire[0:0] mux_2880_nl;
  wire[0:0] and_503_nl;
  wire[0:0] mux_2879_nl;
  wire[0:0] mux_2878_nl;
  wire[0:0] nor_672_nl;
  wire[0:0] nor_673_nl;
  wire[0:0] nor_674_nl;
  wire[0:0] mux_2877_nl;
  wire[0:0] or_2662_nl;
  wire[0:0] mux_2876_nl;
  wire[0:0] or_2659_nl;
  wire[0:0] mux_2875_nl;
  wire[0:0] mux_2874_nl;
  wire[0:0] nor_675_nl;
  wire[0:0] mux_2873_nl;
  wire[0:0] and_505_nl;
  wire[0:0] mux_2872_nl;
  wire[0:0] nor_676_nl;
  wire[0:0] mux_2870_nl;
  wire[0:0] or_2647_nl;
  wire[0:0] mux_2902_nl;
  wire[0:0] mux_2901_nl;
  wire[0:0] and_498_nl;
  wire[0:0] mux_2900_nl;
  wire[0:0] nor_654_nl;
  wire[0:0] mux_2899_nl;
  wire[0:0] nor_655_nl;
  wire[0:0] nor_656_nl;
  wire[0:0] mux_2898_nl;
  wire[0:0] nor_657_nl;
  wire[0:0] and_499_nl;
  wire[0:0] mux_2897_nl;
  wire[0:0] nor_658_nl;
  wire[0:0] mux_2896_nl;
  wire[0:0] or_2699_nl;
  wire[0:0] mux_2895_nl;
  wire[0:0] nor_659_nl;
  wire[0:0] nor_660_nl;
  wire[0:0] mux_2894_nl;
  wire[0:0] mux_2893_nl;
  wire[0:0] nor_661_nl;
  wire[0:0] mux_2892_nl;
  wire[0:0] or_2693_nl;
  wire[0:0] and_500_nl;
  wire[0:0] mux_2891_nl;
  wire[0:0] nor_662_nl;
  wire[0:0] nor_663_nl;
  wire[0:0] mux_2890_nl;
  wire[0:0] nor_664_nl;
  wire[0:0] nor_665_nl;
  wire[0:0] mux_523_nl;
  wire[0:0] or_248_nl;
  wire[0:0] mux_2910_nl;
  wire[0:0] mux_2920_nl;
  wire[0:0] mux_520_nl;
  wire[0:0] mux_3168_nl;
  wire[0:0] nor_627_nl;
  wire[0:0] nor_628_nl;
  wire[0:0] or_3260_nl;
  wire[0:0] mux_3213_nl;
  wire[0:0] or_2886_nl;
  wire[0:0] nand_220_nl;
  wire[0:0] mux_3212_nl;
  wire[0:0] or_2882_nl;
  wire[0:0] mux_3235_nl;
  wire[0:0] or_2905_nl;
  wire[0:0] or_2904_nl;
  wire[0:0] mux_3279_nl;
  wire[0:0] and_436_nl;
  wire[0:0] mux_3368_nl;
  wire[0:0] mux_3354_nl;
  wire[0:0] mux_3353_nl;
  wire[0:0] mux_3352_nl;
  wire[0:0] mux_3351_nl;
  wire[0:0] mux_3350_nl;
  wire[0:0] mux_3382_nl;
  wire[0:0] mux_3381_nl;
  wire[0:0] mux_3380_nl;
  wire[0:0] and_417_nl;
  wire[0:0] mux_3378_nl;
  wire[0:0] mux_3377_nl;
  wire[0:0] nor_591_nl;
  wire[0:0] nor_1295_nl;
  wire[0:0] mux_3376_nl;
  wire[0:0] mux_3375_nl;
  wire[0:0] and_418_nl;
  wire[0:0] mux_3374_nl;
  wire[0:0] nor_594_nl;
  wire[0:0] nor_595_nl;
  wire[0:0] nor_596_nl;
  wire[0:0] mux_3372_nl;
  wire[0:0] mux_3371_nl;
  wire[0:0] nor_1287_nl;
  wire[0:0] and_419_nl;
  wire[0:0] or_3007_nl;
  wire[0:0] or_3006_nl;
  wire[0:0] mux_3409_nl;
  wire[0:0] nor_573_nl;
  wire[0:0] mux_3408_nl;
  wire[0:0] mux_3407_nl;
  wire[0:0] or_3037_nl;
  wire[0:0] mux_3406_nl;
  wire[0:0] mux_3421_nl;
  wire[0:0] nor_568_nl;
  wire[0:0] mux_3613_nl;
  wire[0:0] mux_2664_nl;
  wire[0:0] mux_2663_nl;
  wire[0:0] mux_2662_nl;
  wire[0:0] nor_724_nl;
  wire[0:0] mux_2661_nl;
  wire[0:0] and_521_nl;
  wire[0:0] or_2522_nl;
  wire[2:0] STAGE_LOOP_acc_nl;
  wire[3:0] nl_STAGE_LOOP_acc_nl;
  wire[0:0] and_139_nl;
  wire[0:0] mux_1044_nl;
  wire[0:0] mux_1043_nl;
  wire[0:0] nor_1194_nl;
  wire[0:0] mux_1042_nl;
  wire[0:0] or_533_nl;
  wire[0:0] or_532_nl;
  wire[0:0] mux_1041_nl;
  wire[0:0] or_531_nl;
  wire[0:0] mux_1040_nl;
  wire[0:0] nor_1195_nl;
  wire[0:0] mux_1039_nl;
  wire[0:0] or_527_nl;
  wire[0:0] mux_1038_nl;
  wire[0:0] mux_1037_nl;
  wire[0:0] or_524_nl;
  wire[0:0] or_523_nl;
  wire[0:0] and_660_nl;
  wire[0:0] mux_1036_nl;
  wire[0:0] mux_1035_nl;
  wire[0:0] nor_1196_nl;
  wire[0:0] nor_1197_nl;
  wire[0:0] nor_1198_nl;
  wire[0:0] mux_1034_nl;
  wire[0:0] nor_1199_nl;
  wire[0:0] mux_1033_nl;
  wire[0:0] mux_1032_nl;
  wire[0:0] or_516_nl;
  wire[0:0] or_514_nl;
  wire[0:0] mux_1031_nl;
  wire[0:0] and_661_nl;
  wire[0:0] mux_1030_nl;
  wire[0:0] or_512_nl;
  wire[0:0] nor_1200_nl;
  wire[0:0] and_145_nl;
  wire[0:0] and_153_nl;
  wire[0:0] mux_1046_nl;
  wire[0:0] nor_1191_nl;
  wire[0:0] nor_1192_nl;
  wire[0:0] and_162_nl;
  wire[0:0] mux_1047_nl;
  wire[0:0] nor_1189_nl;
  wire[0:0] nor_1190_nl;
  wire[0:0] and_170_nl;
  wire[0:0] mux_1048_nl;
  wire[0:0] nor_1187_nl;
  wire[0:0] nor_1188_nl;
  wire[0:0] and_179_nl;
  wire[0:0] and_188_nl;
  wire[0:0] mux_1050_nl;
  wire[0:0] nor_1185_nl;
  wire[0:0] nor_1186_nl;
  wire[0:0] and_197_nl;
  wire[0:0] mux_1051_nl;
  wire[0:0] nor_1183_nl;
  wire[0:0] nor_1184_nl;
  wire[0:0] and_205_nl;
  wire[0:0] mux_1052_nl;
  wire[0:0] nor_1181_nl;
  wire[0:0] nor_1182_nl;
  wire[0:0] and_211_nl;
  wire[0:0] mux_1053_nl;
  wire[0:0] nor_1179_nl;
  wire[0:0] nor_1180_nl;
  wire[0:0] and_220_nl;
  wire[0:0] mux_1054_nl;
  wire[0:0] nor_1177_nl;
  wire[0:0] nor_1178_nl;
  wire[0:0] and_231_nl;
  wire[0:0] and_238_nl;
  wire[0:0] mux_1055_nl;
  wire[0:0] nor_1175_nl;
  wire[0:0] nor_1176_nl;
  wire[0:0] and_246_nl;
  wire[0:0] mux_1056_nl;
  wire[0:0] and_817_nl;
  wire[0:0] nor_1174_nl;
  wire[0:0] and_253_nl;
  wire[0:0] mux_1057_nl;
  wire[0:0] and_657_nl;
  wire[0:0] nor_1172_nl;
  wire[0:0] and_261_nl;
  wire[0:0] mux_1098_nl;
  wire[0:0] mux_1097_nl;
  wire[0:0] mux_1096_nl;
  wire[0:0] mux_1095_nl;
  wire[0:0] mux_1094_nl;
  wire[0:0] mux_1093_nl;
  wire[0:0] or_624_nl;
  wire[0:0] mux_1091_nl;
  wire[0:0] mux_1090_nl;
  wire[0:0] or_615_nl;
  wire[0:0] mux_1089_nl;
  wire[0:0] mux_1085_nl;
  wire[0:0] mux_1084_nl;
  wire[0:0] mux_1083_nl;
  wire[0:0] mux_1082_nl;
  wire[0:0] or_605_nl;
  wire[0:0] mux_1081_nl;
  wire[0:0] mux_1079_nl;
  wire[0:0] mux_1078_nl;
  wire[0:0] mux_1077_nl;
  wire[0:0] mux_1076_nl;
  wire[0:0] or_602_nl;
  wire[0:0] mux_1075_nl;
  wire[0:0] mux_1074_nl;
  wire[0:0] or_597_nl;
  wire[0:0] mux_1072_nl;
  wire[0:0] mux_1071_nl;
  wire[0:0] mux_1070_nl;
  wire[0:0] or_594_nl;
  wire[0:0] mux_1069_nl;
  wire[0:0] or_592_nl;
  wire[0:0] or_588_nl;
  wire[0:0] mux_1064_nl;
  wire[0:0] mux_1063_nl;
  wire[0:0] or_581_nl;
  wire[0:0] or_580_nl;
  wire[0:0] mux_1060_nl;
  wire[0:0] mux_1059_nl;
  wire[0:0] mux_1058_nl;
  wire[0:0] or_573_nl;
  wire[0:0] or_570_nl;
  wire[0:0] or_569_nl;
  wire[0:0] mux_1128_nl;
  wire[0:0] mux_1127_nl;
  wire[0:0] and_654_nl;
  wire[0:0] mux_1126_nl;
  wire[0:0] nor_1147_nl;
  wire[0:0] mux_1125_nl;
  wire[0:0] nor_1149_nl;
  wire[0:0] mux_1124_nl;
  wire[0:0] nor_1150_nl;
  wire[0:0] mux_1123_nl;
  wire[0:0] or_670_nl;
  wire[0:0] or_669_nl;
  wire[0:0] mux_1122_nl;
  wire[0:0] nor_1151_nl;
  wire[0:0] nor_1152_nl;
  wire[0:0] mux_1121_nl;
  wire[0:0] mux_1120_nl;
  wire[0:0] nor_1153_nl;
  wire[0:0] mux_1119_nl;
  wire[0:0] nor_1154_nl;
  wire[0:0] mux_1118_nl;
  wire[0:0] or_661_nl;
  wire[0:0] or_659_nl;
  wire[0:0] nor_1155_nl;
  wire[0:0] mux_1117_nl;
  wire[0:0] nor_1156_nl;
  wire[0:0] and_655_nl;
  wire[0:0] mux_1116_nl;
  wire[0:0] nor_1157_nl;
  wire[0:0] mux_1115_nl;
  wire[0:0] nor_1158_nl;
  wire[0:0] mux_1114_nl;
  wire[0:0] mux_1113_nl;
  wire[0:0] nor_1160_nl;
  wire[0:0] mux_1112_nl;
  wire[0:0] mux_1111_nl;
  wire[0:0] or_650_nl;
  wire[0:0] or_649_nl;
  wire[0:0] mux_1110_nl;
  wire[0:0] or_648_nl;
  wire[0:0] or_646_nl;
  wire[0:0] mux_1109_nl;
  wire[0:0] mux_1108_nl;
  wire[0:0] nor_1161_nl;
  wire[0:0] nor_1162_nl;
  wire[0:0] mux_1107_nl;
  wire[0:0] or_641_nl;
  wire[0:0] mux_1106_nl;
  wire[0:0] nor_1163_nl;
  wire[0:0] nor_1164_nl;
  wire[0:0] mux_1105_nl;
  wire[0:0] nor_1165_nl;
  wire[0:0] mux_1104_nl;
  wire[0:0] mux_1103_nl;
  wire[0:0] or_635_nl;
  wire[0:0] mux_1102_nl;
  wire[0:0] or_633_nl;
  wire[0:0] or_630_nl;
  wire[0:0] mux_1101_nl;
  wire[0:0] and_656_nl;
  wire[0:0] mux_1100_nl;
  wire[0:0] nor_1166_nl;
  wire[0:0] mux_1099_nl;
  wire[0:0] nor_1167_nl;
  wire[0:0] nor_1168_nl;
  wire[0:0] nor_1169_nl;
  wire[0:0] mux_1170_nl;
  wire[0:0] mux_1169_nl;
  wire[0:0] mux_1168_nl;
  wire[0:0] mux_1167_nl;
  wire[0:0] or_730_nl;
  wire[0:0] mux_1166_nl;
  wire[0:0] or_728_nl;
  wire[0:0] or_727_nl;
  wire[0:0] mux_1165_nl;
  wire[0:0] mux_1164_nl;
  wire[0:0] or_726_nl;
  wire[0:0] or_725_nl;
  wire[0:0] mux_1163_nl;
  wire[0:0] mux_1162_nl;
  wire[0:0] mux_1161_nl;
  wire[0:0] or_724_nl;
  wire[0:0] or_723_nl;
  wire[0:0] mux_1160_nl;
  wire[0:0] mux_1159_nl;
  wire[0:0] mux_1158_nl;
  wire[0:0] mux_1157_nl;
  wire[0:0] mux_1156_nl;
  wire[0:0] or_722_nl;
  wire[0:0] mux_1154_nl;
  wire[0:0] mux_1153_nl;
  wire[0:0] or_713_nl;
  wire[0:0] mux_1151_nl;
  wire[0:0] mux_1144_nl;
  wire[0:0] mux_1143_nl;
  wire[0:0] mux_1142_nl;
  wire[0:0] mux_1141_nl;
  wire[0:0] or_694_nl;
  wire[0:0] mux_1140_nl;
  wire[0:0] mux_1136_nl;
  wire[0:0] mux_1135_nl;
  wire[0:0] mux_1134_nl;
  wire[0:0] mux_1133_nl;
  wire[0:0] or_685_nl;
  wire[0:0] mux_1132_nl;
  wire[0:0] mux_1131_nl;
  wire[0:0] or_678_nl;
  wire[0:0] nor_224_nl;
  wire[0:0] mux_1200_nl;
  wire[0:0] mux_1199_nl;
  wire[0:0] and_651_nl;
  wire[0:0] mux_1198_nl;
  wire[0:0] nor_1122_nl;
  wire[0:0] mux_1197_nl;
  wire[0:0] nor_1124_nl;
  wire[0:0] mux_1196_nl;
  wire[0:0] nor_1125_nl;
  wire[0:0] mux_1195_nl;
  wire[0:0] or_776_nl;
  wire[0:0] or_775_nl;
  wire[0:0] mux_1194_nl;
  wire[0:0] nor_1126_nl;
  wire[0:0] nor_1127_nl;
  wire[0:0] mux_1193_nl;
  wire[0:0] mux_1192_nl;
  wire[0:0] nor_1128_nl;
  wire[0:0] mux_1191_nl;
  wire[0:0] nor_1129_nl;
  wire[0:0] mux_1190_nl;
  wire[0:0] or_767_nl;
  wire[0:0] or_765_nl;
  wire[0:0] nor_1130_nl;
  wire[0:0] mux_1189_nl;
  wire[0:0] nor_1131_nl;
  wire[0:0] and_652_nl;
  wire[0:0] mux_1188_nl;
  wire[0:0] nor_1132_nl;
  wire[0:0] mux_1187_nl;
  wire[0:0] nor_1133_nl;
  wire[0:0] mux_1186_nl;
  wire[0:0] mux_1185_nl;
  wire[0:0] nor_1135_nl;
  wire[0:0] mux_1184_nl;
  wire[0:0] mux_1183_nl;
  wire[0:0] or_756_nl;
  wire[0:0] or_755_nl;
  wire[0:0] mux_1182_nl;
  wire[0:0] or_754_nl;
  wire[0:0] or_752_nl;
  wire[0:0] mux_1181_nl;
  wire[0:0] mux_1180_nl;
  wire[0:0] nor_1136_nl;
  wire[0:0] nor_1137_nl;
  wire[0:0] mux_1179_nl;
  wire[0:0] or_747_nl;
  wire[0:0] mux_1178_nl;
  wire[0:0] nor_1138_nl;
  wire[0:0] nor_1139_nl;
  wire[0:0] mux_1177_nl;
  wire[0:0] nor_1140_nl;
  wire[0:0] mux_1176_nl;
  wire[0:0] mux_1175_nl;
  wire[0:0] or_741_nl;
  wire[0:0] mux_1174_nl;
  wire[0:0] or_739_nl;
  wire[0:0] or_736_nl;
  wire[0:0] mux_1173_nl;
  wire[0:0] and_653_nl;
  wire[0:0] mux_1172_nl;
  wire[0:0] nor_1141_nl;
  wire[0:0] mux_1171_nl;
  wire[0:0] nor_1142_nl;
  wire[0:0] nor_1143_nl;
  wire[0:0] nor_1144_nl;
  wire[0:0] mux_1242_nl;
  wire[0:0] mux_1241_nl;
  wire[0:0] mux_1240_nl;
  wire[0:0] mux_1239_nl;
  wire[0:0] mux_1238_nl;
  wire[0:0] mux_1237_nl;
  wire[0:0] or_837_nl;
  wire[0:0] mux_1235_nl;
  wire[0:0] mux_1234_nl;
  wire[0:0] or_828_nl;
  wire[0:0] mux_1233_nl;
  wire[0:0] mux_1229_nl;
  wire[0:0] mux_1228_nl;
  wire[0:0] mux_1227_nl;
  wire[0:0] mux_1226_nl;
  wire[0:0] or_818_nl;
  wire[0:0] mux_1225_nl;
  wire[0:0] mux_1223_nl;
  wire[0:0] mux_1222_nl;
  wire[0:0] mux_1221_nl;
  wire[0:0] mux_1220_nl;
  wire[0:0] or_815_nl;
  wire[0:0] mux_1219_nl;
  wire[0:0] mux_1218_nl;
  wire[0:0] or_810_nl;
  wire[0:0] mux_1216_nl;
  wire[0:0] mux_1215_nl;
  wire[0:0] mux_1214_nl;
  wire[0:0] or_807_nl;
  wire[0:0] mux_1213_nl;
  wire[0:0] or_805_nl;
  wire[0:0] or_801_nl;
  wire[0:0] mux_1208_nl;
  wire[0:0] mux_1207_nl;
  wire[0:0] or_794_nl;
  wire[0:0] or_793_nl;
  wire[0:0] mux_1204_nl;
  wire[0:0] mux_1203_nl;
  wire[0:0] mux_1202_nl;
  wire[0:0] or_786_nl;
  wire[0:0] or_783_nl;
  wire[0:0] or_782_nl;
  wire[0:0] mux_1272_nl;
  wire[0:0] mux_1271_nl;
  wire[0:0] and_648_nl;
  wire[0:0] mux_1270_nl;
  wire[0:0] nor_1097_nl;
  wire[0:0] mux_1269_nl;
  wire[0:0] nor_1099_nl;
  wire[0:0] mux_1268_nl;
  wire[0:0] nor_1100_nl;
  wire[0:0] mux_1267_nl;
  wire[0:0] or_883_nl;
  wire[0:0] or_882_nl;
  wire[0:0] mux_1266_nl;
  wire[0:0] nor_1101_nl;
  wire[0:0] nor_1102_nl;
  wire[0:0] mux_1265_nl;
  wire[0:0] mux_1264_nl;
  wire[0:0] nor_1103_nl;
  wire[0:0] mux_1263_nl;
  wire[0:0] nor_1104_nl;
  wire[0:0] mux_1262_nl;
  wire[0:0] or_874_nl;
  wire[0:0] or_872_nl;
  wire[0:0] nor_1105_nl;
  wire[0:0] mux_1261_nl;
  wire[0:0] nor_1106_nl;
  wire[0:0] and_649_nl;
  wire[0:0] mux_1260_nl;
  wire[0:0] nor_1107_nl;
  wire[0:0] mux_1259_nl;
  wire[0:0] nor_1108_nl;
  wire[0:0] mux_1258_nl;
  wire[0:0] mux_1257_nl;
  wire[0:0] nor_1110_nl;
  wire[0:0] mux_1256_nl;
  wire[0:0] mux_1255_nl;
  wire[0:0] or_863_nl;
  wire[0:0] or_862_nl;
  wire[0:0] mux_1254_nl;
  wire[0:0] or_861_nl;
  wire[0:0] or_859_nl;
  wire[0:0] mux_1253_nl;
  wire[0:0] mux_1252_nl;
  wire[0:0] nor_1111_nl;
  wire[0:0] nor_1112_nl;
  wire[0:0] mux_1251_nl;
  wire[0:0] or_854_nl;
  wire[0:0] mux_1250_nl;
  wire[0:0] nor_1113_nl;
  wire[0:0] nor_1114_nl;
  wire[0:0] mux_1249_nl;
  wire[0:0] nor_1115_nl;
  wire[0:0] mux_1248_nl;
  wire[0:0] mux_1247_nl;
  wire[0:0] or_848_nl;
  wire[0:0] mux_1246_nl;
  wire[0:0] or_846_nl;
  wire[0:0] or_843_nl;
  wire[0:0] mux_1245_nl;
  wire[0:0] and_650_nl;
  wire[0:0] mux_1244_nl;
  wire[0:0] nor_1116_nl;
  wire[0:0] mux_1243_nl;
  wire[0:0] nor_1117_nl;
  wire[0:0] nor_1118_nl;
  wire[0:0] nor_1119_nl;
  wire[0:0] mux_1314_nl;
  wire[0:0] mux_1313_nl;
  wire[0:0] mux_1312_nl;
  wire[0:0] mux_1311_nl;
  wire[0:0] or_943_nl;
  wire[0:0] mux_1310_nl;
  wire[0:0] or_941_nl;
  wire[0:0] or_940_nl;
  wire[0:0] mux_1309_nl;
  wire[0:0] mux_1308_nl;
  wire[0:0] or_939_nl;
  wire[0:0] or_938_nl;
  wire[0:0] mux_1307_nl;
  wire[0:0] mux_1306_nl;
  wire[0:0] mux_1305_nl;
  wire[0:0] or_937_nl;
  wire[0:0] or_936_nl;
  wire[0:0] mux_1304_nl;
  wire[0:0] mux_1303_nl;
  wire[0:0] mux_1302_nl;
  wire[0:0] mux_1301_nl;
  wire[0:0] mux_1300_nl;
  wire[0:0] or_935_nl;
  wire[0:0] mux_1298_nl;
  wire[0:0] mux_1297_nl;
  wire[0:0] or_926_nl;
  wire[0:0] mux_1295_nl;
  wire[0:0] mux_1288_nl;
  wire[0:0] mux_1287_nl;
  wire[0:0] mux_1286_nl;
  wire[0:0] mux_1285_nl;
  wire[0:0] or_907_nl;
  wire[0:0] mux_1284_nl;
  wire[0:0] mux_1280_nl;
  wire[0:0] mux_1279_nl;
  wire[0:0] mux_1278_nl;
  wire[0:0] mux_1277_nl;
  wire[0:0] or_898_nl;
  wire[0:0] mux_1276_nl;
  wire[0:0] mux_1275_nl;
  wire[0:0] or_891_nl;
  wire[0:0] nor_231_nl;
  wire[0:0] mux_1344_nl;
  wire[0:0] mux_1343_nl;
  wire[0:0] and_645_nl;
  wire[0:0] mux_1342_nl;
  wire[0:0] nor_1072_nl;
  wire[0:0] mux_1341_nl;
  wire[0:0] nor_1074_nl;
  wire[0:0] mux_1340_nl;
  wire[0:0] nor_1075_nl;
  wire[0:0] mux_1339_nl;
  wire[0:0] or_989_nl;
  wire[0:0] or_988_nl;
  wire[0:0] mux_1338_nl;
  wire[0:0] nor_1076_nl;
  wire[0:0] nor_1077_nl;
  wire[0:0] mux_1337_nl;
  wire[0:0] mux_1336_nl;
  wire[0:0] nor_1078_nl;
  wire[0:0] mux_1335_nl;
  wire[0:0] nor_1079_nl;
  wire[0:0] mux_1334_nl;
  wire[0:0] or_980_nl;
  wire[0:0] or_978_nl;
  wire[0:0] nor_1080_nl;
  wire[0:0] mux_1333_nl;
  wire[0:0] nor_1081_nl;
  wire[0:0] and_646_nl;
  wire[0:0] mux_1332_nl;
  wire[0:0] nor_1082_nl;
  wire[0:0] mux_1331_nl;
  wire[0:0] nor_1083_nl;
  wire[0:0] mux_1330_nl;
  wire[0:0] mux_1329_nl;
  wire[0:0] nor_1085_nl;
  wire[0:0] mux_1328_nl;
  wire[0:0] mux_1327_nl;
  wire[0:0] or_969_nl;
  wire[0:0] or_968_nl;
  wire[0:0] mux_1326_nl;
  wire[0:0] or_967_nl;
  wire[0:0] or_965_nl;
  wire[0:0] mux_1325_nl;
  wire[0:0] mux_1324_nl;
  wire[0:0] nor_1086_nl;
  wire[0:0] nor_1087_nl;
  wire[0:0] mux_1323_nl;
  wire[0:0] or_960_nl;
  wire[0:0] mux_1322_nl;
  wire[0:0] nor_1088_nl;
  wire[0:0] nor_1089_nl;
  wire[0:0] mux_1321_nl;
  wire[0:0] nor_1090_nl;
  wire[0:0] mux_1320_nl;
  wire[0:0] mux_1319_nl;
  wire[0:0] or_954_nl;
  wire[0:0] mux_1318_nl;
  wire[0:0] or_952_nl;
  wire[0:0] or_949_nl;
  wire[0:0] mux_1317_nl;
  wire[0:0] and_647_nl;
  wire[0:0] mux_1316_nl;
  wire[0:0] nor_1091_nl;
  wire[0:0] mux_1315_nl;
  wire[0:0] nor_1092_nl;
  wire[0:0] nor_1093_nl;
  wire[0:0] nor_1094_nl;
  wire[0:0] mux_1386_nl;
  wire[0:0] mux_1385_nl;
  wire[0:0] mux_1384_nl;
  wire[0:0] mux_1383_nl;
  wire[0:0] mux_1382_nl;
  wire[0:0] mux_1381_nl;
  wire[0:0] or_1050_nl;
  wire[0:0] mux_1379_nl;
  wire[0:0] mux_1378_nl;
  wire[0:0] or_1041_nl;
  wire[0:0] mux_1377_nl;
  wire[0:0] mux_1373_nl;
  wire[0:0] mux_1372_nl;
  wire[0:0] mux_1371_nl;
  wire[0:0] mux_1370_nl;
  wire[0:0] or_1031_nl;
  wire[0:0] mux_1369_nl;
  wire[0:0] mux_1367_nl;
  wire[0:0] mux_1366_nl;
  wire[0:0] mux_1365_nl;
  wire[0:0] mux_1364_nl;
  wire[0:0] or_1028_nl;
  wire[0:0] mux_1363_nl;
  wire[0:0] mux_1362_nl;
  wire[0:0] or_1023_nl;
  wire[0:0] mux_1360_nl;
  wire[0:0] mux_1359_nl;
  wire[0:0] mux_1358_nl;
  wire[0:0] or_1020_nl;
  wire[0:0] mux_1357_nl;
  wire[0:0] or_1018_nl;
  wire[0:0] or_1014_nl;
  wire[0:0] mux_1352_nl;
  wire[0:0] mux_1351_nl;
  wire[0:0] or_1007_nl;
  wire[0:0] or_1006_nl;
  wire[0:0] mux_1348_nl;
  wire[0:0] mux_1347_nl;
  wire[0:0] mux_1346_nl;
  wire[0:0] or_999_nl;
  wire[0:0] or_996_nl;
  wire[0:0] or_995_nl;
  wire[0:0] mux_1416_nl;
  wire[0:0] mux_1415_nl;
  wire[0:0] and_642_nl;
  wire[0:0] mux_1414_nl;
  wire[0:0] nor_1047_nl;
  wire[0:0] mux_1413_nl;
  wire[0:0] nor_1049_nl;
  wire[0:0] mux_1412_nl;
  wire[0:0] nor_1050_nl;
  wire[0:0] mux_1411_nl;
  wire[0:0] or_1096_nl;
  wire[0:0] or_1095_nl;
  wire[0:0] mux_1410_nl;
  wire[0:0] nor_1051_nl;
  wire[0:0] nor_1052_nl;
  wire[0:0] mux_1409_nl;
  wire[0:0] mux_1408_nl;
  wire[0:0] nor_1053_nl;
  wire[0:0] mux_1407_nl;
  wire[0:0] nor_1054_nl;
  wire[0:0] mux_1406_nl;
  wire[0:0] or_1087_nl;
  wire[0:0] or_1085_nl;
  wire[0:0] nor_1055_nl;
  wire[0:0] mux_1405_nl;
  wire[0:0] nor_1056_nl;
  wire[0:0] and_643_nl;
  wire[0:0] mux_1404_nl;
  wire[0:0] nor_1057_nl;
  wire[0:0] mux_1403_nl;
  wire[0:0] nor_1058_nl;
  wire[0:0] mux_1402_nl;
  wire[0:0] mux_1401_nl;
  wire[0:0] nor_1060_nl;
  wire[0:0] mux_1400_nl;
  wire[0:0] mux_1399_nl;
  wire[0:0] or_1076_nl;
  wire[0:0] or_1075_nl;
  wire[0:0] mux_1398_nl;
  wire[0:0] or_1074_nl;
  wire[0:0] or_1072_nl;
  wire[0:0] mux_1397_nl;
  wire[0:0] mux_1396_nl;
  wire[0:0] nor_1061_nl;
  wire[0:0] nor_1062_nl;
  wire[0:0] mux_1395_nl;
  wire[0:0] or_1067_nl;
  wire[0:0] mux_1394_nl;
  wire[0:0] nor_1063_nl;
  wire[0:0] nor_1064_nl;
  wire[0:0] mux_1393_nl;
  wire[0:0] nor_1065_nl;
  wire[0:0] mux_1392_nl;
  wire[0:0] mux_1391_nl;
  wire[0:0] or_1061_nl;
  wire[0:0] mux_1390_nl;
  wire[0:0] or_1059_nl;
  wire[0:0] or_1056_nl;
  wire[0:0] mux_1389_nl;
  wire[0:0] and_644_nl;
  wire[0:0] mux_1388_nl;
  wire[0:0] nor_1066_nl;
  wire[0:0] mux_1387_nl;
  wire[0:0] nor_1067_nl;
  wire[0:0] nor_1068_nl;
  wire[0:0] nor_1069_nl;
  wire[0:0] mux_1458_nl;
  wire[0:0] mux_1457_nl;
  wire[0:0] mux_1456_nl;
  wire[0:0] mux_1455_nl;
  wire[0:0] or_1156_nl;
  wire[0:0] mux_1454_nl;
  wire[0:0] or_1154_nl;
  wire[0:0] or_1153_nl;
  wire[0:0] mux_1453_nl;
  wire[0:0] mux_1452_nl;
  wire[0:0] or_1152_nl;
  wire[0:0] or_1151_nl;
  wire[0:0] mux_1451_nl;
  wire[0:0] mux_1450_nl;
  wire[0:0] mux_1449_nl;
  wire[0:0] or_1150_nl;
  wire[0:0] or_1149_nl;
  wire[0:0] mux_1448_nl;
  wire[0:0] mux_1447_nl;
  wire[0:0] mux_1446_nl;
  wire[0:0] mux_1445_nl;
  wire[0:0] mux_1444_nl;
  wire[0:0] or_1148_nl;
  wire[0:0] mux_1442_nl;
  wire[0:0] mux_1441_nl;
  wire[0:0] or_1139_nl;
  wire[0:0] mux_1439_nl;
  wire[0:0] mux_1432_nl;
  wire[0:0] mux_1431_nl;
  wire[0:0] mux_1430_nl;
  wire[0:0] mux_1429_nl;
  wire[0:0] or_1120_nl;
  wire[0:0] mux_1428_nl;
  wire[0:0] mux_1424_nl;
  wire[0:0] mux_1423_nl;
  wire[0:0] mux_1422_nl;
  wire[0:0] mux_1421_nl;
  wire[0:0] or_1111_nl;
  wire[0:0] mux_1420_nl;
  wire[0:0] mux_1419_nl;
  wire[0:0] or_1104_nl;
  wire[0:0] nor_238_nl;
  wire[0:0] mux_1488_nl;
  wire[0:0] mux_1487_nl;
  wire[0:0] and_639_nl;
  wire[0:0] mux_1486_nl;
  wire[0:0] nor_1022_nl;
  wire[0:0] mux_1485_nl;
  wire[0:0] nor_1024_nl;
  wire[0:0] mux_1484_nl;
  wire[0:0] nor_1025_nl;
  wire[0:0] mux_1483_nl;
  wire[0:0] or_1202_nl;
  wire[0:0] or_1201_nl;
  wire[0:0] mux_1482_nl;
  wire[0:0] nor_1026_nl;
  wire[0:0] nor_1027_nl;
  wire[0:0] mux_1481_nl;
  wire[0:0] mux_1480_nl;
  wire[0:0] nor_1028_nl;
  wire[0:0] mux_1479_nl;
  wire[0:0] nor_1029_nl;
  wire[0:0] mux_1478_nl;
  wire[0:0] or_1193_nl;
  wire[0:0] or_1191_nl;
  wire[0:0] nor_1030_nl;
  wire[0:0] mux_1477_nl;
  wire[0:0] nor_1031_nl;
  wire[0:0] and_640_nl;
  wire[0:0] mux_1476_nl;
  wire[0:0] nor_1032_nl;
  wire[0:0] mux_1475_nl;
  wire[0:0] nor_1033_nl;
  wire[0:0] mux_1474_nl;
  wire[0:0] mux_1473_nl;
  wire[0:0] nor_1035_nl;
  wire[0:0] mux_1472_nl;
  wire[0:0] mux_1471_nl;
  wire[0:0] or_1182_nl;
  wire[0:0] or_1181_nl;
  wire[0:0] mux_1470_nl;
  wire[0:0] or_1180_nl;
  wire[0:0] or_1178_nl;
  wire[0:0] mux_1469_nl;
  wire[0:0] mux_1468_nl;
  wire[0:0] nor_1036_nl;
  wire[0:0] nor_1037_nl;
  wire[0:0] mux_1467_nl;
  wire[0:0] or_1173_nl;
  wire[0:0] mux_1466_nl;
  wire[0:0] nor_1038_nl;
  wire[0:0] nor_1039_nl;
  wire[0:0] mux_1465_nl;
  wire[0:0] nor_1040_nl;
  wire[0:0] mux_1464_nl;
  wire[0:0] mux_1463_nl;
  wire[0:0] or_1167_nl;
  wire[0:0] mux_1462_nl;
  wire[0:0] or_1165_nl;
  wire[0:0] or_1162_nl;
  wire[0:0] mux_1461_nl;
  wire[0:0] and_641_nl;
  wire[0:0] mux_1460_nl;
  wire[0:0] nor_1041_nl;
  wire[0:0] mux_1459_nl;
  wire[0:0] nor_1042_nl;
  wire[0:0] nor_1043_nl;
  wire[0:0] nor_1044_nl;
  wire[0:0] mux_1530_nl;
  wire[0:0] mux_1529_nl;
  wire[0:0] mux_1528_nl;
  wire[0:0] mux_1527_nl;
  wire[0:0] mux_1526_nl;
  wire[0:0] mux_1525_nl;
  wire[0:0] or_1263_nl;
  wire[0:0] mux_1523_nl;
  wire[0:0] mux_1522_nl;
  wire[0:0] or_1254_nl;
  wire[0:0] mux_1521_nl;
  wire[0:0] mux_1517_nl;
  wire[0:0] mux_1516_nl;
  wire[0:0] mux_1515_nl;
  wire[0:0] mux_1514_nl;
  wire[0:0] or_1244_nl;
  wire[0:0] mux_1513_nl;
  wire[0:0] mux_1511_nl;
  wire[0:0] mux_1510_nl;
  wire[0:0] mux_1509_nl;
  wire[0:0] mux_1508_nl;
  wire[0:0] or_1241_nl;
  wire[0:0] mux_1507_nl;
  wire[0:0] mux_1506_nl;
  wire[0:0] or_1236_nl;
  wire[0:0] mux_1504_nl;
  wire[0:0] mux_1503_nl;
  wire[0:0] mux_1502_nl;
  wire[0:0] or_1233_nl;
  wire[0:0] mux_1501_nl;
  wire[0:0] or_1231_nl;
  wire[0:0] or_1227_nl;
  wire[0:0] mux_1496_nl;
  wire[0:0] mux_1495_nl;
  wire[0:0] or_1220_nl;
  wire[0:0] or_1219_nl;
  wire[0:0] mux_1492_nl;
  wire[0:0] mux_1491_nl;
  wire[0:0] mux_1490_nl;
  wire[0:0] or_1212_nl;
  wire[0:0] or_1209_nl;
  wire[0:0] or_1208_nl;
  wire[0:0] mux_1560_nl;
  wire[0:0] mux_1559_nl;
  wire[0:0] and_636_nl;
  wire[0:0] mux_1558_nl;
  wire[0:0] nor_997_nl;
  wire[0:0] mux_1557_nl;
  wire[0:0] nor_999_nl;
  wire[0:0] mux_1556_nl;
  wire[0:0] nor_1000_nl;
  wire[0:0] mux_1555_nl;
  wire[0:0] or_1309_nl;
  wire[0:0] or_1308_nl;
  wire[0:0] mux_1554_nl;
  wire[0:0] nor_1001_nl;
  wire[0:0] nor_1002_nl;
  wire[0:0] mux_1553_nl;
  wire[0:0] mux_1552_nl;
  wire[0:0] nor_1003_nl;
  wire[0:0] mux_1551_nl;
  wire[0:0] nor_1004_nl;
  wire[0:0] mux_1550_nl;
  wire[0:0] or_1300_nl;
  wire[0:0] or_1298_nl;
  wire[0:0] nor_1005_nl;
  wire[0:0] mux_1549_nl;
  wire[0:0] nor_1006_nl;
  wire[0:0] and_637_nl;
  wire[0:0] mux_1548_nl;
  wire[0:0] nor_1007_nl;
  wire[0:0] mux_1547_nl;
  wire[0:0] nor_1008_nl;
  wire[0:0] mux_1546_nl;
  wire[0:0] mux_1545_nl;
  wire[0:0] nor_1010_nl;
  wire[0:0] mux_1544_nl;
  wire[0:0] mux_1543_nl;
  wire[0:0] or_1289_nl;
  wire[0:0] or_1288_nl;
  wire[0:0] mux_1542_nl;
  wire[0:0] or_1287_nl;
  wire[0:0] or_1285_nl;
  wire[0:0] mux_1541_nl;
  wire[0:0] mux_1540_nl;
  wire[0:0] nor_1011_nl;
  wire[0:0] nor_1012_nl;
  wire[0:0] mux_1539_nl;
  wire[0:0] or_1280_nl;
  wire[0:0] mux_1538_nl;
  wire[0:0] nor_1013_nl;
  wire[0:0] nor_1014_nl;
  wire[0:0] mux_1537_nl;
  wire[0:0] nor_1015_nl;
  wire[0:0] mux_1536_nl;
  wire[0:0] mux_1535_nl;
  wire[0:0] or_1274_nl;
  wire[0:0] mux_1534_nl;
  wire[0:0] or_1272_nl;
  wire[0:0] or_1269_nl;
  wire[0:0] mux_1533_nl;
  wire[0:0] and_638_nl;
  wire[0:0] mux_1532_nl;
  wire[0:0] nor_1016_nl;
  wire[0:0] mux_1531_nl;
  wire[0:0] nor_1017_nl;
  wire[0:0] nor_1018_nl;
  wire[0:0] nor_1019_nl;
  wire[0:0] mux_1602_nl;
  wire[0:0] mux_1601_nl;
  wire[0:0] mux_1600_nl;
  wire[0:0] mux_1599_nl;
  wire[0:0] or_1369_nl;
  wire[0:0] mux_1598_nl;
  wire[0:0] or_1367_nl;
  wire[0:0] or_1366_nl;
  wire[0:0] mux_1597_nl;
  wire[0:0] mux_1596_nl;
  wire[0:0] nand_336_nl;
  wire[0:0] or_1364_nl;
  wire[0:0] mux_1595_nl;
  wire[0:0] mux_1594_nl;
  wire[0:0] mux_1593_nl;
  wire[0:0] or_1363_nl;
  wire[0:0] or_1362_nl;
  wire[0:0] mux_1592_nl;
  wire[0:0] mux_1591_nl;
  wire[0:0] mux_1590_nl;
  wire[0:0] mux_1589_nl;
  wire[0:0] mux_1588_nl;
  wire[0:0] or_1361_nl;
  wire[0:0] mux_1586_nl;
  wire[0:0] mux_1585_nl;
  wire[0:0] or_1352_nl;
  wire[0:0] mux_1583_nl;
  wire[0:0] mux_1576_nl;
  wire[0:0] mux_1575_nl;
  wire[0:0] mux_1574_nl;
  wire[0:0] mux_1573_nl;
  wire[0:0] nand_338_nl;
  wire[0:0] mux_1572_nl;
  wire[0:0] mux_1568_nl;
  wire[0:0] mux_1567_nl;
  wire[0:0] mux_1566_nl;
  wire[0:0] mux_1565_nl;
  wire[0:0] or_1324_nl;
  wire[0:0] mux_1564_nl;
  wire[0:0] mux_1563_nl;
  wire[0:0] or_1317_nl;
  wire[0:0] and_635_nl;
  wire[0:0] mux_1632_nl;
  wire[0:0] mux_1631_nl;
  wire[0:0] and_630_nl;
  wire[0:0] mux_1630_nl;
  wire[0:0] nor_974_nl;
  wire[0:0] mux_1629_nl;
  wire[0:0] nor_976_nl;
  wire[0:0] mux_1628_nl;
  wire[0:0] nor_977_nl;
  wire[0:0] mux_1627_nl;
  wire[0:0] nand_333_nl;
  wire[0:0] or_1414_nl;
  wire[0:0] mux_1626_nl;
  wire[0:0] nor_978_nl;
  wire[0:0] nor_979_nl;
  wire[0:0] mux_1625_nl;
  wire[0:0] mux_1624_nl;
  wire[0:0] and_631_nl;
  wire[0:0] mux_1623_nl;
  wire[0:0] nor_980_nl;
  wire[0:0] mux_1622_nl;
  wire[0:0] or_1406_nl;
  wire[0:0] or_1404_nl;
  wire[0:0] nor_981_nl;
  wire[0:0] mux_1621_nl;
  wire[0:0] nor_982_nl;
  wire[0:0] and_632_nl;
  wire[0:0] mux_1620_nl;
  wire[0:0] and_828_nl;
  wire[0:0] mux_1619_nl;
  wire[0:0] nor_984_nl;
  wire[0:0] mux_1618_nl;
  wire[0:0] mux_1617_nl;
  wire[0:0] nor_986_nl;
  wire[0:0] mux_1616_nl;
  wire[0:0] mux_1615_nl;
  wire[0:0] or_1395_nl;
  wire[0:0] or_1394_nl;
  wire[0:0] mux_1614_nl;
  wire[0:0] or_1393_nl;
  wire[0:0] or_1391_nl;
  wire[0:0] mux_1613_nl;
  wire[0:0] mux_1612_nl;
  wire[0:0] nor_987_nl;
  wire[0:0] nor_988_nl;
  wire[0:0] mux_1611_nl;
  wire[0:0] or_1386_nl;
  wire[0:0] mux_1610_nl;
  wire[0:0] nor_989_nl;
  wire[0:0] nor_990_nl;
  wire[0:0] mux_1609_nl;
  wire[0:0] nor_991_nl;
  wire[0:0] mux_1608_nl;
  wire[0:0] mux_1607_nl;
  wire[0:0] nand_417_nl;
  wire[0:0] mux_1606_nl;
  wire[0:0] or_1378_nl;
  wire[0:0] or_1375_nl;
  wire[0:0] mux_1605_nl;
  wire[0:0] and_633_nl;
  wire[0:0] mux_1604_nl;
  wire[0:0] nor_992_nl;
  wire[0:0] mux_1603_nl;
  wire[0:0] and_634_nl;
  wire[0:0] nor_993_nl;
  wire[0:0] nor_994_nl;
  wire[0:0] mux_1674_nl;
  wire[0:0] mux_1673_nl;
  wire[0:0] mux_1672_nl;
  wire[0:0] mux_1671_nl;
  wire[0:0] mux_1670_nl;
  wire[0:0] mux_1669_nl;
  wire[0:0] or_1476_nl;
  wire[0:0] mux_1667_nl;
  wire[0:0] mux_1666_nl;
  wire[0:0] or_1467_nl;
  wire[0:0] mux_1665_nl;
  wire[0:0] mux_1661_nl;
  wire[0:0] mux_1660_nl;
  wire[0:0] mux_1659_nl;
  wire[0:0] mux_1658_nl;
  wire[0:0] or_1457_nl;
  wire[0:0] mux_1657_nl;
  wire[0:0] mux_1655_nl;
  wire[0:0] mux_1654_nl;
  wire[0:0] mux_1653_nl;
  wire[0:0] mux_1652_nl;
  wire[0:0] or_1454_nl;
  wire[0:0] mux_1651_nl;
  wire[0:0] mux_1650_nl;
  wire[0:0] or_1449_nl;
  wire[0:0] mux_1648_nl;
  wire[0:0] mux_1647_nl;
  wire[0:0] mux_1646_nl;
  wire[0:0] or_1446_nl;
  wire[0:0] mux_1645_nl;
  wire[0:0] or_1444_nl;
  wire[0:0] or_1440_nl;
  wire[0:0] mux_1640_nl;
  wire[0:0] mux_1639_nl;
  wire[0:0] or_1433_nl;
  wire[0:0] or_1432_nl;
  wire[0:0] mux_1636_nl;
  wire[0:0] mux_1635_nl;
  wire[0:0] mux_1634_nl;
  wire[0:0] or_1425_nl;
  wire[0:0] or_1422_nl;
  wire[0:0] or_1421_nl;
  wire[0:0] mux_1704_nl;
  wire[0:0] mux_1703_nl;
  wire[0:0] and_627_nl;
  wire[0:0] mux_1702_nl;
  wire[0:0] nor_949_nl;
  wire[0:0] mux_1701_nl;
  wire[0:0] nor_951_nl;
  wire[0:0] mux_1700_nl;
  wire[0:0] nor_952_nl;
  wire[0:0] mux_1699_nl;
  wire[0:0] or_1522_nl;
  wire[0:0] or_1521_nl;
  wire[0:0] mux_1698_nl;
  wire[0:0] nor_953_nl;
  wire[0:0] nor_954_nl;
  wire[0:0] mux_1697_nl;
  wire[0:0] mux_1696_nl;
  wire[0:0] nor_955_nl;
  wire[0:0] mux_1695_nl;
  wire[0:0] nor_956_nl;
  wire[0:0] mux_1694_nl;
  wire[0:0] or_1513_nl;
  wire[0:0] or_1511_nl;
  wire[0:0] nor_957_nl;
  wire[0:0] mux_1693_nl;
  wire[0:0] nor_958_nl;
  wire[0:0] and_628_nl;
  wire[0:0] mux_1692_nl;
  wire[0:0] nor_959_nl;
  wire[0:0] mux_1691_nl;
  wire[0:0] nor_960_nl;
  wire[0:0] mux_1690_nl;
  wire[0:0] mux_1689_nl;
  wire[0:0] nor_962_nl;
  wire[0:0] mux_1688_nl;
  wire[0:0] mux_1687_nl;
  wire[0:0] or_1502_nl;
  wire[0:0] or_1501_nl;
  wire[0:0] mux_1686_nl;
  wire[0:0] or_1500_nl;
  wire[0:0] or_1498_nl;
  wire[0:0] mux_1685_nl;
  wire[0:0] mux_1684_nl;
  wire[0:0] nor_963_nl;
  wire[0:0] nor_964_nl;
  wire[0:0] mux_1683_nl;
  wire[0:0] or_1493_nl;
  wire[0:0] mux_1682_nl;
  wire[0:0] nor_965_nl;
  wire[0:0] nor_966_nl;
  wire[0:0] mux_1681_nl;
  wire[0:0] nor_967_nl;
  wire[0:0] mux_1680_nl;
  wire[0:0] mux_1679_nl;
  wire[0:0] or_1487_nl;
  wire[0:0] mux_1678_nl;
  wire[0:0] or_1485_nl;
  wire[0:0] or_1482_nl;
  wire[0:0] mux_1677_nl;
  wire[0:0] and_629_nl;
  wire[0:0] mux_1676_nl;
  wire[0:0] nor_968_nl;
  wire[0:0] mux_1675_nl;
  wire[0:0] nor_969_nl;
  wire[0:0] nor_970_nl;
  wire[0:0] nor_971_nl;
  wire[0:0] mux_1746_nl;
  wire[0:0] mux_1745_nl;
  wire[0:0] mux_1744_nl;
  wire[0:0] mux_1743_nl;
  wire[0:0] or_1582_nl;
  wire[0:0] mux_1742_nl;
  wire[0:0] or_1580_nl;
  wire[0:0] or_1579_nl;
  wire[0:0] mux_1741_nl;
  wire[0:0] mux_1740_nl;
  wire[0:0] or_1578_nl;
  wire[0:0] or_1577_nl;
  wire[0:0] mux_1739_nl;
  wire[0:0] mux_1738_nl;
  wire[0:0] mux_1737_nl;
  wire[0:0] or_1576_nl;
  wire[0:0] or_1575_nl;
  wire[0:0] mux_1736_nl;
  wire[0:0] mux_1735_nl;
  wire[0:0] mux_1734_nl;
  wire[0:0] mux_1733_nl;
  wire[0:0] mux_1732_nl;
  wire[0:0] or_1574_nl;
  wire[0:0] mux_1730_nl;
  wire[0:0] mux_1729_nl;
  wire[0:0] or_1565_nl;
  wire[0:0] mux_1727_nl;
  wire[0:0] mux_1720_nl;
  wire[0:0] mux_1719_nl;
  wire[0:0] mux_1718_nl;
  wire[0:0] mux_1717_nl;
  wire[0:0] or_1546_nl;
  wire[0:0] mux_1716_nl;
  wire[0:0] mux_1712_nl;
  wire[0:0] mux_1711_nl;
  wire[0:0] mux_1710_nl;
  wire[0:0] mux_1709_nl;
  wire[0:0] or_1537_nl;
  wire[0:0] mux_1708_nl;
  wire[0:0] mux_1707_nl;
  wire[0:0] or_1530_nl;
  wire[0:0] nor_252_nl;
  wire[0:0] mux_1776_nl;
  wire[0:0] mux_1775_nl;
  wire[0:0] and_624_nl;
  wire[0:0] mux_1774_nl;
  wire[0:0] nor_924_nl;
  wire[0:0] mux_1773_nl;
  wire[0:0] nor_926_nl;
  wire[0:0] mux_1772_nl;
  wire[0:0] nor_927_nl;
  wire[0:0] mux_1771_nl;
  wire[0:0] or_1628_nl;
  wire[0:0] or_1627_nl;
  wire[0:0] mux_1770_nl;
  wire[0:0] nor_928_nl;
  wire[0:0] nor_929_nl;
  wire[0:0] mux_1769_nl;
  wire[0:0] mux_1768_nl;
  wire[0:0] nor_930_nl;
  wire[0:0] mux_1767_nl;
  wire[0:0] nor_931_nl;
  wire[0:0] mux_1766_nl;
  wire[0:0] or_1619_nl;
  wire[0:0] or_1617_nl;
  wire[0:0] nor_932_nl;
  wire[0:0] mux_1765_nl;
  wire[0:0] nor_933_nl;
  wire[0:0] and_625_nl;
  wire[0:0] mux_1764_nl;
  wire[0:0] nor_934_nl;
  wire[0:0] mux_1763_nl;
  wire[0:0] nor_935_nl;
  wire[0:0] mux_1762_nl;
  wire[0:0] mux_1761_nl;
  wire[0:0] nor_937_nl;
  wire[0:0] mux_1760_nl;
  wire[0:0] mux_1759_nl;
  wire[0:0] or_1608_nl;
  wire[0:0] or_1607_nl;
  wire[0:0] mux_1758_nl;
  wire[0:0] or_1606_nl;
  wire[0:0] or_1604_nl;
  wire[0:0] mux_1757_nl;
  wire[0:0] mux_1756_nl;
  wire[0:0] nor_938_nl;
  wire[0:0] nor_939_nl;
  wire[0:0] mux_1755_nl;
  wire[0:0] or_1599_nl;
  wire[0:0] mux_1754_nl;
  wire[0:0] nor_940_nl;
  wire[0:0] nor_941_nl;
  wire[0:0] mux_1753_nl;
  wire[0:0] nor_942_nl;
  wire[0:0] mux_1752_nl;
  wire[0:0] mux_1751_nl;
  wire[0:0] or_1593_nl;
  wire[0:0] mux_1750_nl;
  wire[0:0] or_1591_nl;
  wire[0:0] or_1588_nl;
  wire[0:0] mux_1749_nl;
  wire[0:0] and_626_nl;
  wire[0:0] mux_1748_nl;
  wire[0:0] nor_943_nl;
  wire[0:0] mux_1747_nl;
  wire[0:0] nor_944_nl;
  wire[0:0] nor_945_nl;
  wire[0:0] nor_946_nl;
  wire[0:0] mux_1818_nl;
  wire[0:0] mux_1817_nl;
  wire[0:0] mux_1816_nl;
  wire[0:0] mux_1815_nl;
  wire[0:0] mux_1814_nl;
  wire[0:0] mux_1813_nl;
  wire[0:0] or_1689_nl;
  wire[0:0] mux_1811_nl;
  wire[0:0] mux_1810_nl;
  wire[0:0] or_1680_nl;
  wire[0:0] mux_1809_nl;
  wire[0:0] mux_1805_nl;
  wire[0:0] mux_1804_nl;
  wire[0:0] mux_1803_nl;
  wire[0:0] mux_1802_nl;
  wire[0:0] or_1670_nl;
  wire[0:0] mux_1801_nl;
  wire[0:0] mux_1799_nl;
  wire[0:0] mux_1798_nl;
  wire[0:0] mux_1797_nl;
  wire[0:0] mux_1796_nl;
  wire[0:0] or_1667_nl;
  wire[0:0] mux_1795_nl;
  wire[0:0] mux_1794_nl;
  wire[0:0] or_1662_nl;
  wire[0:0] mux_1792_nl;
  wire[0:0] mux_1791_nl;
  wire[0:0] mux_1790_nl;
  wire[0:0] or_1659_nl;
  wire[0:0] mux_1789_nl;
  wire[0:0] or_1657_nl;
  wire[0:0] or_1653_nl;
  wire[0:0] mux_1784_nl;
  wire[0:0] mux_1783_nl;
  wire[0:0] or_1646_nl;
  wire[0:0] or_1645_nl;
  wire[0:0] mux_1780_nl;
  wire[0:0] mux_1779_nl;
  wire[0:0] mux_1778_nl;
  wire[0:0] or_1638_nl;
  wire[0:0] or_1635_nl;
  wire[0:0] or_1634_nl;
  wire[0:0] mux_1848_nl;
  wire[0:0] mux_1847_nl;
  wire[0:0] and_621_nl;
  wire[0:0] mux_1846_nl;
  wire[0:0] nor_899_nl;
  wire[0:0] mux_1845_nl;
  wire[0:0] nor_901_nl;
  wire[0:0] mux_1844_nl;
  wire[0:0] nor_902_nl;
  wire[0:0] mux_1843_nl;
  wire[0:0] or_1735_nl;
  wire[0:0] or_1734_nl;
  wire[0:0] mux_1842_nl;
  wire[0:0] nor_903_nl;
  wire[0:0] nor_904_nl;
  wire[0:0] mux_1841_nl;
  wire[0:0] mux_1840_nl;
  wire[0:0] nor_905_nl;
  wire[0:0] mux_1839_nl;
  wire[0:0] nor_906_nl;
  wire[0:0] mux_1838_nl;
  wire[0:0] or_1726_nl;
  wire[0:0] or_1724_nl;
  wire[0:0] nor_907_nl;
  wire[0:0] mux_1837_nl;
  wire[0:0] nor_908_nl;
  wire[0:0] and_622_nl;
  wire[0:0] mux_1836_nl;
  wire[0:0] nor_909_nl;
  wire[0:0] mux_1835_nl;
  wire[0:0] nor_910_nl;
  wire[0:0] mux_1834_nl;
  wire[0:0] mux_1833_nl;
  wire[0:0] nor_912_nl;
  wire[0:0] mux_1832_nl;
  wire[0:0] mux_1831_nl;
  wire[0:0] or_1715_nl;
  wire[0:0] or_1714_nl;
  wire[0:0] mux_1830_nl;
  wire[0:0] or_1713_nl;
  wire[0:0] or_1711_nl;
  wire[0:0] mux_1829_nl;
  wire[0:0] mux_1828_nl;
  wire[0:0] nor_913_nl;
  wire[0:0] nor_914_nl;
  wire[0:0] mux_1827_nl;
  wire[0:0] or_1706_nl;
  wire[0:0] mux_1826_nl;
  wire[0:0] nor_915_nl;
  wire[0:0] nor_916_nl;
  wire[0:0] mux_1825_nl;
  wire[0:0] nor_917_nl;
  wire[0:0] mux_1824_nl;
  wire[0:0] mux_1823_nl;
  wire[0:0] or_1700_nl;
  wire[0:0] mux_1822_nl;
  wire[0:0] or_1698_nl;
  wire[0:0] or_1695_nl;
  wire[0:0] mux_1821_nl;
  wire[0:0] and_623_nl;
  wire[0:0] mux_1820_nl;
  wire[0:0] nor_918_nl;
  wire[0:0] mux_1819_nl;
  wire[0:0] nor_919_nl;
  wire[0:0] nor_920_nl;
  wire[0:0] nor_921_nl;
  wire[0:0] mux_1890_nl;
  wire[0:0] mux_1889_nl;
  wire[0:0] mux_1888_nl;
  wire[0:0] mux_1887_nl;
  wire[0:0] or_1795_nl;
  wire[0:0] mux_1886_nl;
  wire[0:0] or_1793_nl;
  wire[0:0] or_1792_nl;
  wire[0:0] mux_1885_nl;
  wire[0:0] mux_1884_nl;
  wire[0:0] nand_319_nl;
  wire[0:0] or_1790_nl;
  wire[0:0] mux_1883_nl;
  wire[0:0] mux_1882_nl;
  wire[0:0] mux_1881_nl;
  wire[0:0] or_1789_nl;
  wire[0:0] or_1788_nl;
  wire[0:0] mux_1880_nl;
  wire[0:0] mux_1879_nl;
  wire[0:0] mux_1878_nl;
  wire[0:0] mux_1877_nl;
  wire[0:0] mux_1876_nl;
  wire[0:0] or_1787_nl;
  wire[0:0] mux_1874_nl;
  wire[0:0] mux_1873_nl;
  wire[0:0] or_1778_nl;
  wire[0:0] mux_1871_nl;
  wire[0:0] mux_1864_nl;
  wire[0:0] mux_1863_nl;
  wire[0:0] mux_1862_nl;
  wire[0:0] mux_1861_nl;
  wire[0:0] nand_321_nl;
  wire[0:0] mux_1860_nl;
  wire[0:0] mux_1856_nl;
  wire[0:0] mux_1855_nl;
  wire[0:0] mux_1854_nl;
  wire[0:0] mux_1853_nl;
  wire[0:0] or_1750_nl;
  wire[0:0] mux_1852_nl;
  wire[0:0] mux_1851_nl;
  wire[0:0] or_1743_nl;
  wire[0:0] and_620_nl;
  wire[0:0] mux_1920_nl;
  wire[0:0] mux_1919_nl;
  wire[0:0] and_615_nl;
  wire[0:0] mux_1918_nl;
  wire[0:0] nor_876_nl;
  wire[0:0] mux_1917_nl;
  wire[0:0] nor_878_nl;
  wire[0:0] mux_1916_nl;
  wire[0:0] nor_879_nl;
  wire[0:0] mux_1915_nl;
  wire[0:0] nand_316_nl;
  wire[0:0] or_1840_nl;
  wire[0:0] mux_1914_nl;
  wire[0:0] nor_880_nl;
  wire[0:0] nor_881_nl;
  wire[0:0] mux_1913_nl;
  wire[0:0] mux_1912_nl;
  wire[0:0] and_616_nl;
  wire[0:0] mux_1911_nl;
  wire[0:0] nor_882_nl;
  wire[0:0] mux_1910_nl;
  wire[0:0] or_1832_nl;
  wire[0:0] or_1830_nl;
  wire[0:0] nor_883_nl;
  wire[0:0] mux_1909_nl;
  wire[0:0] nor_884_nl;
  wire[0:0] and_617_nl;
  wire[0:0] mux_1908_nl;
  wire[0:0] and_827_nl;
  wire[0:0] mux_1907_nl;
  wire[0:0] nor_886_nl;
  wire[0:0] mux_1906_nl;
  wire[0:0] mux_1905_nl;
  wire[0:0] nor_888_nl;
  wire[0:0] mux_1904_nl;
  wire[0:0] mux_1903_nl;
  wire[0:0] or_1821_nl;
  wire[0:0] or_1820_nl;
  wire[0:0] mux_1902_nl;
  wire[0:0] or_1819_nl;
  wire[0:0] or_1817_nl;
  wire[0:0] mux_1901_nl;
  wire[0:0] mux_1900_nl;
  wire[0:0] nor_889_nl;
  wire[0:0] nor_890_nl;
  wire[0:0] mux_1899_nl;
  wire[0:0] or_1812_nl;
  wire[0:0] mux_1898_nl;
  wire[0:0] nor_891_nl;
  wire[0:0] nor_892_nl;
  wire[0:0] mux_1897_nl;
  wire[0:0] nor_893_nl;
  wire[0:0] mux_1896_nl;
  wire[0:0] mux_1895_nl;
  wire[0:0] nand_415_nl;
  wire[0:0] mux_1894_nl;
  wire[0:0] or_1804_nl;
  wire[0:0] or_1801_nl;
  wire[0:0] mux_1893_nl;
  wire[0:0] and_618_nl;
  wire[0:0] mux_1892_nl;
  wire[0:0] nor_894_nl;
  wire[0:0] mux_1891_nl;
  wire[0:0] and_619_nl;
  wire[0:0] nor_895_nl;
  wire[0:0] nor_896_nl;
  wire[0:0] mux_1963_nl;
  wire[0:0] mux_1962_nl;
  wire[0:0] mux_1961_nl;
  wire[0:0] mux_1960_nl;
  wire[0:0] mux_1959_nl;
  wire[0:0] mux_1958_nl;
  wire[0:0] or_1905_nl;
  wire[0:0] or_1903_nl;
  wire[0:0] or_1902_nl;
  wire[0:0] mux_1957_nl;
  wire[0:0] nand_311_nl;
  wire[0:0] or_1900_nl;
  wire[0:0] mux_1956_nl;
  wire[0:0] mux_1955_nl;
  wire[0:0] mux_1954_nl;
  wire[0:0] or_1898_nl;
  wire[0:0] or_1896_nl;
  wire[0:0] mux_1953_nl;
  wire[0:0] or_1894_nl;
  wire[0:0] mux_1952_nl;
  wire[0:0] nand_437_nl;
  wire[0:0] mux_1951_nl;
  wire[0:0] or_1891_nl;
  wire[0:0] mux_1950_nl;
  wire[0:0] mux_1949_nl;
  wire[0:0] or_1890_nl;
  wire[0:0] mux_1948_nl;
  wire[0:0] or_1889_nl;
  wire[0:0] or_1888_nl;
  wire[0:0] mux_1947_nl;
  wire[0:0] mux_1946_nl;
  wire[0:0] mux_1945_nl;
  wire[0:0] mux_1944_nl;
  wire[0:0] or_1887_nl;
  wire[0:0] or_1886_nl;
  wire[0:0] mux_1943_nl;
  wire[0:0] or_1884_nl;
  wire[0:0] or_1883_nl;
  wire[0:0] mux_1942_nl;
  wire[0:0] mux_1941_nl;
  wire[0:0] mux_1940_nl;
  wire[0:0] or_1882_nl;
  wire[0:0] or_1881_nl;
  wire[0:0] mux_1939_nl;
  wire[0:0] mux_1938_nl;
  wire[0:0] mux_1937_nl;
  wire[0:0] or_1879_nl;
  wire[0:0] or_1876_nl;
  wire[0:0] or_1875_nl;
  wire[0:0] mux_1936_nl;
  wire[0:0] mux_1935_nl;
  wire[0:0] mux_1934_nl;
  wire[0:0] or_1873_nl;
  wire[0:0] mux_1933_nl;
  wire[0:0] mux_1932_nl;
  wire[0:0] or_1871_nl;
  wire[0:0] mux_1931_nl;
  wire[0:0] or_1867_nl;
  wire[0:0] mux_1930_nl;
  wire[0:0] or_1866_nl;
  wire[0:0] mux_1928_nl;
  wire[0:0] or_1862_nl;
  wire[0:0] mux_1924_nl;
  wire[0:0] mux_1923_nl;
  wire[0:0] or_1850_nl;
  wire[0:0] or_1848_nl;
  wire[0:0] or_1847_nl;
  wire[0:0] mux_1993_nl;
  wire[0:0] mux_1992_nl;
  wire[0:0] and_612_nl;
  wire[0:0] mux_1991_nl;
  wire[0:0] nor_849_nl;
  wire[0:0] mux_1990_nl;
  wire[0:0] nor_851_nl;
  wire[0:0] mux_1989_nl;
  wire[0:0] nor_852_nl;
  wire[0:0] mux_1988_nl;
  wire[0:0] or_1951_nl;
  wire[0:0] or_1950_nl;
  wire[0:0] mux_1987_nl;
  wire[0:0] nor_853_nl;
  wire[0:0] nor_854_nl;
  wire[0:0] mux_1986_nl;
  wire[0:0] mux_1985_nl;
  wire[0:0] nor_855_nl;
  wire[0:0] mux_1984_nl;
  wire[0:0] nor_856_nl;
  wire[0:0] mux_1983_nl;
  wire[0:0] or_1942_nl;
  wire[0:0] or_1940_nl;
  wire[0:0] nor_857_nl;
  wire[0:0] mux_1982_nl;
  wire[0:0] nor_858_nl;
  wire[0:0] and_613_nl;
  wire[0:0] mux_1981_nl;
  wire[0:0] nor_859_nl;
  wire[0:0] mux_1980_nl;
  wire[0:0] nor_860_nl;
  wire[0:0] mux_1979_nl;
  wire[0:0] mux_1978_nl;
  wire[0:0] nor_862_nl;
  wire[0:0] mux_1977_nl;
  wire[0:0] mux_1976_nl;
  wire[0:0] or_1931_nl;
  wire[0:0] or_1930_nl;
  wire[0:0] mux_1975_nl;
  wire[0:0] or_1929_nl;
  wire[0:0] or_1927_nl;
  wire[0:0] mux_1974_nl;
  wire[0:0] mux_1973_nl;
  wire[0:0] nor_863_nl;
  wire[0:0] nor_864_nl;
  wire[0:0] mux_1972_nl;
  wire[0:0] or_1922_nl;
  wire[0:0] mux_1971_nl;
  wire[0:0] nor_865_nl;
  wire[0:0] nor_866_nl;
  wire[0:0] mux_1970_nl;
  wire[0:0] nor_867_nl;
  wire[0:0] mux_1969_nl;
  wire[0:0] mux_1968_nl;
  wire[0:0] or_1916_nl;
  wire[0:0] mux_1967_nl;
  wire[0:0] or_1914_nl;
  wire[0:0] or_1911_nl;
  wire[0:0] mux_1966_nl;
  wire[0:0] and_614_nl;
  wire[0:0] mux_1965_nl;
  wire[0:0] nor_868_nl;
  wire[0:0] mux_1964_nl;
  wire[0:0] nor_869_nl;
  wire[0:0] nor_870_nl;
  wire[0:0] nor_871_nl;
  wire[0:0] mux_2035_nl;
  wire[0:0] mux_2034_nl;
  wire[0:0] mux_2033_nl;
  wire[0:0] mux_2032_nl;
  wire[0:0] or_2011_nl;
  wire[0:0] mux_2031_nl;
  wire[0:0] or_2009_nl;
  wire[0:0] or_2008_nl;
  wire[0:0] mux_2030_nl;
  wire[0:0] mux_2029_nl;
  wire[0:0] nand_305_nl;
  wire[0:0] or_2006_nl;
  wire[0:0] mux_2028_nl;
  wire[0:0] mux_2027_nl;
  wire[0:0] mux_2026_nl;
  wire[0:0] or_2005_nl;
  wire[0:0] or_2004_nl;
  wire[0:0] mux_2025_nl;
  wire[0:0] mux_2024_nl;
  wire[0:0] mux_2023_nl;
  wire[0:0] mux_2022_nl;
  wire[0:0] mux_2021_nl;
  wire[0:0] or_2003_nl;
  wire[0:0] mux_2019_nl;
  wire[0:0] mux_2018_nl;
  wire[0:0] or_1994_nl;
  wire[0:0] mux_2016_nl;
  wire[0:0] mux_2009_nl;
  wire[0:0] mux_2008_nl;
  wire[0:0] mux_2007_nl;
  wire[0:0] mux_2006_nl;
  wire[0:0] nand_307_nl;
  wire[0:0] mux_2005_nl;
  wire[0:0] mux_2001_nl;
  wire[0:0] mux_2000_nl;
  wire[0:0] mux_1999_nl;
  wire[0:0] mux_1998_nl;
  wire[0:0] or_1966_nl;
  wire[0:0] mux_1997_nl;
  wire[0:0] mux_1996_nl;
  wire[0:0] or_1959_nl;
  wire[0:0] and_611_nl;
  wire[0:0] mux_2065_nl;
  wire[0:0] mux_2064_nl;
  wire[0:0] and_606_nl;
  wire[0:0] mux_2063_nl;
  wire[0:0] nor_826_nl;
  wire[0:0] mux_2062_nl;
  wire[0:0] nor_828_nl;
  wire[0:0] mux_2061_nl;
  wire[0:0] nor_829_nl;
  wire[0:0] mux_2060_nl;
  wire[0:0] nand_302_nl;
  wire[0:0] or_2056_nl;
  wire[0:0] mux_2059_nl;
  wire[0:0] nor_830_nl;
  wire[0:0] nor_831_nl;
  wire[0:0] mux_2058_nl;
  wire[0:0] mux_2057_nl;
  wire[0:0] and_607_nl;
  wire[0:0] mux_2056_nl;
  wire[0:0] nor_832_nl;
  wire[0:0] mux_2055_nl;
  wire[0:0] or_2048_nl;
  wire[0:0] or_2046_nl;
  wire[0:0] nor_833_nl;
  wire[0:0] mux_2054_nl;
  wire[0:0] nor_834_nl;
  wire[0:0] and_608_nl;
  wire[0:0] mux_2053_nl;
  wire[0:0] and_826_nl;
  wire[0:0] mux_2052_nl;
  wire[0:0] nor_836_nl;
  wire[0:0] mux_2051_nl;
  wire[0:0] mux_2050_nl;
  wire[0:0] nor_838_nl;
  wire[0:0] mux_2049_nl;
  wire[0:0] mux_2048_nl;
  wire[0:0] or_2037_nl;
  wire[0:0] or_2036_nl;
  wire[0:0] mux_2047_nl;
  wire[0:0] or_2035_nl;
  wire[0:0] or_2033_nl;
  wire[0:0] mux_2046_nl;
  wire[0:0] mux_2045_nl;
  wire[0:0] nor_839_nl;
  wire[0:0] nor_840_nl;
  wire[0:0] mux_2044_nl;
  wire[0:0] or_2028_nl;
  wire[0:0] mux_2043_nl;
  wire[0:0] nor_841_nl;
  wire[0:0] nor_842_nl;
  wire[0:0] mux_2042_nl;
  wire[0:0] nor_843_nl;
  wire[0:0] mux_2041_nl;
  wire[0:0] mux_2040_nl;
  wire[0:0] nand_413_nl;
  wire[0:0] mux_2039_nl;
  wire[0:0] or_2020_nl;
  wire[0:0] or_2017_nl;
  wire[0:0] mux_2038_nl;
  wire[0:0] and_609_nl;
  wire[0:0] mux_2037_nl;
  wire[0:0] nor_844_nl;
  wire[0:0] mux_2036_nl;
  wire[0:0] and_610_nl;
  wire[0:0] nor_845_nl;
  wire[0:0] nor_846_nl;
  wire[0:0] mux_2107_nl;
  wire[0:0] mux_2106_nl;
  wire[0:0] mux_2105_nl;
  wire[0:0] mux_2104_nl;
  wire[0:0] mux_2103_nl;
  wire[0:0] mux_2102_nl;
  wire[0:0] or_2118_nl;
  wire[0:0] mux_2100_nl;
  wire[0:0] mux_2099_nl;
  wire[0:0] or_2109_nl;
  wire[0:0] mux_2098_nl;
  wire[0:0] mux_2094_nl;
  wire[0:0] mux_2093_nl;
  wire[0:0] mux_2092_nl;
  wire[0:0] mux_2091_nl;
  wire[0:0] nand_297_nl;
  wire[0:0] mux_2090_nl;
  wire[0:0] mux_2088_nl;
  wire[0:0] mux_2087_nl;
  wire[0:0] mux_2086_nl;
  wire[0:0] mux_2085_nl;
  wire[0:0] or_2096_nl;
  wire[0:0] mux_2084_nl;
  wire[0:0] mux_2083_nl;
  wire[0:0] or_2091_nl;
  wire[0:0] mux_2081_nl;
  wire[0:0] mux_2080_nl;
  wire[0:0] mux_2079_nl;
  wire[0:0] or_2088_nl;
  wire[0:0] mux_2078_nl;
  wire[0:0] or_2086_nl;
  wire[0:0] or_2082_nl;
  wire[0:0] mux_2073_nl;
  wire[0:0] mux_2072_nl;
  wire[0:0] nand_298_nl;
  wire[0:0] or_2074_nl;
  wire[0:0] mux_2069_nl;
  wire[0:0] mux_2068_nl;
  wire[0:0] mux_2067_nl;
  wire[0:0] or_2067_nl;
  wire[0:0] or_2064_nl;
  wire[0:0] nand_299_nl;
  wire[0:0] mux_2137_nl;
  wire[0:0] mux_2136_nl;
  wire[0:0] and_601_nl;
  wire[0:0] mux_2135_nl;
  wire[0:0] nor_803_nl;
  wire[0:0] mux_2134_nl;
  wire[0:0] nor_805_nl;
  wire[0:0] mux_2133_nl;
  wire[0:0] nor_806_nl;
  wire[0:0] mux_2132_nl;
  wire[0:0] nand_293_nl;
  wire[0:0] or_2163_nl;
  wire[0:0] mux_2131_nl;
  wire[0:0] nor_807_nl;
  wire[0:0] nor_808_nl;
  wire[0:0] mux_2130_nl;
  wire[0:0] mux_2129_nl;
  wire[0:0] and_602_nl;
  wire[0:0] mux_2128_nl;
  wire[0:0] nor_809_nl;
  wire[0:0] mux_2127_nl;
  wire[0:0] or_2155_nl;
  wire[0:0] or_2153_nl;
  wire[0:0] nor_810_nl;
  wire[0:0] mux_2126_nl;
  wire[0:0] nor_811_nl;
  wire[0:0] and_603_nl;
  wire[0:0] mux_2125_nl;
  wire[0:0] and_825_nl;
  wire[0:0] mux_2124_nl;
  wire[0:0] nor_813_nl;
  wire[0:0] mux_2123_nl;
  wire[0:0] mux_2122_nl;
  wire[0:0] nor_815_nl;
  wire[0:0] mux_2121_nl;
  wire[0:0] mux_2120_nl;
  wire[0:0] or_2144_nl;
  wire[0:0] or_2143_nl;
  wire[0:0] mux_2119_nl;
  wire[0:0] or_2142_nl;
  wire[0:0] or_2140_nl;
  wire[0:0] mux_2118_nl;
  wire[0:0] mux_2117_nl;
  wire[0:0] nor_816_nl;
  wire[0:0] nor_817_nl;
  wire[0:0] mux_2116_nl;
  wire[0:0] or_2135_nl;
  wire[0:0] mux_2115_nl;
  wire[0:0] nor_818_nl;
  wire[0:0] nor_819_nl;
  wire[0:0] mux_2114_nl;
  wire[0:0] nor_820_nl;
  wire[0:0] mux_2113_nl;
  wire[0:0] mux_2112_nl;
  wire[0:0] nand_411_nl;
  wire[0:0] mux_2111_nl;
  wire[0:0] or_2127_nl;
  wire[0:0] or_2124_nl;
  wire[0:0] mux_2110_nl;
  wire[0:0] and_604_nl;
  wire[0:0] mux_2109_nl;
  wire[0:0] nor_821_nl;
  wire[0:0] mux_2108_nl;
  wire[0:0] and_605_nl;
  wire[0:0] nor_822_nl;
  wire[0:0] nor_823_nl;
  wire[0:0] mux_2179_nl;
  wire[0:0] mux_2178_nl;
  wire[0:0] mux_2177_nl;
  wire[0:0] mux_2176_nl;
  wire[0:0] or_2224_nl;
  wire[0:0] mux_2175_nl;
  wire[0:0] or_2222_nl;
  wire[0:0] or_2221_nl;
  wire[0:0] mux_2174_nl;
  wire[0:0] mux_2173_nl;
  wire[0:0] nand_284_nl;
  wire[0:0] or_2219_nl;
  wire[0:0] mux_2172_nl;
  wire[0:0] mux_2171_nl;
  wire[0:0] mux_2170_nl;
  wire[0:0] or_2218_nl;
  wire[0:0] or_2217_nl;
  wire[0:0] mux_2169_nl;
  wire[0:0] mux_2168_nl;
  wire[0:0] mux_2167_nl;
  wire[0:0] mux_2166_nl;
  wire[0:0] mux_2165_nl;
  wire[0:0] nand_438_nl;
  wire[0:0] mux_2163_nl;
  wire[0:0] mux_2162_nl;
  wire[0:0] or_2207_nl;
  wire[0:0] mux_2160_nl;
  wire[0:0] mux_2153_nl;
  wire[0:0] mux_2152_nl;
  wire[0:0] mux_2151_nl;
  wire[0:0] mux_2150_nl;
  wire[0:0] nand_286_nl;
  wire[0:0] mux_2149_nl;
  wire[0:0] mux_2145_nl;
  wire[0:0] mux_2144_nl;
  wire[0:0] mux_2143_nl;
  wire[0:0] mux_2142_nl;
  wire[0:0] or_2179_nl;
  wire[0:0] mux_2141_nl;
  wire[0:0] mux_2140_nl;
  wire[0:0] or_2172_nl;
  wire[0:0] and_600_nl;
  wire[0:0] mux_2209_nl;
  wire[0:0] mux_2208_nl;
  wire[0:0] and_590_nl;
  wire[0:0] mux_2207_nl;
  wire[0:0] and_823_nl;
  wire[0:0] mux_2206_nl;
  wire[0:0] nor_786_nl;
  wire[0:0] mux_2205_nl;
  wire[0:0] nor_787_nl;
  wire[0:0] mux_2204_nl;
  wire[0:0] nand_269_nl;
  wire[0:0] or_2269_nl;
  wire[0:0] mux_2203_nl;
  wire[0:0] nor_788_nl;
  wire[0:0] nor_789_nl;
  wire[0:0] mux_2202_nl;
  wire[0:0] mux_2201_nl;
  wire[0:0] and_592_nl;
  wire[0:0] mux_2200_nl;
  wire[0:0] nor_790_nl;
  wire[0:0] mux_2199_nl;
  wire[0:0] nand_436_nl;
  wire[0:0] nand_434_nl;
  wire[0:0] nor_791_nl;
  wire[0:0] mux_2198_nl;
  wire[0:0] nor_792_nl;
  wire[0:0] and_593_nl;
  wire[0:0] mux_2197_nl;
  wire[0:0] and_824_nl;
  wire[0:0] mux_2196_nl;
  wire[0:0] and_594_nl;
  wire[0:0] mux_2195_nl;
  wire[0:0] mux_2194_nl;
  wire[0:0] nor_794_nl;
  wire[0:0] mux_2193_nl;
  wire[0:0] mux_2192_nl;
  wire[0:0] nand_274_nl;
  wire[0:0] nand_275_nl;
  wire[0:0] mux_2191_nl;
  wire[0:0] or_2248_nl;
  wire[0:0] nand_277_nl;
  wire[0:0] mux_2190_nl;
  wire[0:0] mux_2189_nl;
  wire[0:0] nor_795_nl;
  wire[0:0] nor_796_nl;
  wire[0:0] mux_2188_nl;
  wire[0:0] or_2241_nl;
  wire[0:0] mux_2187_nl;
  wire[0:0] nor_797_nl;
  wire[0:0] and_596_nl;
  wire[0:0] mux_2186_nl;
  wire[0:0] nor_798_nl;
  wire[0:0] mux_2185_nl;
  wire[0:0] mux_2184_nl;
  wire[0:0] nand_409_nl;
  wire[0:0] mux_2183_nl;
  wire[0:0] or_2233_nl;
  wire[0:0] or_2230_nl;
  wire[0:0] mux_2182_nl;
  wire[0:0] and_597_nl;
  wire[0:0] mux_2181_nl;
  wire[0:0] and_598_nl;
  wire[0:0] mux_2180_nl;
  wire[0:0] and_599_nl;
  wire[0:0] nor_799_nl;
  wire[0:0] nor_800_nl;
  wire[0:0] nand_450_nl;
  wire[0:0] or_3357_nl;
  wire[0:0] mux_3723_nl;
  wire[0:0] mux_3722_nl;
  wire[0:0] mux_3721_nl;
  wire[0:0] nand_439_nl;
  wire[0:0] or_3373_nl;
  wire[0:0] mux_3720_nl;
  wire[0:0] or_3371_nl;
  wire[0:0] or_3369_nl;
  wire[0:0] or_3368_nl;
  wire[0:0] mux_3719_nl;
  wire[0:0] mux_3718_nl;
  wire[0:0] or_3367_nl;
  wire[0:0] or_3366_nl;
  wire[0:0] or_3365_nl;
  wire[0:0] mux_3717_nl;
  wire[0:0] nand_445_nl;
  wire[0:0] mux_3716_nl;
  wire[0:0] mux_3715_nl;
  wire[0:0] nor_1381_nl;
  wire[0:0] nor_1382_nl;
  wire[0:0] nor_1383_nl;
  wire[0:0] mux_3714_nl;
  wire[0:0] or_3358_nl;
  wire[0:0] mux_3713_nl;
  wire[0:0] mux_3712_nl;
  wire[0:0] or_3356_nl;
  wire[0:0] or_3355_nl;
  wire[0:0] nand_455_nl;
  wire[0:0] or_3396_nl;
  wire[0:0] or_3406_nl;
  wire[0:0] or_3409_nl;
  wire[0:0] mux_3771_nl;
  wire[0:0] or_3413_nl;
  wire[0:0] mux_3787_nl;
  wire[0:0] mux_3786_nl;
  wire[0:0] mux_3785_nl;
  wire[0:0] mux_3784_nl;
  wire[0:0] mux_3783_nl;
  wire[0:0] or_3420_nl;
  wire[0:0] mux_3782_nl;
  wire[0:0] or_3418_nl;
  wire[0:0] mux_3781_nl;
  wire[0:0] mux_3780_nl;
  wire[0:0] mux_3779_nl;
  wire[0:0] mux_3778_nl;
  wire[0:0] mux_3777_nl;
  wire[0:0] or_3417_nl;
  wire[0:0] mux_3776_nl;
  wire[0:0] or_3415_nl;
  wire[0:0] mux_3775_nl;
  wire[0:0] mux_3774_nl;
  wire[0:0] mux_3773_nl;
  wire[0:0] mux_3770_nl;
  wire[0:0] mux_3769_nl;
  wire[0:0] mux_3768_nl;
  wire[0:0] or_3411_nl;
  wire[0:0] mux_3767_nl;
  wire[0:0] mux_3766_nl;
  wire[0:0] mux_3765_nl;
  wire[0:0] mux_3764_nl;
  wire[0:0] mux_3762_nl;
  wire[0:0] mux_3761_nl;
  wire[0:0] mux_3760_nl;
  wire[0:0] or_3407_nl;
  wire[0:0] mux_3759_nl;
  wire[0:0] mux_3758_nl;
  wire[0:0] mux_3757_nl;
  wire[0:0] mux_3756_nl;
  wire[0:0] mux_3755_nl;
  wire[0:0] mux_3753_nl;
  wire[0:0] mux_3751_nl;
  wire[0:0] or_3403_nl;
  wire[0:0] mux_3750_nl;
  wire[0:0] mux_3749_nl;
  wire[0:0] mux_3748_nl;
  wire[0:0] or_3401_nl;
  wire[0:0] mux_3747_nl;
  wire[0:0] mux_3746_nl;
  wire[0:0] mux_3745_nl;
  wire[0:0] mux_3742_nl;
  wire[0:0] mux_3741_nl;
  wire[0:0] mux_3740_nl;
  wire[0:0] or_3395_nl;
  wire[0:0] mux_3739_nl;
  wire[0:0] or_3392_nl;
  wire[0:0] mux_3737_nl;
  wire[0:0] mux_3735_nl;
  wire[0:0] mux_3733_nl;
  wire[0:0] mux_3732_nl;
  wire[0:0] mux_3731_nl;
  wire[0:0] mux_3730_nl;
  wire[0:0] or_3384_nl;
  wire[0:0] mux_3728_nl;
  wire[0:0] mux_3727_nl;
  wire[0:0] or_3376_nl;
  wire[0:0] mux_3801_nl;
  wire[0:0] and_1248_nl;
  wire[0:0] mux_3800_nl;
  wire[0:0] nor_1369_nl;
  wire[0:0] and_1249_nl;
  wire[0:0] mux_3799_nl;
  wire[0:0] nor_1370_nl;
  wire[0:0] nor_1371_nl;
  wire[0:0] nor_1372_nl;
  wire[0:0] mux_3798_nl;
  wire[0:0] or_3441_nl;
  wire[0:0] mux_3797_nl;
  wire[0:0] or_3439_nl;
  wire[0:0] or_3438_nl;
  wire[0:0] mux_3796_nl;
  wire[0:0] mux_3795_nl;
  wire[0:0] mux_3794_nl;
  wire[0:0] mux_3793_nl;
  wire[0:0] nor_1373_nl;
  wire[0:0] nor_1374_nl;
  wire[0:0] nor_1375_nl;
  wire[0:0] nor_1376_nl;
  wire[0:0] mux_3792_nl;
  wire[0:0] or_3431_nl;
  wire[0:0] or_3430_nl;
  wire[0:0] mux_3791_nl;
  wire[0:0] and_1250_nl;
  wire[0:0] mux_3790_nl;
  wire[0:0] nor_1378_nl;
  wire[0:0] nor_1379_nl;
  wire[0:0] mux_3789_nl;
  wire[0:0] or_3424_nl;
  wire[0:0] or_3422_nl;
  wire[0:0] nor_1460_nl;
  wire[0:0] and_1267_nl;
  wire[0:0] mux_3898_nl;
  wire[0:0] or_3516_nl;
  wire[0:0] mux_3902_nl;
  wire[0:0] nand_470_nl;
  wire[0:0] or_3531_nl;
  wire[0:0] or_3530_nl;
  wire[0:0] mux_3906_nl;
  wire[10:0] acc_nl;
  wire[11:0] nl_acc_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_15_nl;
  wire[8:0] COMP_LOOP_COMP_LOOP_mux_18_nl;
  wire[0:0] COMP_LOOP_or_77_nl;
  wire[4:0] COMP_LOOP_COMP_LOOP_mux_19_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_16_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_17_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_18_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_19_nl;
  wire[9:0] COMP_LOOP_mux_84_nl;
  wire[4:0] COMP_LOOP_COMP_LOOP_mux_20_nl;
  wire[1:0] COMP_LOOP_COMP_LOOP_or_20_nl;
  wire[1:0] COMP_LOOP_mux_85_nl;
  wire[3:0] COMP_LOOP_mux1h_585_nl;
  wire[0:0] and_1278_nl;
  wire[0:0] and_1279_nl;
  wire[0:0] and_1280_nl;
  wire[1:0] COMP_LOOP_or_78_nl;
  wire[1:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_53_nl;
  wire[1:0] COMP_LOOP_mux_86_nl;
  wire[0:0] and_1281_nl;
  wire[0:0] and_1282_nl;
  wire[3:0] COMP_LOOP_mux1h_586_nl;
  wire[0:0] and_1283_nl;
  wire[0:0] and_1284_nl;
  wire[0:0] and_1285_nl;
  wire[63:0] COMP_LOOP_mux1h_587_nl;
  wire[63:0] COMP_LOOP_mux1h_588_nl;
  wire[63:0] operator_64_false_1_mux1h_2_nl;
  wire[63:0] operator_64_false_1_or_1_nl;
  wire[63:0] operator_64_false_1_mux1h_3_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_21_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_54_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_55_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_56_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_57_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_58_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_59_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_60_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_61_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_62_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_63_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_64_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_65_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_66_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_67_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_68_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_69_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_70_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_71_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_72_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_73_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_74_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_75_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_76_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_77_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_78_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_79_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_80_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_81_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_82_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_83_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_84_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_85_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_86_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_87_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_88_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_89_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_90_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_91_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_92_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_93_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_94_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_95_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_96_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_97_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_98_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_99_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_100_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_101_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_102_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_103_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_104_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_105_nl;
  wire[11:0] COMP_LOOP_mux1h_589_nl;
  wire[0:0] COMP_LOOP_or_79_nl;
  wire[6:0] COMP_LOOP_and_285_nl;
  wire[6:0] COMP_LOOP_mux1h_590_nl;
  wire[0:0] not_8636_nl;
  wire[2:0] COMP_LOOP_mux1h_591_nl;
  wire[0:0] COMP_LOOP_or_80_nl;
  wire[9:0] acc_8_nl;
  wire[10:0] nl_acc_8_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_22_nl;
  wire[0:0] COMP_LOOP_mux_87_nl;
  wire[0:0] COMP_LOOP_mux1h_592_nl;
  wire[0:0] COMP_LOOP_mux1h_593_nl;
  wire[0:0] COMP_LOOP_mux1h_594_nl;
  wire[0:0] COMP_LOOP_mux1h_595_nl;
  wire[0:0] COMP_LOOP_mux1h_596_nl;
  wire[0:0] COMP_LOOP_mux1h_597_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_mux_21_nl;
  wire[0:0] COMP_LOOP_or_81_nl;
  wire[0:0] COMP_LOOP_or_82_nl;
  wire[4:0] COMP_LOOP_COMP_LOOP_and_990_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_23_nl;
  wire[7:0] acc_9_nl;
  wire[8:0] nl_acc_9_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_24_nl;
  wire[5:0] COMP_LOOP_mux1h_598_nl;
  wire[0:0] COMP_LOOP_or_83_nl;
  wire[4:0] COMP_LOOP_COMP_LOOP_mux_22_nl;
  wire[0:0] COMP_LOOP_or_84_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_25_nl;
  wire[63:0] modExp_while_if_mux_1_nl;
  wire[0:0] mux_3954_nl;
  wire[0:0] mux_3955_nl;
  wire[0:0] mux_3956_nl;
  wire[0:0] mux_3957_nl;
  wire[0:0] mux_3958_nl;
  wire[0:0] nor_1463_nl;
  wire[0:0] nor_1464_nl;
  wire[0:0] nor_1465_nl;
  wire[0:0] mux_3959_nl;
  wire[0:0] nor_1466_nl;
  wire[0:0] mux_3960_nl;
  wire[0:0] nor_1467_nl;
  wire[0:0] nor_1468_nl;
  wire[0:0] mux_3961_nl;
  wire[0:0] mux_3962_nl;
  wire[0:0] nor_1469_nl;
  wire[0:0] nor_1470_nl;
  wire[0:0] mux_3963_nl;
  wire[0:0] nor_1471_nl;
  wire[0:0] nor_1472_nl;
  wire[0:0] mux_3964_nl;
  wire[0:0] or_3612_nl;
  wire[0:0] or_3613_nl;
  wire[0:0] mux_3965_nl;
  wire[0:0] mux_3966_nl;
  wire[0:0] and_1286_nl;
  wire[0:0] mux_3967_nl;
  wire[0:0] nor_1473_nl;
  wire[0:0] nor_1474_nl;
  wire[0:0] nor_1475_nl;
  wire[0:0] mux_3968_nl;
  wire[0:0] nor_1476_nl;
  wire[0:0] mux_3969_nl;
  wire[0:0] and_1287_nl;
  wire[0:0] nor_1477_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [10:0] nl_operator_66_true_div_cmp_b;
  assign nl_operator_66_true_div_cmp_b = {1'b0, operator_66_true_div_cmp_b_9_0};
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_8_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_8_tr0 = ~ (z_out_7[64]);
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_1_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_1_tr0 = ~ COMP_LOOP_nor_11_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_62_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_62_tr0 = ~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_2_modExp_1_while_C_38_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_2_modExp_1_while_C_38_tr0
      = ~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_124_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_124_tr0 = ~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_3_modExp_1_while_C_38_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_3_modExp_1_while_C_38_tr0
      = ~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_186_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_186_tr0 = ~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_4_modExp_1_while_C_38_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_4_modExp_1_while_C_38_tr0
      = ~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_248_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_248_tr0 = ~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_5_modExp_1_while_C_38_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_5_modExp_1_while_C_38_tr0
      = ~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_310_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_310_tr0 = ~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_6_modExp_1_while_C_38_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_6_modExp_1_while_C_38_tr0
      = ~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_372_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_372_tr0 = ~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_7_modExp_1_while_C_38_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_7_modExp_1_while_C_38_tr0
      = ~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_434_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_434_tr0 = ~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_8_modExp_1_while_C_38_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_8_modExp_1_while_C_38_tr0
      = ~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_496_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_496_tr0 = ~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_9_modExp_1_while_C_38_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_9_modExp_1_while_C_38_tr0
      = ~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_558_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_558_tr0 = ~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_10_modExp_1_while_C_38_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_10_modExp_1_while_C_38_tr0
      = ~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_620_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_620_tr0 = ~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_11_modExp_1_while_C_38_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_11_modExp_1_while_C_38_tr0
      = ~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_682_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_682_tr0 = ~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_12_modExp_1_while_C_38_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_12_modExp_1_while_C_38_tr0
      = ~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_744_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_744_tr0 = ~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_13_modExp_1_while_C_38_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_13_modExp_1_while_C_38_tr0
      = ~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_806_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_806_tr0 = ~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_14_modExp_1_while_C_38_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_14_modExp_1_while_C_38_tr0
      = ~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_868_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_868_tr0 = ~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_15_modExp_1_while_C_38_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_15_modExp_1_while_C_38_tr0
      = ~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_930_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_930_tr0 = ~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_16_modExp_1_while_C_38_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_16_modExp_1_while_C_38_tr0
      = ~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_C_0_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_C_0_tr0 = z_out_6[12];
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_9_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_9_tr0 = ~ STAGE_LOOP_acc_itm_2_1;
  ccs_in_v1 #(.rscid(32'sd2),
  .width(32'sd64)) p_rsci (
      .dat(p_rsc_dat),
      .idat(p_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd3),
  .width(32'sd64)) r_rsci (
      .dat(r_rsc_dat),
      .idat(r_rsci_idat)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_15_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_15_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_14_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_14_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_13_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_13_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_12_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_12_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_11_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_11_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_10_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_10_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_9_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_9_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_8_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_8_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_7_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_7_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_6_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_6_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_5_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_5_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_4_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_4_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_3_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_3_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_2_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_2_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_1_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_1_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_0_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_0_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) p_rsc_triosy_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(p_rsc_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) r_rsc_triosy_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(r_rsc_triosy_lz)
    );
  mgc_rem #(.width_a(32'sd64),
  .width_b(32'sd64),
  .signd(32'sd1)) modulo_result_rem_cmp (
      .a(modulo_result_rem_cmp_a),
      .b(modulo_result_rem_cmp_b),
      .z(modulo_result_rem_cmp_z)
    );
  mgc_div #(.width_a(32'sd65),
  .width_b(32'sd11),
  .signd(32'sd1)) operator_66_true_div_cmp (
      .a(operator_66_true_div_cmp_a),
      .b(nl_operator_66_true_div_cmp_b[10:0]),
      .z(operator_66_true_div_cmp_z)
    );
  mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd10)) STAGE_LOOP_lshift_rg (
      .a(1'b1),
      .s(STAGE_LOOP_i_3_0_sva),
      .z(STAGE_LOOP_lshift_psp_sva_mx0w0)
    );
  inPlaceNTT_DIT_core_core_fsm inPlaceNTT_DIT_core_core_fsm_inst (
      .clk(clk),
      .rst(rst),
      .fsm_output(fsm_output),
      .STAGE_LOOP_C_8_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_8_tr0[0:0]),
      .modExp_while_C_38_tr0(COMP_LOOP_COMP_LOOP_and_137_itm),
      .COMP_LOOP_C_1_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_1_tr0[0:0]),
      .COMP_LOOP_1_modExp_1_while_C_38_tr0(COMP_LOOP_COMP_LOOP_and_137_itm),
      .COMP_LOOP_C_62_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_62_tr0[0:0]),
      .COMP_LOOP_2_modExp_1_while_C_38_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_2_modExp_1_while_C_38_tr0[0:0]),
      .COMP_LOOP_C_124_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_124_tr0[0:0]),
      .COMP_LOOP_3_modExp_1_while_C_38_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_3_modExp_1_while_C_38_tr0[0:0]),
      .COMP_LOOP_C_186_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_186_tr0[0:0]),
      .COMP_LOOP_4_modExp_1_while_C_38_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_4_modExp_1_while_C_38_tr0[0:0]),
      .COMP_LOOP_C_248_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_248_tr0[0:0]),
      .COMP_LOOP_5_modExp_1_while_C_38_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_5_modExp_1_while_C_38_tr0[0:0]),
      .COMP_LOOP_C_310_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_310_tr0[0:0]),
      .COMP_LOOP_6_modExp_1_while_C_38_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_6_modExp_1_while_C_38_tr0[0:0]),
      .COMP_LOOP_C_372_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_372_tr0[0:0]),
      .COMP_LOOP_7_modExp_1_while_C_38_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_7_modExp_1_while_C_38_tr0[0:0]),
      .COMP_LOOP_C_434_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_434_tr0[0:0]),
      .COMP_LOOP_8_modExp_1_while_C_38_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_8_modExp_1_while_C_38_tr0[0:0]),
      .COMP_LOOP_C_496_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_496_tr0[0:0]),
      .COMP_LOOP_9_modExp_1_while_C_38_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_9_modExp_1_while_C_38_tr0[0:0]),
      .COMP_LOOP_C_558_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_558_tr0[0:0]),
      .COMP_LOOP_10_modExp_1_while_C_38_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_10_modExp_1_while_C_38_tr0[0:0]),
      .COMP_LOOP_C_620_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_620_tr0[0:0]),
      .COMP_LOOP_11_modExp_1_while_C_38_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_11_modExp_1_while_C_38_tr0[0:0]),
      .COMP_LOOP_C_682_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_682_tr0[0:0]),
      .COMP_LOOP_12_modExp_1_while_C_38_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_12_modExp_1_while_C_38_tr0[0:0]),
      .COMP_LOOP_C_744_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_744_tr0[0:0]),
      .COMP_LOOP_13_modExp_1_while_C_38_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_13_modExp_1_while_C_38_tr0[0:0]),
      .COMP_LOOP_C_806_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_806_tr0[0:0]),
      .COMP_LOOP_14_modExp_1_while_C_38_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_14_modExp_1_while_C_38_tr0[0:0]),
      .COMP_LOOP_C_868_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_868_tr0[0:0]),
      .COMP_LOOP_15_modExp_1_while_C_38_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_15_modExp_1_while_C_38_tr0[0:0]),
      .COMP_LOOP_C_930_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_930_tr0[0:0]),
      .COMP_LOOP_16_modExp_1_while_C_38_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_16_modExp_1_while_C_38_tr0[0:0]),
      .COMP_LOOP_C_992_tr0(COMP_LOOP_COMP_LOOP_and_10_itm),
      .VEC_LOOP_C_0_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_C_0_tr0[0:0]),
      .STAGE_LOOP_C_9_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_9_tr0[0:0])
    );
  assign nand_360_nl = ~((fsm_output[3]) & (fsm_output[6]) & (fsm_output[9]) & (fsm_output[8])
      & (~ (fsm_output[10])));
  assign or_619_nl = (fsm_output[3]) | (~ (fsm_output[6])) | (fsm_output[9]) | not_tmp_51;
  assign mux_1092_nl = MUX_s_1_2_2(nand_360_nl, or_619_nl, fsm_output[0]);
  assign or_621_cse = (fsm_output[5]) | mux_1092_nl;
  assign or_596_cse = (~ (fsm_output[5])) | (fsm_output[0]) | (fsm_output[3]) | (fsm_output[6])
      | (fsm_output[9]) | not_tmp_51;
  assign nor_223_cse = ~((fsm_output[7:6]!=2'b10));
  assign and_574_cse = (fsm_output[6]) & (fsm_output[0]) & (fsm_output[1]);
  assign or_2348_cse = (fsm_output[1:0]!=2'b00);
  assign and_573_cse = (fsm_output[1:0]==2'b11);
  assign and_563_cse = (fsm_output[2:1]==2'b11);
  assign or_2385_cse = (fsm_output[2:1]!=2'b00);
  assign and_565_cse = (fsm_output[2:0]==3'b111);
  assign nand_257_cse = ~((fsm_output[8]) & (fsm_output[6]));
  assign nand_375_cse = ~((fsm_output[7]) & (fsm_output[9]) & (fsm_output[10]));
  assign or_495_cse = (fsm_output[6:2]!=5'b00000);
  assign nand_376_cse = ~((fsm_output[10:9]==2'b11));
  assign nor_412_cse = ~((fsm_output[1:0]!=2'b10));
  assign and_528_cse = (fsm_output[6]) & (fsm_output[3]);
  assign nor_422_cse = ~((fsm_output[3]) | (~ (fsm_output[6])));
  assign and_472_cse = (fsm_output[9]) & (fsm_output[4]);
  assign or_2778_nl = (fsm_output[7]) | (~ (fsm_output[2])) | (~ (fsm_output[4]))
      | (fsm_output[10]);
  assign mux_3143_cse = MUX_s_1_2_2(or_tmp_2516, or_2778_nl, fsm_output[9]);
  assign nor_637_nl = ~((~ (fsm_output[9])) | (~ (fsm_output[7])) | (fsm_output[2])
      | (~ (fsm_output[4])) | (fsm_output[10]));
  assign nor_638_nl = ~((fsm_output[9]) | (fsm_output[7]) | (~ (fsm_output[2])) |
      (fsm_output[4]) | (~ (fsm_output[10])));
  assign mux_3145_nl = MUX_s_1_2_2(nor_637_nl, nor_638_nl, fsm_output[5]);
  assign and_466_nl = (fsm_output[1]) & mux_3145_nl;
  assign nor_639_nl = ~((fsm_output[1]) | (~ (fsm_output[5])) | (fsm_output[9]) |
      (~ (fsm_output[7])) | (fsm_output[2]) | nand_398_cse);
  assign mux_3146_nl = MUX_s_1_2_2(and_466_nl, nor_639_nl, fsm_output[6]);
  assign and_467_nl = (fsm_output[6]) & (fsm_output[1]) & (fsm_output[5]) & (~ (fsm_output[9]))
      & (fsm_output[7]) & (fsm_output[2]) & (fsm_output[4]) & (~ (fsm_output[10]));
  assign mux_3147_nl = MUX_s_1_2_2(mux_3146_nl, and_467_nl, fsm_output[3]);
  assign nor_640_nl = ~((~ (fsm_output[1])) | (~ (fsm_output[5])) | (fsm_output[9])
      | (~ (fsm_output[7])) | (fsm_output[2]) | nand_398_cse);
  assign nor_641_nl = ~((fsm_output[1]) | (fsm_output[5]) | mux_3143_cse);
  assign mux_3144_nl = MUX_s_1_2_2(nor_640_nl, nor_641_nl, fsm_output[6]);
  assign and_468_nl = (fsm_output[3]) & mux_3144_nl;
  assign mux_3148_nl = MUX_s_1_2_2(mux_3147_nl, and_468_nl, fsm_output[8]);
  assign nor_642_nl = ~((~ (fsm_output[1])) | (~ (fsm_output[5])) | (fsm_output[9])
      | (fsm_output[7]) | (fsm_output[2]) | (~ (fsm_output[4])) | (fsm_output[10]));
  assign and_469_nl = (fsm_output[1]) & (fsm_output[5]) & (fsm_output[9]) & (fsm_output[7])
      & (fsm_output[2]) & (fsm_output[4]) & (~ (fsm_output[10]));
  assign mux_3140_nl = MUX_s_1_2_2(nor_642_nl, and_469_nl, fsm_output[6]);
  assign or_2773_nl = (fsm_output[9]) | (~ (fsm_output[7])) | (fsm_output[2]) | (~
      (fsm_output[4])) | (fsm_output[10]);
  assign or_2772_nl = (~ (fsm_output[9])) | (fsm_output[7]) | (~ (fsm_output[2]))
      | (fsm_output[4]) | (fsm_output[10]);
  assign mux_3138_nl = MUX_s_1_2_2(or_2773_nl, or_2772_nl, fsm_output[5]);
  assign or_2770_nl = (~ (fsm_output[7])) | (fsm_output[2]) | (fsm_output[4]) | (~
      (fsm_output[10]));
  assign mux_3137_nl = MUX_s_1_2_2(or_2770_nl, or_tmp_2707, fsm_output[9]);
  assign or_2771_nl = (fsm_output[5]) | mux_3137_nl;
  assign mux_3139_nl = MUX_s_1_2_2(mux_3138_nl, or_2771_nl, fsm_output[1]);
  assign nor_643_nl = ~((fsm_output[6]) | mux_3139_nl);
  assign mux_3141_nl = MUX_s_1_2_2(mux_3140_nl, nor_643_nl, fsm_output[3]);
  assign mux_3135_nl = MUX_s_1_2_2(or_tmp_2707, or_tmp_2516, fsm_output[9]);
  assign nor_644_nl = ~((fsm_output[5]) | mux_3135_nl);
  assign nor_645_nl = ~((~ (fsm_output[5])) | (fsm_output[9]) | (fsm_output[7]) |
      (fsm_output[2]) | (fsm_output[4]) | (fsm_output[10]));
  assign mux_3136_nl = MUX_s_1_2_2(nor_644_nl, nor_645_nl, fsm_output[1]);
  assign and_470_nl = nor_422_cse & mux_3136_nl;
  assign mux_3142_nl = MUX_s_1_2_2(mux_3141_nl, and_470_nl, fsm_output[8]);
  assign mux_3149_nl = MUX_s_1_2_2(mux_3148_nl, mux_3142_nl, fsm_output[0]);
  assign and_353_nl = mux_3149_nl & COMP_LOOP_nor_11_itm;
  assign modExp_while_if_and_nl = modExp_while_and_3 & not_tmp_646;
  assign modExp_while_if_and_1_nl = modExp_while_and_5 & not_tmp_646;
  assign modExp_while_if_mux1h_nl = MUX1HOT_v_64_6_2(z_out_10, 64'b0000000000000000000000000000000000000000000000000000000000000001,
      COMP_LOOP_1_modExp_1_while_if_mul_mut_1, modulo_result_rem_cmp_z, (z_out_6[63:0]),
      z_out_5, {and_dcpl_260 , not_tmp_596 , and_353_nl , modExp_while_if_and_nl
      , modExp_while_if_and_1_nl , (~ mux_2475_itm)});
  assign and_284_nl = and_dcpl_118 & and_dcpl_98;
  assign mux_2560_nl = MUX_s_1_2_2(not_tmp_529, mux_tmp_2502, fsm_output[1]);
  assign mux_2559_nl = MUX_s_1_2_2(mux_tmp_2519, nor_tmp_342, and_573_cse);
  assign mux_2561_nl = MUX_s_1_2_2(mux_2560_nl, mux_2559_nl, fsm_output[9]);
  assign and_532_nl = (fsm_output[1]) & (fsm_output[2]) & (fsm_output[3]) & (fsm_output[10]);
  assign and_533_nl = (and_565_cse | (fsm_output[3])) & (fsm_output[10]);
  assign mux_2558_nl = MUX_s_1_2_2(and_532_nl, and_533_nl, fsm_output[9]);
  assign mux_2562_nl = MUX_s_1_2_2(mux_2561_nl, mux_2558_nl, fsm_output[6]);
  assign mux_2556_nl = MUX_s_1_2_2(and_dcpl_101, nor_tmp_6, or_3308_cse);
  assign or_2494_nl = (fsm_output[9]) | (~ mux_2556_nl);
  assign mux_2553_nl = MUX_s_1_2_2(mux_tmp_2519, nor_tmp_342, fsm_output[1]);
  assign and_535_nl = (and_563_cse | (fsm_output[3])) & (fsm_output[10]);
  assign mux_2554_nl = MUX_s_1_2_2(mux_2553_nl, and_535_nl, fsm_output[0]);
  assign or_2491_nl = nor_784_cse | (~ (fsm_output[2])) | (~ (fsm_output[3])) | (fsm_output[10]);
  assign mux_2555_nl = MUX_s_1_2_2((~ mux_2554_nl), or_2491_nl, fsm_output[9]);
  assign mux_2557_nl = MUX_s_1_2_2(or_2494_nl, mux_2555_nl, fsm_output[6]);
  assign mux_2563_nl = MUX_s_1_2_2(mux_2562_nl, mux_2557_nl, fsm_output[7]);
  assign mux_2551_nl = MUX_s_1_2_2(and_816_cse, mux_tmp_2549, fsm_output[6]);
  assign nor_731_nl = ~(and_563_cse | (fsm_output[3]) | (fsm_output[10]));
  assign mux_2548_nl = MUX_s_1_2_2(nor_731_nl, (fsm_output[10]), fsm_output[9]);
  assign mux_2550_nl = MUX_s_1_2_2(mux_tmp_2549, mux_2548_nl, fsm_output[6]);
  assign mux_2552_nl = MUX_s_1_2_2(mux_2551_nl, mux_2550_nl, fsm_output[7]);
  assign mux_2564_nl = MUX_s_1_2_2(mux_2563_nl, mux_2552_nl, fsm_output[8]);
  assign mux_2544_nl = MUX_s_1_2_2(nor_tmp_342, or_tmp_2429, fsm_output[9]);
  assign mux_2542_nl = MUX_s_1_2_2(nor_tmp_338, or_tmp_2416, fsm_output[0]);
  assign mux_2543_nl = MUX_s_1_2_2((~ mux_2542_nl), mux_tmp_2502, fsm_output[9]);
  assign mux_2545_nl = MUX_s_1_2_2((~ mux_2544_nl), mux_2543_nl, fsm_output[6]);
  assign mux_2540_nl = MUX_s_1_2_2(and_dcpl_101, nor_tmp_6, and_563_cse);
  assign or_2484_nl = (fsm_output[9]) | (~ mux_2540_nl);
  assign mux_2541_nl = MUX_s_1_2_2(and_816_cse, or_2484_nl, fsm_output[6]);
  assign mux_2546_nl = MUX_s_1_2_2(mux_2545_nl, mux_2541_nl, fsm_output[7]);
  assign mux_2536_nl = MUX_s_1_2_2(mux_tmp_2502, mux_tmp_2523, fsm_output[1]);
  assign mux_2537_nl = MUX_s_1_2_2(mux_2536_nl, mux_tmp_2525, fsm_output[0]);
  assign or_2483_nl = (fsm_output[9]) | (~ mux_2537_nl);
  assign nor_732_nl = ~((fsm_output[0]) | (fsm_output[1]) | (fsm_output[2]) | (fsm_output[3])
      | (fsm_output[10]));
  assign mux_2535_nl = MUX_s_1_2_2(nor_732_nl, (fsm_output[10]), fsm_output[9]);
  assign mux_2538_nl = MUX_s_1_2_2(or_2483_nl, mux_2535_nl, fsm_output[6]);
  assign or_2480_nl = (or_3308_cse & (fsm_output[3])) | (fsm_output[10]);
  assign mux_2534_nl = MUX_s_1_2_2(nor_tmp_338, or_2480_nl, fsm_output[9]);
  assign mux_2539_nl = MUX_s_1_2_2(mux_2538_nl, mux_2534_nl, fsm_output[7]);
  assign mux_2547_nl = MUX_s_1_2_2(mux_2546_nl, mux_2539_nl, fsm_output[8]);
  assign mux_2565_nl = MUX_s_1_2_2(mux_2564_nl, mux_2547_nl, fsm_output[5]);
  assign mux_2528_nl = MUX_s_1_2_2(and_dcpl_101, nor_tmp_6, and_540_cse);
  assign mux_2529_nl = MUX_s_1_2_2(not_tmp_529, mux_2528_nl, fsm_output[9]);
  assign mux_2524_nl = MUX_s_1_2_2(mux_tmp_2523, mux_tmp_2519, fsm_output[1]);
  assign mux_2526_nl = MUX_s_1_2_2(mux_tmp_2525, mux_2524_nl, fsm_output[0]);
  assign mux_2527_nl = MUX_s_1_2_2(not_tmp_529, mux_2526_nl, fsm_output[9]);
  assign mux_2530_nl = MUX_s_1_2_2(mux_2529_nl, mux_2527_nl, fsm_output[6]);
  assign nor_733_nl = ~(and_565_cse | (fsm_output[3]) | (fsm_output[10]));
  assign mux_2521_nl = MUX_s_1_2_2(nor_733_nl, (fsm_output[10]), fsm_output[9]);
  assign mux_2520_nl = MUX_s_1_2_2(mux_tmp_2519, or_tmp_2419, fsm_output[9]);
  assign mux_2522_nl = MUX_s_1_2_2(mux_2521_nl, mux_2520_nl, fsm_output[6]);
  assign mux_2531_nl = MUX_s_1_2_2((~ mux_2530_nl), mux_2522_nl, fsm_output[7]);
  assign mux_2516_nl = MUX_s_1_2_2(nor_tmp_6, or_tmp_2419, fsm_output[9]);
  assign or_2475_nl = (~((fsm_output[2:1]!=2'b00))) | (~ (fsm_output[3])) | (fsm_output[10]);
  assign mux_2515_nl = MUX_s_1_2_2((~ nor_tmp_330), or_2475_nl, fsm_output[9]);
  assign mux_2517_nl = MUX_s_1_2_2(mux_2516_nl, mux_2515_nl, fsm_output[6]);
  assign or_2472_nl = (~(and_565_cse | (fsm_output[3]))) | (fsm_output[10]);
  assign mux_2513_nl = MUX_s_1_2_2((~ or_tmp_2416), or_2472_nl, fsm_output[9]);
  assign mux_2514_nl = MUX_s_1_2_2(mux_2513_nl, and_816_cse, fsm_output[6]);
  assign mux_2518_nl = MUX_s_1_2_2(mux_2517_nl, mux_2514_nl, fsm_output[7]);
  assign mux_2532_nl = MUX_s_1_2_2(mux_2531_nl, mux_2518_nl, fsm_output[8]);
  assign mux_2510_nl = MUX_s_1_2_2(nor_1203_cse, mux_tmp_2508, fsm_output[6]);
  assign or_2466_nl = (~(and_540_cse | (fsm_output[3]))) | (fsm_output[10]);
  assign mux_2507_nl = MUX_s_1_2_2(not_tmp_529, or_2466_nl, fsm_output[9]);
  assign mux_2509_nl = MUX_s_1_2_2(mux_tmp_2508, mux_2507_nl, fsm_output[6]);
  assign mux_2511_nl = MUX_s_1_2_2(mux_2510_nl, mux_2509_nl, fsm_output[7]);
  assign mux_2503_nl = MUX_s_1_2_2(not_tmp_529, mux_tmp_2502, or_2348_cse);
  assign or_2460_nl = nor_738_cse | (fsm_output[10]);
  assign mux_2504_nl = MUX_s_1_2_2(mux_2503_nl, or_2460_nl, fsm_output[9]);
  assign and_544_nl = or_2348_cse & (fsm_output[2]) & (fsm_output[3]) & (fsm_output[10]);
  assign mux_2500_nl = MUX_s_1_2_2(and_544_nl, (fsm_output[10]), fsm_output[9]);
  assign mux_2505_nl = MUX_s_1_2_2(mux_2504_nl, mux_2500_nl, fsm_output[6]);
  assign nand_247_nl = ~((fsm_output[0]) & (fsm_output[1]) & (fsm_output[2]) & (fsm_output[3])
      & (~ (fsm_output[10])));
  assign mux_2498_nl = MUX_s_1_2_2((~ nor_tmp_6), nand_247_nl, fsm_output[9]);
  assign nand_248_nl = ~((and_540_cse | (fsm_output[3])) & (fsm_output[10]));
  assign or_2454_nl = (~ (fsm_output[2])) | (~ (fsm_output[3])) | (fsm_output[10]);
  assign mux_2497_nl = MUX_s_1_2_2(nand_248_nl, or_2454_nl, fsm_output[9]);
  assign mux_2499_nl = MUX_s_1_2_2(mux_2498_nl, mux_2497_nl, fsm_output[6]);
  assign mux_2506_nl = MUX_s_1_2_2(mux_2505_nl, mux_2499_nl, fsm_output[7]);
  assign mux_2512_nl = MUX_s_1_2_2(mux_2511_nl, mux_2506_nl, fsm_output[8]);
  assign mux_2533_nl = MUX_s_1_2_2(mux_2532_nl, mux_2512_nl, fsm_output[5]);
  assign mux_2566_nl = MUX_s_1_2_2(mux_2565_nl, mux_2533_nl, fsm_output[4]);
  assign operator_64_false_mux1h_2_rgt = MUX1HOT_v_65_3_2(z_out_6, ({2'b00 , operator_64_false_slc_modExp_exp_63_1_3}),
      ({1'b0 , modExp_while_if_mux1h_nl}), {and_284_nl , and_dcpl_273 , (~ mux_2566_nl)});
  assign and_1262_cse = (fsm_output[3]) & (fsm_output[9]);
  assign nor_1450_cse = ~((~ (fsm_output[1])) | COMP_LOOP_nor_11_itm);
  assign or_3328_cse = (fsm_output[9:8]!=2'b00);
  assign or_2520_cse = (fsm_output[7:6]!=2'b00);
  assign and_754_cse = or_3328_cse & (fsm_output[10]);
  assign and_300_m1c = and_dcpl_191 & and_dcpl_279;
  assign and_816_cse = (fsm_output[10:9]==2'b11);
  assign and_815_cse = (fsm_output[7]) & (fsm_output[9]) & (fsm_output[10]);
  assign modExp_result_and_rgt = (~ modExp_while_and_5) & and_300_m1c;
  assign modExp_result_and_1_rgt = modExp_while_and_5 & and_300_m1c;
  assign or_15_cse = (~((fsm_output[6]) | (~ (fsm_output[3])))) | (fsm_output[10]);
  assign nand_402_cse = ~((fsm_output[3]) & (fsm_output[0]) & (fsm_output[1]) & (~
      (fsm_output[10])));
  assign mux_28_cse = MUX_s_1_2_2((~ (fsm_output[10])), or_tmp_21, fsm_output[6]);
  assign or_36_cse = (fsm_output[6]) | (~ nor_tmp_6);
  assign mux_3_cse = MUX_s_1_2_2(or_tmp_4, or_tmp_3, fsm_output[7]);
  assign mux_7_cse = MUX_s_1_2_2(or_tmp_9, (fsm_output[10]), fsm_output[6]);
  assign mux_9_cse = MUX_s_1_2_2((fsm_output[10]), nand_402_cse, fsm_output[6]);
  assign nand_240_cse = ~((fsm_output[7]) & (fsm_output[4]) & (fsm_output[10]));
  assign or_2591_nl = (~ (fsm_output[5])) | (~ (fsm_output[1])) | (fsm_output[9])
      | (fsm_output[2]) | nand_240_cse;
  assign or_2588_nl = (~ (fsm_output[9])) | (~ (fsm_output[2])) | (fsm_output[7])
      | (fsm_output[4]) | (~ (fsm_output[10]));
  assign mux_2767_nl = MUX_s_1_2_2(mux_3143_cse, or_2588_nl, fsm_output[1]);
  assign or_2589_nl = (fsm_output[5]) | mux_2767_nl;
  assign mux_2768_nl = MUX_s_1_2_2(or_2591_nl, or_2589_nl, fsm_output[6]);
  assign nor_694_nl = ~((fsm_output[3]) | mux_2768_nl);
  assign nor_695_nl = ~((fsm_output[5]) | (~ (fsm_output[1])) | mux_3143_cse);
  assign nor_696_nl = ~((~ (fsm_output[5])) | (fsm_output[1]) | mux_tmp_2758);
  assign mux_2766_nl = MUX_s_1_2_2(nor_695_nl, nor_696_nl, fsm_output[6]);
  assign and_513_nl = (fsm_output[3]) & mux_2766_nl;
  assign mux_2769_nl = MUX_s_1_2_2(nor_694_nl, and_513_nl, fsm_output[8]);
  assign nor_697_nl = ~((~ (fsm_output[5])) | (fsm_output[1]) | (~ (fsm_output[9]))
      | (fsm_output[2]) | (~ (fsm_output[7])) | (~ (fsm_output[4])) | (fsm_output[10]));
  assign or_2581_nl = (fsm_output[9]) | (~ (fsm_output[2])) | (fsm_output[7]) | (fsm_output[4])
      | (~ (fsm_output[10]));
  assign or_2579_nl = (fsm_output[9]) | (fsm_output[2]) | (fsm_output[7]) | (~ (fsm_output[4]))
      | (fsm_output[10]);
  assign mux_2762_nl = MUX_s_1_2_2(or_2581_nl, or_2579_nl, fsm_output[1]);
  assign nor_698_nl = ~((fsm_output[5]) | mux_2762_nl);
  assign mux_2763_nl = MUX_s_1_2_2(nor_697_nl, nor_698_nl, fsm_output[6]);
  assign and_514_nl = (fsm_output[3]) & mux_2763_nl;
  assign and_515_nl = (fsm_output[1]) & (~ mux_tmp_2758);
  assign nor_699_nl = ~((fsm_output[1]) | (fsm_output[9]) | (~ (fsm_output[2])) |
      (fsm_output[7]) | (fsm_output[4]) | (fsm_output[10]));
  assign mux_2759_nl = MUX_s_1_2_2(and_515_nl, nor_699_nl, fsm_output[5]);
  assign nor_700_nl = ~((~ (fsm_output[5])) | (fsm_output[1]) | (fsm_output[9]) |
      (fsm_output[2]) | (~ (fsm_output[7])) | (fsm_output[4]) | (~ (fsm_output[10])));
  assign mux_2760_nl = MUX_s_1_2_2(mux_2759_nl, nor_700_nl, fsm_output[6]);
  assign nor_701_nl = ~((~ (fsm_output[6])) | (~ (fsm_output[5])) | (~ (fsm_output[1]))
      | (fsm_output[9]) | (~ (fsm_output[2])) | (~ (fsm_output[7])) | (fsm_output[4])
      | (fsm_output[10]));
  assign mux_2761_nl = MUX_s_1_2_2(mux_2760_nl, nor_701_nl, fsm_output[3]);
  assign mux_2764_nl = MUX_s_1_2_2(and_514_nl, mux_2761_nl, fsm_output[8]);
  assign mux_2770_m1c = MUX_s_1_2_2(mux_2769_nl, mux_2764_nl, fsm_output[0]);
  assign and_517_cse = (fsm_output[6]) & (fsm_output[0]) & (fsm_output[3]);
  assign nand_398_cse = ~((fsm_output[4]) & (fsm_output[10]));
  assign nand_237_cse = ~((fsm_output[1:0]==2'b11));
  assign modulo_result_mux_1_cse = MUX_v_64_2_2(modulo_result_rem_cmp_z, (z_out_6[63:0]),
      modulo_result_rem_cmp_z[63]);
  assign nor_1302_nl = ~((fsm_output[7]) | (~ (fsm_output[9])) | (fsm_output[8])
      | (fsm_output[4]) | (fsm_output[10]));
  assign and_801_nl = (fsm_output[7]) & (fsm_output[9]) & (fsm_output[8]) & (fsm_output[4])
      & (~ (fsm_output[10]));
  assign mux_71_cse = MUX_s_1_2_2(nor_1302_nl, and_801_nl, fsm_output[2]);
  assign nor_715_nl = ~((fsm_output[6]) | (fsm_output[0]) | (fsm_output[3]));
  assign mux_2742_nl = MUX_s_1_2_2(and_517_cse, nor_715_nl, fsm_output[5]);
  assign and_345_m1c = mux_2742_nl & and_dcpl_26 & (~ (fsm_output[7])) & (~ (fsm_output[2]))
      & (~ (fsm_output[8])) & and_dcpl_30;
  assign or_2679_cse = (fsm_output[8]) | (~ (fsm_output[9])) | (fsm_output[5]) |
      (fsm_output[10]);
  assign nor_381_cse = ~((fsm_output[4]) | (~ (fsm_output[2])) | (~ (fsm_output[6])));
  assign nor_670_cse = ~((~ (fsm_output[8])) | (fsm_output[9]) | (fsm_output[5])
      | (fsm_output[10]));
  assign or_212_cse = (fsm_output[8]) | (fsm_output[4]);
  assign and_491_cse = (fsm_output[4]) & (fsm_output[10]);
  assign or_2729_cse = (fsm_output[8]) | and_491_cse;
  assign or_199_nl = (fsm_output[8]) | (~ or_tmp_182);
  assign mux_384_cse = MUX_s_1_2_2(or_199_nl, nand_tmp_12, fsm_output[6]);
  assign mux_382_cse = MUX_s_1_2_2(mux_tmp_381, mux_tmp_379, fsm_output[1]);
  assign COMP_LOOP_or_32_cse = and_dcpl_126 | and_dcpl_141 | and_dcpl_147 | and_dcpl_158
      | and_dcpl_164 | and_dcpl_175 | and_dcpl_182 | and_dcpl_192 | and_dcpl_198
      | and_dcpl_206 | and_dcpl_217 | and_dcpl_225 | and_dcpl_232 | and_dcpl_242
      | and_dcpl_247 | and_dcpl_255;
  assign or_2824_cse = (fsm_output[3]) | (~ (fsm_output[1])) | (~ (fsm_output[9]))
      | (~ (fsm_output[4])) | (fsm_output[10]);
  assign nand_226_cse = ~((fsm_output[3]) & (fsm_output[1]) & (fsm_output[9]) & (fsm_output[4])
      & (fsm_output[10]));
  assign or_2826_cse = (fsm_output[3]) | (fsm_output[1]) | (fsm_output[9]) | (fsm_output[4])
      | (~ (fsm_output[10]));
  assign or_2839_cse = (~ (fsm_output[0])) | (~ (fsm_output[3])) | (~ (fsm_output[1]))
      | (fsm_output[9]) | (fsm_output[4]) | (fsm_output[10]);
  assign and_464_cse = (fsm_output[0]) & (fsm_output[3]) & (fsm_output[1]) & (fsm_output[9])
      & (fsm_output[4]) & (~ (fsm_output[10]));
  assign or_2819_cse = (fsm_output[0]) | (fsm_output[3]) | (fsm_output[1]) | (fsm_output[9])
      | nand_398_cse;
  assign or_2894_cse = (fsm_output[3:1]!=3'b000);
  assign and_458_cse = (fsm_output[3:1]==3'b111);
  assign and_459_cse = (fsm_output[3:2]==2'b11);
  assign and_359_cse = (fsm_output[5:4]==2'b11) & or_2894_cse;
  assign and_456_cse = (fsm_output[5:4]==2'b11);
  assign or_2898_cse = (fsm_output[3]) | (fsm_output[6]);
  assign and_450_cse = (fsm_output[7:6]==2'b11);
  assign or_2902_cse = and_573_cse | (fsm_output[3]);
  assign nor_1316_cse = ~((fsm_output[8:6]!=3'b000));
  assign nor_610_cse = ~((fsm_output[9:8]!=2'b00));
  assign and_440_cse = (fsm_output[3:0]==4'b1111);
  assign or_2935_cse = (fsm_output[8:7]!=2'b00);
  assign mux_726_cse = MUX_s_1_2_2((~ (fsm_output[10])), (fsm_output[10]), fsm_output[9]);
  assign or_3308_cse = (fsm_output[2:0]!=3'b000);
  assign or_2951_cse = (fsm_output[8:6]!=3'b000);
  assign nor_1203_cse = ~((fsm_output[2]) | (fsm_output[1]) | (fsm_output[3]) | (fsm_output[9])
      | (fsm_output[10]));
  assign nor_601_cse = ~((fsm_output[10:9]!=2'b00));
  assign or_3002_cse = (fsm_output[2]) | (fsm_output[7]) | (fsm_output[8]) | (~ (fsm_output[4]))
      | (fsm_output[10]);
  assign or_3018_cse = (~ (fsm_output[5])) | (fsm_output[1]) | (fsm_output[2]) |
      (~ (fsm_output[7])) | (fsm_output[8]) | nand_398_cse;
  assign or_3016_cse = (fsm_output[1]) | (~ (fsm_output[2])) | (fsm_output[7]) |
      not_tmp_34;
  assign or_3014_nl = (~ (fsm_output[1])) | (fsm_output[2]) | (fsm_output[7]) | (~
      (fsm_output[8])) | (fsm_output[4]) | (fsm_output[10]);
  assign mux_3393_nl = MUX_s_1_2_2(or_3016_cse, or_3014_nl, fsm_output[5]);
  assign mux_3394_cse = MUX_s_1_2_2(or_3018_cse, mux_3393_nl, fsm_output[0]);
  assign or_3004_nl = (~ (fsm_output[2])) | (fsm_output[7]) | (fsm_output[8]) | (fsm_output[4])
      | (~ (fsm_output[10]));
  assign mux_3384_nl = MUX_s_1_2_2(or_3004_nl, or_3002_cse, fsm_output[1]);
  assign or_3001_nl = (~ (fsm_output[1])) | (~ (fsm_output[2])) | (~ (fsm_output[7]))
      | (~ (fsm_output[8])) | (fsm_output[4]) | (fsm_output[10]);
  assign mux_3385_cse = MUX_s_1_2_2(mux_3384_nl, or_3001_nl, fsm_output[5]);
  assign nor_581_nl = ~((fsm_output[0]) | mux_tmp_3386);
  assign nor_582_nl = ~((~ (fsm_output[5])) | (~ (fsm_output[1])) | (fsm_output[2])
      | (fsm_output[7]) | not_tmp_34);
  assign nor_583_nl = ~((fsm_output[7]) | (fsm_output[8]) | (fsm_output[4]) | (~
      (fsm_output[10])));
  assign and_415_nl = (fsm_output[7]) & (fsm_output[8]) & (fsm_output[4]) & (fsm_output[10]);
  assign mux_3389_nl = MUX_s_1_2_2(nor_583_nl, and_415_nl, fsm_output[2]);
  assign and_414_nl = (fsm_output[1]) & mux_3389_nl;
  assign nor_584_nl = ~((fsm_output[1]) | (~ (fsm_output[2])) | (~ (fsm_output[7]))
      | (~ (fsm_output[8])) | (fsm_output[4]) | (fsm_output[10]));
  assign mux_3390_nl = MUX_s_1_2_2(and_414_nl, nor_584_nl, fsm_output[5]);
  assign mux_3391_nl = MUX_s_1_2_2(nor_582_nl, mux_3390_nl, fsm_output[0]);
  assign mux_3392_cse = MUX_s_1_2_2(nor_581_nl, mux_3391_nl, fsm_output[6]);
  assign and_416_nl = (fsm_output[0]) & (~ mux_tmp_3386);
  assign nor_585_nl = ~((fsm_output[0]) | mux_3385_cse);
  assign mux_3387_nl = MUX_s_1_2_2(and_416_nl, nor_585_nl, fsm_output[6]);
  assign nor_586_nl = ~((fsm_output[6]) | (fsm_output[0]) | (fsm_output[5]) | (fsm_output[1])
      | (~ (fsm_output[2])) | (fsm_output[7]) | (~ (fsm_output[8])) | (~ (fsm_output[4]))
      | (fsm_output[10]));
  assign mux_3388_cse = MUX_s_1_2_2(mux_3387_nl, nor_586_nl, fsm_output[3]);
  assign or_3241_nl = (fsm_output[7]) | (fsm_output[8]) | (fsm_output[4]) | (~ (fsm_output[10]));
  assign nand_205_nl = ~((fsm_output[7]) & (fsm_output[8]) & (fsm_output[4]) & (fsm_output[10]));
  assign mux_3498_cse = MUX_s_1_2_2(or_3241_nl, nand_205_nl, fsm_output[2]);
  assign mux_3556_nl = MUX_s_1_2_2(nand_tmp_157, nand_tmp_12, fsm_output[1]);
  assign mux_3557_cse = MUX_s_1_2_2(or_tmp_191, mux_3556_nl, fsm_output[6]);
  assign mux_3056_nl = MUX_s_1_2_2(and_491_cse, (fsm_output[4]), fsm_output[9]);
  assign or_3120_nl = (fsm_output[8]) | mux_3056_nl;
  assign mux_3572_nl = MUX_s_1_2_2(or_2729_cse, or_3120_nl, fsm_output[1]);
  assign mux_3573_nl = MUX_s_1_2_2(nand_tmp_157, mux_3572_nl, fsm_output[6]);
  assign mux_433_nl = MUX_s_1_2_2((~ mux_tmp_380), or_tmp_182, fsm_output[8]);
  assign or_3119_nl = (fsm_output[8]) | (~ mux_tmp_380);
  assign mux_3569_nl = MUX_s_1_2_2(mux_433_nl, or_3119_nl, and_573_cse);
  assign mux_3567_nl = MUX_s_1_2_2(nand_tmp_14, nand_tmp_157, fsm_output[1]);
  assign mux_3570_nl = MUX_s_1_2_2(mux_3569_nl, mux_3567_nl, fsm_output[6]);
  assign mux_3574_nl = MUX_s_1_2_2(mux_3573_nl, mux_3570_nl, fsm_output[5]);
  assign mux_437_nl = MUX_s_1_2_2(mux_tmp_399, mux_tmp_375, or_2348_cse);
  assign mux_438_nl = MUX_s_1_2_2(mux_437_nl, nand_tmp_14, fsm_output[6]);
  assign mux_431_nl = MUX_s_1_2_2(or_tmp_189, mux_tmp_399, fsm_output[6]);
  assign mux_3566_nl = MUX_s_1_2_2(mux_438_nl, mux_431_nl, fsm_output[5]);
  assign mux_3575_cse = MUX_s_1_2_2(mux_3574_nl, mux_3566_nl, fsm_output[7]);
  assign mux_3554_nl = MUX_s_1_2_2(mux_tmp_373, nand_tmp_157, fsm_output[6]);
  assign mux_419_nl = MUX_s_1_2_2(or_tmp_188, mux_tmp_381, or_2348_cse);
  assign mux_420_nl = MUX_s_1_2_2(mux_419_nl, mux_tmp_375, fsm_output[6]);
  assign mux_3555_cse = MUX_s_1_2_2(mux_3554_nl, mux_420_nl, fsm_output[5]);
  assign nand_201_cse = ~((fsm_output[9]) & (fsm_output[4]) & (fsm_output[10]));
  assign mux_3547_nl = MUX_s_1_2_2(nand_tmp_157, nand_tmp_12, or_2348_cse);
  assign mux_3548_nl = MUX_s_1_2_2(mux_3547_nl, mux_tmp_381, fsm_output[6]);
  assign or_3115_nl = (fsm_output[8]) | (~ mux_tmp_378);
  assign mux_403_nl = MUX_s_1_2_2(or_3115_nl, or_tmp_191, or_2348_cse);
  assign mux_3546_nl = MUX_s_1_2_2(mux_403_nl, nand_tmp_157, fsm_output[6]);
  assign mux_3549_nl = MUX_s_1_2_2(mux_3548_nl, mux_3546_nl, fsm_output[5]);
  assign mux_3542_nl = MUX_s_1_2_2(nand_tmp_14, nand_tmp_157, and_573_cse);
  assign mux_3543_nl = MUX_s_1_2_2(mux_tmp_375, mux_3542_nl, fsm_output[6]);
  assign mux_401_nl = MUX_s_1_2_2(or_tmp_189, or_tmp_188, and_573_cse);
  assign mux_400_nl = MUX_s_1_2_2(mux_tmp_399, mux_tmp_375, fsm_output[1]);
  assign mux_402_nl = MUX_s_1_2_2(mux_401_nl, mux_400_nl, fsm_output[6]);
  assign mux_3544_nl = MUX_s_1_2_2(mux_3543_nl, mux_402_nl, fsm_output[5]);
  assign mux_3550_nl = MUX_s_1_2_2(mux_3549_nl, mux_3544_nl, fsm_output[7]);
  assign nand_173_nl = ~((fsm_output[8]) & (~ mux_tmp_380));
  assign mux_3532_nl = MUX_s_1_2_2(nand_201_cse, mux_tmp_380, fsm_output[8]);
  assign mux_3533_nl = MUX_s_1_2_2(nand_173_nl, mux_3532_nl, fsm_output[1]);
  assign mux_3534_nl = MUX_s_1_2_2(mux_3533_nl, mux_tmp_3323, fsm_output[6]);
  assign mux_3535_nl = MUX_s_1_2_2(mux_3534_nl, mux_384_cse, fsm_output[5]);
  assign mux_3527_nl = MUX_s_1_2_2(nand_tmp_157, nand_tmp_12, and_573_cse);
  assign mux_3528_nl = MUX_s_1_2_2(or_tmp_180, mux_3527_nl, fsm_output[6]);
  assign mux_376_nl = MUX_s_1_2_2(mux_tmp_375, or_tmp_181, fsm_output[1]);
  assign mux_377_nl = MUX_s_1_2_2(mux_376_nl, mux_tmp_373, fsm_output[0]);
  assign mux_383_nl = MUX_s_1_2_2(mux_382_cse, mux_377_nl, fsm_output[6]);
  assign mux_3529_nl = MUX_s_1_2_2(mux_3528_nl, mux_383_nl, fsm_output[5]);
  assign mux_3536_nl = MUX_s_1_2_2(mux_3535_nl, mux_3529_nl, fsm_output[7]);
  assign mux_3551_cse = MUX_s_1_2_2(mux_3550_nl, mux_3536_nl, fsm_output[3]);
  assign nor_544_cse = ~((~ (fsm_output[3])) | (~ (fsm_output[7])) | (~ (fsm_output[2]))
      | (fsm_output[9]) | (fsm_output[8]) | (fsm_output[4]) | (~ (fsm_output[10])));
  assign nor_539_cse = ~((fsm_output[7]) | (~ (fsm_output[2])) | (fsm_output[9])
      | (fsm_output[8]) | (fsm_output[4]) | (~ (fsm_output[10])));
  assign nor_515_cse = ~((fsm_output[5]) | (~ (fsm_output[3])));
  assign nor_540_nl = ~((~ (fsm_output[7])) | (fsm_output[2]) | (fsm_output[9]) |
      not_tmp_34);
  assign mux_3603_cse = MUX_s_1_2_2(nor_539_cse, nor_540_nl, fsm_output[3]);
  assign nor_545_cse = ~((fsm_output[5]) | (fsm_output[3]) | (fsm_output[7]) | (fsm_output[2])
      | (fsm_output[9]) | not_tmp_34);
  assign nl_STAGE_LOOP_i_3_0_sva_2 = STAGE_LOOP_i_3_0_sva + 4'b0001;
  assign STAGE_LOOP_i_3_0_sva_2 = nl_STAGE_LOOP_i_3_0_sva_2[3:0];
  assign nl_COMP_LOOP_acc_psp_sva_1 = (VEC_LOOP_j_sva_11_0[11:4]) + conv_u2u_5_8(COMP_LOOP_k_9_4_sva_4_0);
  assign COMP_LOOP_acc_psp_sva_1 = nl_COMP_LOOP_acc_psp_sva_1[7:0];
  assign or_529_cse = (fsm_output[1]) | (~ (fsm_output[9])) | (~ (fsm_output[3]))
      | (fsm_output[4]) | (fsm_output[10]);
  assign or_525_cse = (~ (fsm_output[1])) | (~ (fsm_output[9])) | (~ (fsm_output[3]))
      | (fsm_output[4]) | (fsm_output[10]);
  assign nl_COMP_LOOP_1_modExp_1_while_if_mul_mut_1 = $signed(operator_64_false_acc_mut_63_0)
      * $signed(COMP_LOOP_10_mul_mut);
  assign COMP_LOOP_1_modExp_1_while_if_mul_mut_1 = nl_COMP_LOOP_1_modExp_1_while_if_mul_mut_1[63:0];
  assign operator_64_false_slc_modExp_exp_63_1_3 = MUX_v_63_2_2((operator_66_true_div_cmp_z[63:1]),
      (tmp_10_lpi_4_dfm[63:1]), and_dcpl_281);
  assign nor_1276_cse = ~((fsm_output[2]) | (~ (fsm_output[7])) | (fsm_output[3])
      | (fsm_output[8]) | (~ (fsm_output[4])) | (~ (fsm_output[9])) | (fsm_output[10]));
  assign nor_1279_cse = ~((~ (fsm_output[5])) | (~ (fsm_output[2])) | (~ (fsm_output[7]))
      | (~ (fsm_output[3])) | (fsm_output[8]) | (~ (fsm_output[4])) | (fsm_output[9])
      | (fsm_output[10]));
  assign nl_COMP_LOOP_acc_1_cse_6_sva_1 = VEC_LOOP_j_sva_11_0 + conv_u2u_9_12({COMP_LOOP_k_9_4_sva_4_0
      , 4'b0101});
  assign COMP_LOOP_acc_1_cse_6_sva_1 = nl_COMP_LOOP_acc_1_cse_6_sva_1[11:0];
  assign nl_COMP_LOOP_acc_1_cse_2_sva_1 = VEC_LOOP_j_sva_11_0 + conv_u2u_9_12({COMP_LOOP_k_9_4_sva_4_0
      , 4'b0001});
  assign COMP_LOOP_acc_1_cse_2_sva_1 = nl_COMP_LOOP_acc_1_cse_2_sva_1[11:0];
  assign or_163_cse = (fsm_output[4]) | (~ (fsm_output[8])) | (fsm_output[10]);
  assign nl_COMP_LOOP_k_9_4_sva_2 = conv_u2u_5_6(COMP_LOOP_k_9_4_sva_4_0) + 6'b000001;
  assign COMP_LOOP_k_9_4_sva_2 = nl_COMP_LOOP_k_9_4_sva_2[5:0];
  assign modExp_while_and_3 = (~ (modulo_result_rem_cmp_z[63])) & COMP_LOOP_nor_11_itm;
  assign modExp_while_and_5 = (modulo_result_rem_cmp_z[63]) & COMP_LOOP_nor_11_itm;
  assign or_tmp_3 = (~ (fsm_output[6])) | (fsm_output[3]) | (fsm_output[10]);
  assign or_tmp_4 = (~ (fsm_output[6])) | (fsm_output[10]);
  assign or_tmp_8 = nor_422_cse | (fsm_output[10]);
  assign or_tmp_9 = (fsm_output[3]) | (fsm_output[1]) | (fsm_output[10]);
  assign or_tmp_14 = (fsm_output[6]) | (fsm_output[10]);
  assign nor_tmp_6 = (fsm_output[3]) & (fsm_output[10]);
  assign or_tmp_21 = (fsm_output[3]) | (fsm_output[10]);
  assign nor_tmp_9 = ((fsm_output[0]) | (fsm_output[1]) | (fsm_output[3])) & (fsm_output[10]);
  assign not_tmp_34 = ~((fsm_output[8]) & (fsm_output[4]) & (fsm_output[10]));
  assign not_tmp_45 = ~((fsm_output[5]) & (fsm_output[10]));
  assign or_tmp_110 = (fsm_output[8]) | (fsm_output[10]);
  assign not_tmp_51 = ~((fsm_output[8]) & (fsm_output[10]));
  assign or_tmp_118 = (~ (fsm_output[8])) | (fsm_output[10]);
  assign or_tmp_141 = (fsm_output[4]) | (fsm_output[8]) | (fsm_output[10]);
  assign or_154_cse = (~ (fsm_output[4])) | (fsm_output[8]) | (fsm_output[10]);
  assign mux_tmp_207 = MUX_s_1_2_2(or_154_cse, or_tmp_141, fsm_output[5]);
  assign mux_tmp_226 = MUX_s_1_2_2(or_tmp_141, or_tmp_118, fsm_output[5]);
  assign or_tmp_150 = (~ (fsm_output[4])) | (fsm_output[8]);
  assign or_tmp_178 = (~ (fsm_output[4])) | (fsm_output[10]);
  assign or_tmp_179 = (fsm_output[4]) | (fsm_output[10]);
  assign mux_371_nl = MUX_s_1_2_2((~ or_tmp_179), or_tmp_178, fsm_output[9]);
  assign or_tmp_180 = (fsm_output[8]) | mux_371_nl;
  assign mux_372_nl = MUX_s_1_2_2((~ (fsm_output[4])), or_tmp_178, fsm_output[9]);
  assign or_tmp_181 = (fsm_output[8]) | mux_372_nl;
  assign mux_tmp_373 = MUX_s_1_2_2(or_tmp_181, or_tmp_180, fsm_output[1]);
  assign or_tmp_182 = (fsm_output[9]) | (fsm_output[4]) | (fsm_output[10]);
  assign mux_tmp_374 = MUX_s_1_2_2((~ and_491_cse), or_tmp_178, fsm_output[9]);
  assign mux_tmp_375 = MUX_s_1_2_2(mux_tmp_374, or_tmp_182, fsm_output[8]);
  assign or_tmp_183 = (fsm_output[9]) | (~ and_491_cse);
  assign mux_tmp_378 = MUX_s_1_2_2((fsm_output[4]), or_tmp_179, fsm_output[9]);
  assign mux_tmp_379 = MUX_s_1_2_2(mux_tmp_378, or_tmp_183, fsm_output[8]);
  assign mux_tmp_380 = MUX_s_1_2_2(and_491_cse, or_tmp_179, fsm_output[9]);
  assign mux_tmp_381 = MUX_s_1_2_2(mux_tmp_380, or_tmp_183, fsm_output[8]);
  assign or_2747_cse = (fsm_output[9]) | (fsm_output[4]);
  assign nor_tmp_46 = or_2747_cse & (fsm_output[10]);
  assign nand_tmp_12 = ~((fsm_output[8]) & (~ nor_tmp_46));
  assign nand_tmp_13 = ~((fsm_output[8]) & (~ and_816_cse));
  assign or_tmp_187 = (fsm_output[10:9]!=2'b00);
  assign mux_tmp_399 = MUX_s_1_2_2(or_tmp_183, or_tmp_179, fsm_output[8]);
  assign or_tmp_188 = (fsm_output[8]) | mux_tmp_380;
  assign or_tmp_189 = (fsm_output[8]) | nor_tmp_46;
  assign or_tmp_191 = (fsm_output[8]) | (~ or_tmp_179);
  assign mux_406_nl = MUX_s_1_2_2(or_tmp_179, (~ (fsm_output[10])), fsm_output[9]);
  assign nand_tmp_14 = ~((fsm_output[8]) & mux_406_nl);
  assign or_tmp_195 = (fsm_output[9]) | (~ (fsm_output[4])) | (fsm_output[10]);
  assign mux_tmp_412 = MUX_s_1_2_2(or_tmp_195, nor_tmp_46, fsm_output[8]);
  assign mux_tmp_413 = MUX_s_1_2_2(or_tmp_195, and_816_cse, fsm_output[8]);
  assign and_dcpl = ~((fsm_output[4]) | (fsm_output[9]));
  assign and_dcpl_1 = (fsm_output[5]) & (fsm_output[2]);
  assign and_dcpl_2 = and_dcpl_1 & (~ (fsm_output[8]));
  assign or_tmp_237 = (~ (fsm_output[3])) | (fsm_output[10]);
  assign nor_tmp_116 = (fsm_output[9:8]==2'b11);
  assign mux_tmp_741 = MUX_s_1_2_2((~ (fsm_output[10])), (fsm_output[10]), or_3328_cse);
  assign or_tmp_434 = (fsm_output[6]) | (~ (fsm_output[10]));
  assign mux_tmp_893 = MUX_s_1_2_2((~ (fsm_output[10])), (fsm_output[10]), fsm_output[6]);
  assign mux_tmp_917 = MUX_s_1_2_2(or_tmp_434, or_tmp_4, fsm_output[8]);
  assign and_dcpl_21 = (~ (fsm_output[5])) & (fsm_output[2]);
  assign and_dcpl_22 = and_dcpl_21 & (fsm_output[8]);
  assign and_dcpl_26 = ~((fsm_output[10]) | (fsm_output[1]));
  assign and_dcpl_30 = (fsm_output[4]) & (~ (fsm_output[9]));
  assign and_dcpl_31 = (fsm_output[5]) & (~ (fsm_output[2]));
  assign and_dcpl_32 = and_dcpl_31 & (fsm_output[8]);
  assign and_dcpl_40 = and_dcpl_21 & (~ (fsm_output[8]));
  assign and_dcpl_46 = and_dcpl_31 & (~ (fsm_output[8]));
  assign and_dcpl_50 = (~ (fsm_output[4])) & (fsm_output[9]);
  assign or_3295_nl = (fsm_output[0]) | (fsm_output[1]) | (fsm_output[7]) | (fsm_output[9])
      | (fsm_output[10]);
  assign mux_1027_nl = MUX_s_1_2_2(or_3295_nl, nand_375_cse, or_495_cse);
  assign not_tmp_219 = MUX_s_1_2_2(mux_1027_nl, nand_376_cse, fsm_output[8]);
  assign and_dcpl_96 = ~((fsm_output[5]) | (fsm_output[2]));
  assign and_dcpl_97 = and_dcpl_96 & (~ (fsm_output[8]));
  assign and_dcpl_98 = and_dcpl_97 & and_dcpl;
  assign and_dcpl_99 = ~((fsm_output[0]) | (fsm_output[6]));
  assign and_dcpl_100 = and_dcpl_99 & (~ (fsm_output[7]));
  assign and_dcpl_101 = ~((fsm_output[10]) | (fsm_output[3]));
  assign and_dcpl_102 = and_dcpl_101 & (~ (fsm_output[1]));
  assign and_dcpl_103 = and_dcpl_102 & and_dcpl_100;
  assign and_dcpl_106 = and_dcpl_97 & and_dcpl_50;
  assign and_dcpl_107 = (fsm_output[0]) & (~ (fsm_output[6]));
  assign and_dcpl_108 = and_dcpl_107 & (fsm_output[7]);
  assign and_dcpl_109 = (fsm_output[10]) & (~ (fsm_output[3]));
  assign and_dcpl_110 = and_dcpl_109 & (fsm_output[1]);
  assign and_dcpl_111 = and_dcpl_110 & and_dcpl_108;
  assign and_dcpl_116 = and_dcpl_46 & and_dcpl_30;
  assign and_dcpl_117 = and_dcpl_107 & (~ (fsm_output[7]));
  assign and_dcpl_118 = and_dcpl_102 & and_dcpl_117;
  assign and_dcpl_119 = and_dcpl_118 & and_dcpl_116;
  assign and_dcpl_121 = (~ (fsm_output[0])) & (fsm_output[6]);
  assign and_dcpl_122 = and_dcpl_121 & (~ (fsm_output[7]));
  assign and_dcpl_123 = (~ (fsm_output[10])) & (fsm_output[3]);
  assign and_dcpl_124 = and_dcpl_123 & (fsm_output[1]);
  assign and_dcpl_125 = and_dcpl_124 & and_dcpl_122;
  assign and_dcpl_126 = and_dcpl_125 & and_dcpl_97 & and_dcpl_30;
  assign and_dcpl_127 = and_dcpl_99 & (fsm_output[7]);
  assign and_dcpl_128 = and_dcpl_101 & (fsm_output[1]);
  assign and_dcpl_129 = and_dcpl_128 & and_dcpl_127;
  assign or_tmp_453 = (fsm_output[1]) | (~ (fsm_output[9])) | (~ (fsm_output[3]))
      | (~ (fsm_output[4])) | (fsm_output[10]);
  assign and_659_nl = (fsm_output[5]) & (fsm_output[6]) & (fsm_output[0]);
  assign nor_1193_nl = ~((fsm_output[5]) | (fsm_output[6]) | (fsm_output[0]));
  assign not_tmp_240 = MUX_s_1_2_2(and_659_nl, nor_1193_nl, fsm_output[4]);
  assign and_dcpl_139 = and_dcpl_2 & and_dcpl_30;
  assign and_dcpl_140 = and_dcpl_124 & and_dcpl_108;
  assign and_dcpl_141 = and_dcpl_140 & and_dcpl_139;
  assign and_dcpl_145 = and_dcpl_1 & (fsm_output[8]);
  assign and_dcpl_146 = and_dcpl_145 & and_dcpl;
  assign and_dcpl_147 = and_dcpl_103 & and_dcpl_146;
  assign and_dcpl_148 = (fsm_output[9:8]==2'b01);
  assign and_dcpl_154 = and_dcpl_96 & (fsm_output[8]);
  assign and_dcpl_156 = and_dcpl_123 & (~ (fsm_output[1]));
  assign and_dcpl_158 = and_dcpl_156 & and_dcpl_108 & and_dcpl_154 & and_dcpl;
  assign and_dcpl_162 = and_dcpl_121 & (fsm_output[7]);
  assign and_dcpl_164 = and_dcpl_124 & and_dcpl_162 & and_dcpl_146;
  assign and_dcpl_165 = (fsm_output[9:8]==2'b10);
  assign nor_tmp_217 = (fsm_output[6]) & (fsm_output[0]);
  assign mux_tmp_1049 = MUX_s_1_2_2(and_dcpl_99, nor_tmp_217, fsm_output[4]);
  assign and_dcpl_172 = and_dcpl_97 & and_472_cse;
  assign and_dcpl_173 = nor_tmp_217 & (~ (fsm_output[7]));
  assign and_dcpl_175 = and_dcpl_128 & and_dcpl_173 & and_dcpl_172;
  assign and_dcpl_182 = and_dcpl_156 & and_dcpl_127 & and_dcpl_46 & and_472_cse;
  assign and_dcpl_191 = and_dcpl_156 & and_dcpl_117;
  assign and_dcpl_192 = and_dcpl_191 & and_dcpl_22 & and_472_cse;
  assign and_dcpl_198 = and_dcpl_129 & and_dcpl_154 & and_dcpl_50;
  assign and_dcpl_204 = nor_tmp_217 & (fsm_output[7]);
  assign and_dcpl_206 = and_dcpl_128 & and_dcpl_204 & and_dcpl_145 & and_dcpl_50;
  assign and_dcpl_215 = nor_tmp_6 & (~ (fsm_output[1]));
  assign and_dcpl_217 = and_dcpl_215 & and_dcpl_122 & and_dcpl_40 & and_dcpl;
  assign and_dcpl_223 = and_dcpl_109 & (~ (fsm_output[1]));
  assign and_dcpl_225 = and_dcpl_223 & and_dcpl_108 & and_dcpl_116;
  assign and_dcpl_232 = and_dcpl_110 & and_dcpl_100 & and_dcpl_22 & and_dcpl_30;
  assign and_dcpl_239 = and_dcpl_32 & and_dcpl_30;
  assign and_dcpl_240 = nor_tmp_6 & (fsm_output[1]);
  assign and_dcpl_242 = and_dcpl_240 & and_dcpl_173 & and_dcpl_239;
  assign and_dcpl_243 = (fsm_output[10]) & (~ (fsm_output[6]));
  assign and_dcpl_245 = and_dcpl_32 & and_dcpl;
  assign and_dcpl_247 = and_dcpl_223 & and_dcpl_162 & and_dcpl_245;
  assign and_dcpl_255 = and_dcpl_223 & and_dcpl_173 & and_dcpl_40 & and_dcpl_50;
  assign or_tmp_515 = (COMP_LOOP_acc_19_psp_sva[1:0]!=2'b00) | (fsm_output[0]) |
      (VEC_LOOP_j_sva_11_0[1:0]!=2'b00) | (~ (fsm_output[3])) | (fsm_output[6]) |
      (fsm_output[9]) | not_tmp_51;
  assign or_tmp_518 = (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b0000) | (fsm_output[5])
      | (~ (fsm_output[0])) | (~ (fsm_output[3])) | (fsm_output[6]) | (fsm_output[9])
      | (fsm_output[8]) | (~ (fsm_output[10]));
  assign or_579_nl = (VEC_LOOP_j_sva_11_0[3]) | (fsm_output[0]) | (VEC_LOOP_j_sva_11_0[2:0]!=3'b000)
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[9]) | (fsm_output[8]) | (fsm_output[10]);
  assign or_578_nl = (COMP_LOOP_acc_16_psp_sva[0]) | (VEC_LOOP_j_sva_11_0[2:0]!=3'b000)
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[9])) | (~ (fsm_output[8]))
      | (fsm_output[10]);
  assign or_577_nl = (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b0000) | (fsm_output[3])
      | (fsm_output[6]) | (fsm_output[9]) | not_tmp_51;
  assign mux_1061_nl = MUX_s_1_2_2(or_578_nl, or_577_nl, fsm_output[0]);
  assign mux_tmp_1062 = MUX_s_1_2_2(or_579_nl, mux_1061_nl, fsm_output[5]);
  assign or_587_nl = (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b000) | (VEC_LOOP_j_sva_11_0[0])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[9]) | (~ (fsm_output[8]))
      | (fsm_output[10]);
  assign or_586_nl = (COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b0000) | (fsm_output[3])
      | (~ (fsm_output[6])) | (~ (fsm_output[9])) | (~ (fsm_output[8])) | (fsm_output[10]);
  assign mux_1065_nl = MUX_s_1_2_2(or_587_nl, or_586_nl, fsm_output[0]);
  assign or_585_nl = (COMP_LOOP_acc_1_cse_sva[3:0]!=4'b0000) | (~ (fsm_output[0]))
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (~ (fsm_output[9])) | (fsm_output[8])
      | (~ (fsm_output[10]));
  assign mux_1066_nl = MUX_s_1_2_2(mux_1065_nl, or_585_nl, fsm_output[5]);
  assign or_583_nl = (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b000) | (~ (fsm_output[5]))
      | (fsm_output[0]) | (VEC_LOOP_j_sva_11_0[0]) | (fsm_output[3]) | (~ (fsm_output[6]))
      | (fsm_output[9]) | (fsm_output[8]) | (~ (fsm_output[10]));
  assign mux_tmp_1067 = MUX_s_1_2_2(mux_1066_nl, or_583_nl, fsm_output[4]);
  assign or_591_nl = (COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b0000) | (~ (fsm_output[0]))
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[9]) | (fsm_output[8])
      | (~ (fsm_output[10]));
  assign or_589_nl = (~ (fsm_output[0])) | (fsm_output[3]) | (fsm_output[6]) | (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b0000)
      | (fsm_output[10:8]!=3'b001);
  assign mux_tmp_1068 = MUX_s_1_2_2(or_591_nl, or_589_nl, fsm_output[5]);
  assign or_622_cse = (~ (fsm_output[0])) | (~ (fsm_output[3])) | (fsm_output[6])
      | (~ (fsm_output[9])) | (fsm_output[8]) | (fsm_output[10]);
  assign or_617_cse = (fsm_output[0]) | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[9]))
      | (fsm_output[8]) | (~ (fsm_output[10]));
  assign or_614_nl = (fsm_output[0]) | (fsm_output[3]) | (~ (fsm_output[6])) | (fsm_output[9])
      | (~ (fsm_output[8])) | (fsm_output[10]);
  assign or_613_nl = (fsm_output[0]) | (~ (fsm_output[3])) | (~ (fsm_output[6]))
      | (fsm_output[9]) | (fsm_output[8]) | (~ (fsm_output[10]));
  assign mux_1087_nl = MUX_s_1_2_2(or_614_nl, or_613_nl, fsm_output[5]);
  assign or_611_nl = (~ (fsm_output[0])) | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[9])
      | (fsm_output[8]) | (fsm_output[10]);
  assign or_610_nl = (~ (fsm_output[0])) | (~ (fsm_output[3])) | (fsm_output[6])
      | (~ (fsm_output[9])) | (~ (fsm_output[8])) | (fsm_output[10]);
  assign mux_1086_nl = MUX_s_1_2_2(or_611_nl, or_610_nl, fsm_output[5]);
  assign mux_1088_cse = MUX_s_1_2_2(mux_1087_nl, mux_1086_nl, fsm_output[4]);
  assign or_609_cse = (~ (fsm_output[5])) | (fsm_output[0]) | (fsm_output[3]) | (fsm_output[6])
      | (fsm_output[9]) | (fsm_output[8]) | (~ (fsm_output[10]));
  assign or_607_cse = (~ (fsm_output[0])) | (~ (fsm_output[3])) | (fsm_output[6])
      | (~ (fsm_output[9])) | (fsm_output[8]) | (~ (fsm_output[10]));
  assign nor_1170_nl = ~((~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[9])
      | (fsm_output[8]) | (fsm_output[10]));
  assign nor_1171_nl = ~((fsm_output[3]) | (~ (fsm_output[6])) | (~ (fsm_output[9]))
      | (fsm_output[8]) | (fsm_output[10]));
  assign mux_1080_nl = MUX_s_1_2_2(nor_1170_nl, nor_1171_nl, fsm_output[0]);
  assign nand_25_cse = ~((fsm_output[5]) & mux_1080_nl);
  assign or_601_cse = (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[9])
      | (~ (fsm_output[8])) | (fsm_output[10]);
  assign or_600_nl = (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[9]))
      | (fsm_output[8]) | (fsm_output[10]);
  assign or_599_nl = (fsm_output[3]) | (fsm_output[6]) | (fsm_output[9]) | (fsm_output[8])
      | (~ (fsm_output[10]));
  assign mux_1073_cse = MUX_s_1_2_2(or_600_nl, or_599_nl, fsm_output[0]);
  assign not_tmp_260 = ~((fsm_output[1]) & (fsm_output[10]));
  assign or_tmp_626 = (COMP_LOOP_acc_19_psp_sva[1:0]!=2'b00) | (fsm_output[0]) |
      (VEC_LOOP_j_sva_11_0[1:0]!=2'b01) | (~ (fsm_output[3])) | (fsm_output[6]) |
      (fsm_output[9]) | not_tmp_51;
  assign or_tmp_630 = (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b0001) | (fsm_output[5])
      | (~ (fsm_output[0])) | (~ (fsm_output[3])) | (fsm_output[6]) | (fsm_output[9])
      | (fsm_output[8]) | (~ (fsm_output[10]));
  assign or_693_nl = (VEC_LOOP_j_sva_11_0[3]) | (fsm_output[0]) | (VEC_LOOP_j_sva_11_0[2:0]!=3'b001)
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[9]) | (fsm_output[8]) | (fsm_output[10]);
  assign or_692_nl = (COMP_LOOP_acc_16_psp_sva[0]) | (VEC_LOOP_j_sva_11_0[2:0]!=3'b001)
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[9])) | (~ (fsm_output[8]))
      | (fsm_output[10]);
  assign or_691_nl = (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b0001) | (fsm_output[3])
      | (fsm_output[6]) | (fsm_output[9]) | not_tmp_51;
  assign mux_1138_nl = MUX_s_1_2_2(or_692_nl, or_691_nl, fsm_output[0]);
  assign mux_tmp_1139 = MUX_s_1_2_2(or_693_nl, mux_1138_nl, fsm_output[5]);
  assign or_709_nl = (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b000) | (~ (VEC_LOOP_j_sva_11_0[0]))
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[9]) | (~ (fsm_output[8]))
      | (fsm_output[10]);
  assign or_708_nl = (COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b0001) | (fsm_output[3])
      | (~ (fsm_output[6])) | (~ (fsm_output[9])) | (~ (fsm_output[8])) | (fsm_output[10]);
  assign mux_1148_nl = MUX_s_1_2_2(or_709_nl, or_708_nl, fsm_output[0]);
  assign or_707_nl = (COMP_LOOP_acc_1_cse_sva[3:0]!=4'b0001) | (~ (fsm_output[0]))
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (~ (fsm_output[9])) | (fsm_output[8])
      | (~ (fsm_output[10]));
  assign mux_1149_nl = MUX_s_1_2_2(mux_1148_nl, or_707_nl, fsm_output[5]);
  assign or_705_nl = (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b000) | (~ (fsm_output[5]))
      | (fsm_output[0]) | (~ (VEC_LOOP_j_sva_11_0[0])) | (fsm_output[3]) | (~ (fsm_output[6]))
      | (fsm_output[9]) | (fsm_output[8]) | (~ (fsm_output[10]));
  assign mux_tmp_1150 = MUX_s_1_2_2(mux_1149_nl, or_705_nl, fsm_output[4]);
  assign or_712_nl = (COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b0001) | (~ (fsm_output[0]))
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[9]) | (fsm_output[8])
      | (~ (fsm_output[10]));
  assign or_710_nl = (~ (fsm_output[0])) | (fsm_output[3]) | (fsm_output[6]) | (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b0001)
      | (fsm_output[10:8]!=3'b001);
  assign mux_tmp_1152 = MUX_s_1_2_2(or_712_nl, or_710_nl, fsm_output[5]);
  assign or_tmp_728 = (COMP_LOOP_acc_19_psp_sva[1:0]!=2'b00) | (fsm_output[0]) |
      (VEC_LOOP_j_sva_11_0[1:0]!=2'b10) | (~ (fsm_output[3])) | (fsm_output[6]) |
      (fsm_output[9]) | not_tmp_51;
  assign or_tmp_731 = (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b0010) | (fsm_output[5])
      | (~ (fsm_output[0])) | (~ (fsm_output[3])) | (fsm_output[6]) | (fsm_output[9])
      | (fsm_output[8]) | (~ (fsm_output[10]));
  assign or_792_nl = (VEC_LOOP_j_sva_11_0[3]) | (fsm_output[0]) | (VEC_LOOP_j_sva_11_0[2:0]!=3'b010)
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[9]) | (fsm_output[8]) | (fsm_output[10]);
  assign or_791_nl = (COMP_LOOP_acc_16_psp_sva[0]) | (VEC_LOOP_j_sva_11_0[2:0]!=3'b010)
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[9])) | (~ (fsm_output[8]))
      | (fsm_output[10]);
  assign or_790_nl = (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b0010) | (fsm_output[3])
      | (fsm_output[6]) | (fsm_output[9]) | not_tmp_51;
  assign mux_1205_nl = MUX_s_1_2_2(or_791_nl, or_790_nl, fsm_output[0]);
  assign mux_tmp_1206 = MUX_s_1_2_2(or_792_nl, mux_1205_nl, fsm_output[5]);
  assign or_800_nl = (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b001) | (VEC_LOOP_j_sva_11_0[0])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[9]) | (~ (fsm_output[8]))
      | (fsm_output[10]);
  assign or_799_nl = (COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b0010) | (fsm_output[3])
      | (~ (fsm_output[6])) | (~ (fsm_output[9])) | (~ (fsm_output[8])) | (fsm_output[10]);
  assign mux_1209_nl = MUX_s_1_2_2(or_800_nl, or_799_nl, fsm_output[0]);
  assign or_798_nl = (COMP_LOOP_acc_1_cse_sva[3:0]!=4'b0010) | (~ (fsm_output[0]))
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (~ (fsm_output[9])) | (fsm_output[8])
      | (~ (fsm_output[10]));
  assign mux_1210_nl = MUX_s_1_2_2(mux_1209_nl, or_798_nl, fsm_output[5]);
  assign or_796_nl = (~ (fsm_output[5])) | (fsm_output[0]) | (VEC_LOOP_j_sva_11_0[0])
      | (fsm_output[3]) | (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b001) | (~ (fsm_output[6]))
      | (fsm_output[9]) | (fsm_output[8]) | (~ (fsm_output[10]));
  assign mux_tmp_1211 = MUX_s_1_2_2(mux_1210_nl, or_796_nl, fsm_output[4]);
  assign or_804_nl = (COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b0010) | (~ (fsm_output[0]))
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[9]) | (fsm_output[8])
      | (~ (fsm_output[10]));
  assign or_802_nl = (~ (fsm_output[0])) | (fsm_output[3]) | (fsm_output[6]) | (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b0010)
      | (fsm_output[10:8]!=3'b001);
  assign mux_tmp_1212 = MUX_s_1_2_2(or_804_nl, or_802_nl, fsm_output[5]);
  assign or_tmp_839 = (COMP_LOOP_acc_19_psp_sva[1:0]!=2'b00) | (fsm_output[0]) |
      (VEC_LOOP_j_sva_11_0[1:0]!=2'b11) | (~ (fsm_output[3])) | (fsm_output[6]) |
      (fsm_output[9]) | not_tmp_51;
  assign or_tmp_843 = (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b0011) | (fsm_output[5])
      | (~ (fsm_output[0])) | (~ (fsm_output[3])) | (fsm_output[6]) | (fsm_output[9])
      | (fsm_output[8]) | (~ (fsm_output[10]));
  assign or_906_nl = (VEC_LOOP_j_sva_11_0[3]) | (fsm_output[0]) | (VEC_LOOP_j_sva_11_0[2:0]!=3'b011)
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[9]) | (fsm_output[8]) | (fsm_output[10]);
  assign or_905_nl = (COMP_LOOP_acc_16_psp_sva[0]) | (VEC_LOOP_j_sva_11_0[2:0]!=3'b011)
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[9])) | (~ (fsm_output[8]))
      | (fsm_output[10]);
  assign or_904_nl = (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b0011) | (fsm_output[3])
      | (fsm_output[6]) | (fsm_output[9]) | not_tmp_51;
  assign mux_1282_nl = MUX_s_1_2_2(or_905_nl, or_904_nl, fsm_output[0]);
  assign mux_tmp_1283 = MUX_s_1_2_2(or_906_nl, mux_1282_nl, fsm_output[5]);
  assign or_922_nl = (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b001) | (~ (VEC_LOOP_j_sva_11_0[0]))
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[9]) | (~ (fsm_output[8]))
      | (fsm_output[10]);
  assign or_921_nl = (COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b0011) | (fsm_output[3])
      | (~ (fsm_output[6])) | (~ (fsm_output[9])) | (~ (fsm_output[8])) | (fsm_output[10]);
  assign mux_1292_nl = MUX_s_1_2_2(or_922_nl, or_921_nl, fsm_output[0]);
  assign nand_433_nl = ~((COMP_LOOP_acc_1_cse_sva[3:0]==4'b0011) & (fsm_output[0])
      & (fsm_output[3]) & (fsm_output[6]) & (fsm_output[9]) & (~ (fsm_output[8]))
      & (fsm_output[10]));
  assign mux_1293_nl = MUX_s_1_2_2(mux_1292_nl, nand_433_nl, fsm_output[5]);
  assign or_918_nl = (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b001) | (~ (fsm_output[5]))
      | (fsm_output[0]) | (~ (VEC_LOOP_j_sva_11_0[0])) | (fsm_output[3]) | (~ (fsm_output[6]))
      | (fsm_output[9]) | (fsm_output[8]) | (~ (fsm_output[10]));
  assign mux_tmp_1294 = MUX_s_1_2_2(mux_1293_nl, or_918_nl, fsm_output[4]);
  assign or_925_nl = (COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b0011) | (~ (fsm_output[0]))
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[9]) | (fsm_output[8])
      | (~ (fsm_output[10]));
  assign or_923_nl = (~ (fsm_output[0])) | (fsm_output[3]) | (fsm_output[6]) | (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b0011)
      | (fsm_output[10:8]!=3'b001);
  assign mux_tmp_1296 = MUX_s_1_2_2(or_925_nl, or_923_nl, fsm_output[5]);
  assign or_tmp_941 = (COMP_LOOP_acc_19_psp_sva[1:0]!=2'b01) | (fsm_output[0]) |
      (VEC_LOOP_j_sva_11_0[1:0]!=2'b00) | (~ (fsm_output[3])) | (fsm_output[6]) |
      (fsm_output[9]) | not_tmp_51;
  assign or_tmp_944 = (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b0100) | (fsm_output[5])
      | (~ (fsm_output[0])) | (~ (fsm_output[3])) | (fsm_output[6]) | (fsm_output[9])
      | (fsm_output[8]) | (~ (fsm_output[10]));
  assign or_1005_nl = (VEC_LOOP_j_sva_11_0[3]) | (fsm_output[0]) | (VEC_LOOP_j_sva_11_0[2:0]!=3'b100)
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[9]) | (fsm_output[8]) | (fsm_output[10]);
  assign or_1004_nl = (COMP_LOOP_acc_16_psp_sva[0]) | (VEC_LOOP_j_sva_11_0[2:0]!=3'b100)
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[9])) | (~ (fsm_output[8]))
      | (fsm_output[10]);
  assign or_1003_nl = (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b0100) | (fsm_output[3])
      | (fsm_output[6]) | (fsm_output[9]) | not_tmp_51;
  assign mux_1349_nl = MUX_s_1_2_2(or_1004_nl, or_1003_nl, fsm_output[0]);
  assign mux_tmp_1350 = MUX_s_1_2_2(or_1005_nl, mux_1349_nl, fsm_output[5]);
  assign or_1013_nl = (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b010) | (VEC_LOOP_j_sva_11_0[0])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[9]) | (~ (fsm_output[8]))
      | (fsm_output[10]);
  assign or_1012_nl = (COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b0100) | (fsm_output[3])
      | (~ (fsm_output[6])) | (~ (fsm_output[9])) | (~ (fsm_output[8])) | (fsm_output[10]);
  assign mux_1353_nl = MUX_s_1_2_2(or_1013_nl, or_1012_nl, fsm_output[0]);
  assign or_1011_nl = (COMP_LOOP_acc_1_cse_sva[3:0]!=4'b0100) | (~ (fsm_output[0]))
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (~ (fsm_output[9])) | (fsm_output[8])
      | (~ (fsm_output[10]));
  assign mux_1354_nl = MUX_s_1_2_2(mux_1353_nl, or_1011_nl, fsm_output[5]);
  assign or_1009_nl = (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b010) | (~ (fsm_output[5]))
      | (fsm_output[0]) | (VEC_LOOP_j_sva_11_0[0]) | (fsm_output[3]) | (~ (fsm_output[6]))
      | (fsm_output[9]) | (fsm_output[8]) | (~ (fsm_output[10]));
  assign mux_tmp_1355 = MUX_s_1_2_2(mux_1354_nl, or_1009_nl, fsm_output[4]);
  assign or_1017_nl = (COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b0100) | (~ (fsm_output[0]))
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[9]) | (fsm_output[8])
      | (~ (fsm_output[10]));
  assign or_1015_nl = (~ (fsm_output[0])) | (fsm_output[3]) | (fsm_output[6]) | (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b0100)
      | (fsm_output[10:8]!=3'b001);
  assign mux_tmp_1356 = MUX_s_1_2_2(or_1017_nl, or_1015_nl, fsm_output[5]);
  assign or_tmp_1052 = (COMP_LOOP_acc_19_psp_sva[1:0]!=2'b01) | (fsm_output[0]) |
      (VEC_LOOP_j_sva_11_0[1:0]!=2'b01) | (~ (fsm_output[3])) | (fsm_output[6]) |
      (fsm_output[9]) | not_tmp_51;
  assign or_tmp_1056 = (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b0101) | (fsm_output[5])
      | (~ (fsm_output[0])) | (~ (fsm_output[3])) | (fsm_output[6]) | (fsm_output[9])
      | (fsm_output[8]) | (~ (fsm_output[10]));
  assign or_1119_nl = (VEC_LOOP_j_sva_11_0[3]) | (fsm_output[0]) | (VEC_LOOP_j_sva_11_0[2:0]!=3'b101)
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[9]) | (fsm_output[8]) | (fsm_output[10]);
  assign or_1118_nl = (COMP_LOOP_acc_16_psp_sva[0]) | (VEC_LOOP_j_sva_11_0[2:0]!=3'b101)
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[9])) | (~ (fsm_output[8]))
      | (fsm_output[10]);
  assign or_1117_nl = (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b0101) | (fsm_output[3])
      | (fsm_output[6]) | (fsm_output[9]) | not_tmp_51;
  assign mux_1426_nl = MUX_s_1_2_2(or_1118_nl, or_1117_nl, fsm_output[0]);
  assign mux_tmp_1427 = MUX_s_1_2_2(or_1119_nl, mux_1426_nl, fsm_output[5]);
  assign or_1135_nl = (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b010) | (~ (VEC_LOOP_j_sva_11_0[0]))
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[9]) | (~ (fsm_output[8]))
      | (fsm_output[10]);
  assign or_1134_nl = (COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b0101) | (fsm_output[3])
      | (~ (fsm_output[6])) | (~ (fsm_output[9])) | (~ (fsm_output[8])) | (fsm_output[10]);
  assign mux_1436_nl = MUX_s_1_2_2(or_1135_nl, or_1134_nl, fsm_output[0]);
  assign nand_432_nl = ~((COMP_LOOP_acc_1_cse_sva[3:0]==4'b0101) & (fsm_output[0])
      & (fsm_output[3]) & (fsm_output[6]) & (fsm_output[9]) & (~ (fsm_output[8]))
      & (fsm_output[10]));
  assign mux_1437_nl = MUX_s_1_2_2(mux_1436_nl, nand_432_nl, fsm_output[5]);
  assign or_1131_nl = (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b010) | (~ (fsm_output[5]))
      | (fsm_output[0]) | (~ (VEC_LOOP_j_sva_11_0[0])) | (fsm_output[3]) | (~ (fsm_output[6]))
      | (fsm_output[9]) | (fsm_output[8]) | (~ (fsm_output[10]));
  assign mux_tmp_1438 = MUX_s_1_2_2(mux_1437_nl, or_1131_nl, fsm_output[4]);
  assign or_1138_nl = (COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b0101) | (~ (fsm_output[0]))
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[9]) | (fsm_output[8])
      | (~ (fsm_output[10]));
  assign or_1136_nl = (~ (fsm_output[0])) | (fsm_output[3]) | (fsm_output[6]) | (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b0101)
      | (fsm_output[10:8]!=3'b001);
  assign mux_tmp_1440 = MUX_s_1_2_2(or_1138_nl, or_1136_nl, fsm_output[5]);
  assign or_tmp_1154 = (COMP_LOOP_acc_19_psp_sva[1:0]!=2'b01) | (fsm_output[0]) |
      (VEC_LOOP_j_sva_11_0[1:0]!=2'b10) | (~ (fsm_output[3])) | (fsm_output[6]) |
      (fsm_output[9]) | not_tmp_51;
  assign or_tmp_1157 = (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b0110) | (fsm_output[5])
      | (~ (fsm_output[0])) | (~ (fsm_output[3])) | (fsm_output[6]) | (fsm_output[9])
      | (fsm_output[8]) | (~ (fsm_output[10]));
  assign or_1218_nl = (VEC_LOOP_j_sva_11_0[3]) | (fsm_output[0]) | (VEC_LOOP_j_sva_11_0[2:0]!=3'b110)
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[9]) | (fsm_output[8]) | (fsm_output[10]);
  assign or_1217_nl = (COMP_LOOP_acc_16_psp_sva[0]) | (VEC_LOOP_j_sva_11_0[2:0]!=3'b110)
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[9])) | (~ (fsm_output[8]))
      | (fsm_output[10]);
  assign or_1216_nl = (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b0110) | (fsm_output[3])
      | (fsm_output[6]) | (fsm_output[9]) | not_tmp_51;
  assign mux_1493_nl = MUX_s_1_2_2(or_1217_nl, or_1216_nl, fsm_output[0]);
  assign mux_tmp_1494 = MUX_s_1_2_2(or_1218_nl, mux_1493_nl, fsm_output[5]);
  assign or_1226_nl = (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b011) | (VEC_LOOP_j_sva_11_0[0])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[9]) | (~ (fsm_output[8]))
      | (fsm_output[10]);
  assign or_1225_nl = (COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b0110) | (fsm_output[3])
      | (~ (fsm_output[6])) | (~ (fsm_output[9])) | (~ (fsm_output[8])) | (fsm_output[10]);
  assign mux_1497_nl = MUX_s_1_2_2(or_1226_nl, or_1225_nl, fsm_output[0]);
  assign nand_431_nl = ~((COMP_LOOP_acc_1_cse_sva[3:0]==4'b0110) & (fsm_output[0])
      & (fsm_output[3]) & (fsm_output[6]) & (fsm_output[9]) & (~ (fsm_output[8]))
      & (fsm_output[10]));
  assign mux_1498_nl = MUX_s_1_2_2(mux_1497_nl, nand_431_nl, fsm_output[5]);
  assign or_1222_nl = (~ (fsm_output[5])) | (fsm_output[0]) | (VEC_LOOP_j_sva_11_0[0])
      | (fsm_output[3]) | (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b011) | (~ (fsm_output[6]))
      | (fsm_output[9]) | (fsm_output[8]) | (~ (fsm_output[10]));
  assign mux_tmp_1499 = MUX_s_1_2_2(mux_1498_nl, or_1222_nl, fsm_output[4]);
  assign or_1230_nl = (COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b0110) | (~ (fsm_output[0]))
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[9]) | (fsm_output[8])
      | (~ (fsm_output[10]));
  assign or_1228_nl = (~ (fsm_output[0])) | (fsm_output[3]) | (fsm_output[6]) | (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b0110)
      | (fsm_output[10:8]!=3'b001);
  assign mux_tmp_1500 = MUX_s_1_2_2(or_1230_nl, or_1228_nl, fsm_output[5]);
  assign or_tmp_1265 = (COMP_LOOP_acc_19_psp_sva[1:0]!=2'b01) | (fsm_output[0]) |
      (VEC_LOOP_j_sva_11_0[1:0]!=2'b11) | (~ (fsm_output[3])) | (fsm_output[6]) |
      (fsm_output[9]) | not_tmp_51;
  assign or_tmp_1269 = (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b0111) | (fsm_output[5])
      | (~ (fsm_output[0])) | (~ (fsm_output[3])) | (fsm_output[6]) | (fsm_output[9])
      | (fsm_output[8]) | (~ (fsm_output[10]));
  assign or_1332_nl = (VEC_LOOP_j_sva_11_0[3]) | (fsm_output[0]) | (VEC_LOOP_j_sva_11_0[2:0]!=3'b111)
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[9]) | (fsm_output[8]) | (fsm_output[10]);
  assign or_1331_nl = (COMP_LOOP_acc_16_psp_sva[0]) | (VEC_LOOP_j_sva_11_0[2:0]!=3'b111)
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[9])) | (~ (fsm_output[8]))
      | (fsm_output[10]);
  assign or_1330_nl = (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b0111) | (fsm_output[3])
      | (fsm_output[6]) | (fsm_output[9]) | not_tmp_51;
  assign mux_1570_nl = MUX_s_1_2_2(or_1331_nl, or_1330_nl, fsm_output[0]);
  assign mux_tmp_1571 = MUX_s_1_2_2(or_1332_nl, mux_1570_nl, fsm_output[5]);
  assign or_1348_nl = (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b011) | (~ (VEC_LOOP_j_sva_11_0[0]))
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[9]) | (~ (fsm_output[8]))
      | (fsm_output[10]);
  assign or_1347_nl = (COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b0111) | (fsm_output[3])
      | (~ (fsm_output[6])) | (~ (fsm_output[9])) | (~ (fsm_output[8])) | (fsm_output[10]);
  assign mux_1580_nl = MUX_s_1_2_2(or_1348_nl, or_1347_nl, fsm_output[0]);
  assign nand_430_nl = ~((COMP_LOOP_acc_1_cse_sva[3:0]==4'b0111) & (fsm_output[0])
      & (fsm_output[3]) & (fsm_output[6]) & (fsm_output[9]) & (~ (fsm_output[8]))
      & (fsm_output[10]));
  assign mux_1581_nl = MUX_s_1_2_2(mux_1580_nl, nand_430_nl, fsm_output[5]);
  assign or_1344_nl = (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b011) | (~ (fsm_output[5]))
      | (fsm_output[0]) | (~ (VEC_LOOP_j_sva_11_0[0])) | (fsm_output[3]) | (~ (fsm_output[6]))
      | (fsm_output[9]) | (fsm_output[8]) | (~ (fsm_output[10]));
  assign mux_tmp_1582 = MUX_s_1_2_2(mux_1581_nl, or_1344_nl, fsm_output[4]);
  assign nand_418_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]==4'b0111) & (fsm_output[0])
      & (fsm_output[3]) & (fsm_output[6]) & (~ (fsm_output[9])) & (~ (fsm_output[8]))
      & (fsm_output[10]));
  assign or_1349_nl = (~ (fsm_output[0])) | (fsm_output[3]) | (fsm_output[6]) | (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b0111)
      | (fsm_output[10:8]!=3'b001);
  assign mux_tmp_1584 = MUX_s_1_2_2(nand_418_nl, or_1349_nl, fsm_output[5]);
  assign or_tmp_1367 = (COMP_LOOP_acc_19_psp_sva[1:0]!=2'b10) | (fsm_output[0]) |
      (VEC_LOOP_j_sva_11_0[1:0]!=2'b00) | (~ (fsm_output[3])) | (fsm_output[6]) |
      (fsm_output[9]) | not_tmp_51;
  assign or_tmp_1370 = (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b1000) | (fsm_output[5])
      | (~ (fsm_output[0])) | (~ (fsm_output[3])) | (fsm_output[6]) | (fsm_output[9])
      | (fsm_output[8]) | (~ (fsm_output[10]));
  assign or_1431_nl = (~ (VEC_LOOP_j_sva_11_0[3])) | (fsm_output[0]) | (VEC_LOOP_j_sva_11_0[2:0]!=3'b000)
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[9]) | (fsm_output[8]) | (fsm_output[10]);
  assign or_1430_nl = (~ (COMP_LOOP_acc_16_psp_sva[0])) | (VEC_LOOP_j_sva_11_0[2:0]!=3'b000)
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[9])) | (~ (fsm_output[8]))
      | (fsm_output[10]);
  assign or_1429_nl = (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b1000) | (fsm_output[3])
      | (fsm_output[6]) | (fsm_output[9]) | not_tmp_51;
  assign mux_1637_nl = MUX_s_1_2_2(or_1430_nl, or_1429_nl, fsm_output[0]);
  assign mux_tmp_1638 = MUX_s_1_2_2(or_1431_nl, mux_1637_nl, fsm_output[5]);
  assign or_1439_nl = (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b100) | (VEC_LOOP_j_sva_11_0[0])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[9]) | (~ (fsm_output[8]))
      | (fsm_output[10]);
  assign or_1438_nl = (COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b1000) | (fsm_output[3])
      | (~ (fsm_output[6])) | (~ (fsm_output[9])) | (~ (fsm_output[8])) | (fsm_output[10]);
  assign mux_1641_nl = MUX_s_1_2_2(or_1439_nl, or_1438_nl, fsm_output[0]);
  assign or_1437_nl = (COMP_LOOP_acc_1_cse_sva[3:0]!=4'b1000) | (~ (fsm_output[0]))
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (~ (fsm_output[9])) | (fsm_output[8])
      | (~ (fsm_output[10]));
  assign mux_1642_nl = MUX_s_1_2_2(mux_1641_nl, or_1437_nl, fsm_output[5]);
  assign or_1435_nl = (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b100) | (~ (fsm_output[5]))
      | (fsm_output[0]) | (VEC_LOOP_j_sva_11_0[0]) | (fsm_output[3]) | (~ (fsm_output[6]))
      | (fsm_output[9]) | (fsm_output[8]) | (~ (fsm_output[10]));
  assign mux_tmp_1643 = MUX_s_1_2_2(mux_1642_nl, or_1435_nl, fsm_output[4]);
  assign or_1443_nl = (COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b1000) | (~ (fsm_output[0]))
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[9]) | (fsm_output[8])
      | (~ (fsm_output[10]));
  assign or_1441_nl = (~ (fsm_output[0])) | (fsm_output[3]) | (fsm_output[6]) | (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b1000)
      | (fsm_output[10:8]!=3'b001);
  assign mux_tmp_1644 = MUX_s_1_2_2(or_1443_nl, or_1441_nl, fsm_output[5]);
  assign or_tmp_1478 = (COMP_LOOP_acc_19_psp_sva[1:0]!=2'b10) | (fsm_output[0]) |
      (VEC_LOOP_j_sva_11_0[1:0]!=2'b01) | (~ (fsm_output[3])) | (fsm_output[6]) |
      (fsm_output[9]) | not_tmp_51;
  assign or_tmp_1482 = (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b1001) | (fsm_output[5])
      | (~ (fsm_output[0])) | (~ (fsm_output[3])) | (fsm_output[6]) | (fsm_output[9])
      | (fsm_output[8]) | (~ (fsm_output[10]));
  assign or_1545_nl = (~ (VEC_LOOP_j_sva_11_0[3])) | (fsm_output[0]) | (VEC_LOOP_j_sva_11_0[2:0]!=3'b001)
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[9]) | (fsm_output[8]) | (fsm_output[10]);
  assign or_1544_nl = (~ (COMP_LOOP_acc_16_psp_sva[0])) | (VEC_LOOP_j_sva_11_0[2:0]!=3'b001)
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[9])) | (~ (fsm_output[8]))
      | (fsm_output[10]);
  assign or_1543_nl = (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b1001) | (fsm_output[3])
      | (fsm_output[6]) | (fsm_output[9]) | not_tmp_51;
  assign mux_1714_nl = MUX_s_1_2_2(or_1544_nl, or_1543_nl, fsm_output[0]);
  assign mux_tmp_1715 = MUX_s_1_2_2(or_1545_nl, mux_1714_nl, fsm_output[5]);
  assign or_1561_nl = (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b100) | (~ (VEC_LOOP_j_sva_11_0[0]))
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[9]) | (~ (fsm_output[8]))
      | (fsm_output[10]);
  assign or_1560_nl = (COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b1001) | (fsm_output[3])
      | (~ (fsm_output[6])) | (~ (fsm_output[9])) | (~ (fsm_output[8])) | (fsm_output[10]);
  assign mux_1724_nl = MUX_s_1_2_2(or_1561_nl, or_1560_nl, fsm_output[0]);
  assign nand_429_nl = ~((COMP_LOOP_acc_1_cse_sva[3:0]==4'b1001) & (fsm_output[0])
      & (fsm_output[3]) & (fsm_output[6]) & (fsm_output[9]) & (~ (fsm_output[8]))
      & (fsm_output[10]));
  assign mux_1725_nl = MUX_s_1_2_2(mux_1724_nl, nand_429_nl, fsm_output[5]);
  assign or_1557_nl = (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b100) | (~ (fsm_output[5]))
      | (fsm_output[0]) | (~ (VEC_LOOP_j_sva_11_0[0])) | (fsm_output[3]) | (~ (fsm_output[6]))
      | (fsm_output[9]) | (fsm_output[8]) | (~ (fsm_output[10]));
  assign mux_tmp_1726 = MUX_s_1_2_2(mux_1725_nl, or_1557_nl, fsm_output[4]);
  assign or_1564_nl = (COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b1001) | (~ (fsm_output[0]))
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[9]) | (fsm_output[8])
      | (~ (fsm_output[10]));
  assign or_1562_nl = (~ (fsm_output[0])) | (fsm_output[3]) | (fsm_output[6]) | (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b1001)
      | (fsm_output[10:8]!=3'b001);
  assign mux_tmp_1728 = MUX_s_1_2_2(or_1564_nl, or_1562_nl, fsm_output[5]);
  assign or_tmp_1580 = (COMP_LOOP_acc_19_psp_sva[1:0]!=2'b10) | (fsm_output[0]) |
      (VEC_LOOP_j_sva_11_0[1:0]!=2'b10) | (~ (fsm_output[3])) | (fsm_output[6]) |
      (fsm_output[9]) | not_tmp_51;
  assign or_tmp_1583 = (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b1010) | (fsm_output[5])
      | (~ (fsm_output[0])) | (~ (fsm_output[3])) | (fsm_output[6]) | (fsm_output[9])
      | (fsm_output[8]) | (~ (fsm_output[10]));
  assign or_1644_nl = (~ (VEC_LOOP_j_sva_11_0[3])) | (fsm_output[0]) | (VEC_LOOP_j_sva_11_0[2:0]!=3'b010)
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[9]) | (fsm_output[8]) | (fsm_output[10]);
  assign or_1643_nl = (~ (COMP_LOOP_acc_16_psp_sva[0])) | (VEC_LOOP_j_sva_11_0[2:0]!=3'b010)
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[9])) | (~ (fsm_output[8]))
      | (fsm_output[10]);
  assign or_1642_nl = (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b1010) | (fsm_output[3])
      | (fsm_output[6]) | (fsm_output[9]) | not_tmp_51;
  assign mux_1781_nl = MUX_s_1_2_2(or_1643_nl, or_1642_nl, fsm_output[0]);
  assign mux_tmp_1782 = MUX_s_1_2_2(or_1644_nl, mux_1781_nl, fsm_output[5]);
  assign or_1652_nl = (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b101) | (VEC_LOOP_j_sva_11_0[0])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[9]) | (~ (fsm_output[8]))
      | (fsm_output[10]);
  assign or_1651_nl = (COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b1010) | (fsm_output[3])
      | (~ (fsm_output[6])) | (~ (fsm_output[9])) | (~ (fsm_output[8])) | (fsm_output[10]);
  assign mux_1785_nl = MUX_s_1_2_2(or_1652_nl, or_1651_nl, fsm_output[0]);
  assign nand_428_nl = ~((COMP_LOOP_acc_1_cse_sva[3:0]==4'b1010) & (fsm_output[0])
      & (fsm_output[3]) & (fsm_output[6]) & (fsm_output[9]) & (~ (fsm_output[8]))
      & (fsm_output[10]));
  assign mux_1786_nl = MUX_s_1_2_2(mux_1785_nl, nand_428_nl, fsm_output[5]);
  assign or_1648_nl = (~ (fsm_output[5])) | (fsm_output[0]) | (VEC_LOOP_j_sva_11_0[0])
      | (fsm_output[3]) | (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b101) | (~ (fsm_output[6]))
      | (fsm_output[9]) | (fsm_output[8]) | (~ (fsm_output[10]));
  assign mux_tmp_1787 = MUX_s_1_2_2(mux_1786_nl, or_1648_nl, fsm_output[4]);
  assign or_1656_nl = (COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b1010) | (~ (fsm_output[0]))
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[9]) | (fsm_output[8])
      | (~ (fsm_output[10]));
  assign or_1654_nl = (~ (fsm_output[0])) | (fsm_output[3]) | (fsm_output[6]) | (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b1010)
      | (fsm_output[10:8]!=3'b001);
  assign mux_tmp_1788 = MUX_s_1_2_2(or_1656_nl, or_1654_nl, fsm_output[5]);
  assign or_tmp_1691 = (COMP_LOOP_acc_19_psp_sva[1:0]!=2'b10) | (fsm_output[0]) |
      (VEC_LOOP_j_sva_11_0[1:0]!=2'b11) | (~ (fsm_output[3])) | (fsm_output[6]) |
      (fsm_output[9]) | not_tmp_51;
  assign or_tmp_1695 = (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b1011) | (fsm_output[5])
      | (~ (fsm_output[0])) | (~ (fsm_output[3])) | (fsm_output[6]) | (fsm_output[9])
      | (fsm_output[8]) | (~ (fsm_output[10]));
  assign or_1758_nl = (~ (VEC_LOOP_j_sva_11_0[3])) | (fsm_output[0]) | (VEC_LOOP_j_sva_11_0[2:0]!=3'b011)
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[9]) | (fsm_output[8]) | (fsm_output[10]);
  assign or_1757_nl = (~ (COMP_LOOP_acc_16_psp_sva[0])) | (VEC_LOOP_j_sva_11_0[2:0]!=3'b011)
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[9])) | (~ (fsm_output[8]))
      | (fsm_output[10]);
  assign or_1756_nl = (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b1011) | (fsm_output[3])
      | (fsm_output[6]) | (fsm_output[9]) | not_tmp_51;
  assign mux_1858_nl = MUX_s_1_2_2(or_1757_nl, or_1756_nl, fsm_output[0]);
  assign mux_tmp_1859 = MUX_s_1_2_2(or_1758_nl, mux_1858_nl, fsm_output[5]);
  assign or_1774_nl = (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b101) | (~ (VEC_LOOP_j_sva_11_0[0]))
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[9]) | (~ (fsm_output[8]))
      | (fsm_output[10]);
  assign or_1773_nl = (COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b1011) | (fsm_output[3])
      | (~ (fsm_output[6])) | (~ (fsm_output[9])) | (~ (fsm_output[8])) | (fsm_output[10]);
  assign mux_1868_nl = MUX_s_1_2_2(or_1774_nl, or_1773_nl, fsm_output[0]);
  assign nand_427_nl = ~((COMP_LOOP_acc_1_cse_sva[3:0]==4'b1011) & (fsm_output[0])
      & (fsm_output[3]) & (fsm_output[6]) & (fsm_output[9]) & (~ (fsm_output[8]))
      & (fsm_output[10]));
  assign mux_1869_nl = MUX_s_1_2_2(mux_1868_nl, nand_427_nl, fsm_output[5]);
  assign or_1770_nl = (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b101) | (~ (fsm_output[5]))
      | (fsm_output[0]) | (~ (VEC_LOOP_j_sva_11_0[0])) | (fsm_output[3]) | (~ (fsm_output[6]))
      | (fsm_output[9]) | (fsm_output[8]) | (~ (fsm_output[10]));
  assign mux_tmp_1870 = MUX_s_1_2_2(mux_1869_nl, or_1770_nl, fsm_output[4]);
  assign nand_416_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]==4'b1011) & (fsm_output[0])
      & (fsm_output[3]) & (fsm_output[6]) & (~ (fsm_output[9])) & (~ (fsm_output[8]))
      & (fsm_output[10]));
  assign or_1775_nl = (~ (fsm_output[0])) | (fsm_output[3]) | (fsm_output[6]) | (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b1011)
      | (fsm_output[10:8]!=3'b001);
  assign mux_tmp_1872 = MUX_s_1_2_2(nand_416_nl, or_1775_nl, fsm_output[5]);
  assign or_1853_nl = (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b11) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b00)
      | (~ (fsm_output[4])) | (~ (fsm_output[9])) | (fsm_output[3]) | (fsm_output[6])
      | (fsm_output[10]);
  assign or_1852_nl = (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b1100) | (fsm_output[4])
      | (fsm_output[9]) | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[10]));
  assign mux_1922_nl = MUX_s_1_2_2(or_1853_nl, or_1852_nl, fsm_output[0]);
  assign or_tmp_1797 = (fsm_output[5]) | mux_1922_nl;
  assign not_tmp_378 = ~((fsm_output[6]) & (fsm_output[10]));
  assign nor_874_nl = ~((COMP_LOOP_acc_17_psp_sva[2:0]!=3'b110) | (VEC_LOOP_j_sva_11_0[0])
      | (~ (fsm_output[4])) | (fsm_output[9]) | (fsm_output[3]) | not_tmp_378);
  assign nor_875_nl = ~((COMP_LOOP_acc_1_cse_sva[3:0]!=4'b1100) | (fsm_output[4])
      | (~((fsm_output[9]) & (fsm_output[3]) & (fsm_output[6]) & (fsm_output[10]))));
  assign mux_1926_nl = MUX_s_1_2_2(nor_874_nl, nor_875_nl, fsm_output[0]);
  assign nand_73_nl = ~((fsm_output[5]) & mux_1926_nl);
  assign or_1856_nl = (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b110) | (VEC_LOOP_j_sva_11_0[0])
      | (fsm_output[4]) | (fsm_output[9]) | (~ (fsm_output[3])) | (~ (fsm_output[6]))
      | (fsm_output[10]);
  assign or_1855_nl = (COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b1100) | (fsm_output[4])
      | (~ (fsm_output[9])) | (fsm_output[3]) | (~ (fsm_output[6])) | (fsm_output[10]);
  assign mux_1925_nl = MUX_s_1_2_2(or_1856_nl, or_1855_nl, fsm_output[0]);
  assign or_1857_nl = (fsm_output[5]) | mux_1925_nl;
  assign mux_tmp_1927 = MUX_s_1_2_2(nand_73_nl, or_1857_nl, fsm_output[8]);
  assign nor_872_nl = ~((~ (COMP_LOOP_acc_16_psp_sva[0])) | (VEC_LOOP_j_sva_11_0[2:0]!=3'b100)
      | (fsm_output[4]) | (~ (fsm_output[9])) | (~ (fsm_output[3])) | (fsm_output[6])
      | (fsm_output[10]));
  assign nor_873_nl = ~((COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b1100) | (fsm_output[4])
      | (fsm_output[9]) | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[10])));
  assign mux_1929_nl = MUX_s_1_2_2(nor_872_nl, nor_873_nl, fsm_output[0]);
  assign nand_tmp_74 = ~((fsm_output[5]) & mux_1929_nl);
  assign or_tmp_1811 = (~ (fsm_output[5])) | (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b1100)
      | (~ (fsm_output[0])) | (~ (fsm_output[4])) | (fsm_output[9]) | (fsm_output[3])
      | (fsm_output[6]) | (fsm_output[10]);
  assign or_tmp_1812 = (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b110) | (fsm_output[0])
      | (VEC_LOOP_j_sva_11_0[0]) | (fsm_output[4]) | (~ (fsm_output[9])) | (fsm_output[3])
      | (~ (fsm_output[6])) | (fsm_output[10]);
  assign not_tmp_381 = ~((fsm_output[3]) & (fsm_output[6]) & (fsm_output[10]));
  assign or_tmp_1821 = (fsm_output[4]) | (fsm_output[9]) | (fsm_output[3]) | (fsm_output[6])
      | (~ (fsm_output[10]));
  assign or_tmp_1907 = (COMP_LOOP_acc_19_psp_sva[1:0]!=2'b11) | (fsm_output[0]) |
      (VEC_LOOP_j_sva_11_0[1:0]!=2'b01) | (~ (fsm_output[3])) | (fsm_output[6]) |
      (fsm_output[9]) | not_tmp_51;
  assign or_tmp_1911 = (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b1101) | (fsm_output[5])
      | (~ (fsm_output[0])) | (~ (fsm_output[3])) | (fsm_output[6]) | (fsm_output[9])
      | (fsm_output[8]) | (~ (fsm_output[10]));
  assign or_1974_nl = (~ (VEC_LOOP_j_sva_11_0[3])) | (fsm_output[0]) | (VEC_LOOP_j_sva_11_0[2:0]!=3'b101)
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[9]) | (fsm_output[8]) | (fsm_output[10]);
  assign or_1973_nl = (~ (COMP_LOOP_acc_16_psp_sva[0])) | (VEC_LOOP_j_sva_11_0[2:0]!=3'b101)
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[9])) | (~ (fsm_output[8]))
      | (fsm_output[10]);
  assign or_1972_nl = (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b1101) | (fsm_output[3])
      | (fsm_output[6]) | (fsm_output[9]) | not_tmp_51;
  assign mux_2003_nl = MUX_s_1_2_2(or_1973_nl, or_1972_nl, fsm_output[0]);
  assign mux_tmp_2004 = MUX_s_1_2_2(or_1974_nl, mux_2003_nl, fsm_output[5]);
  assign or_1990_nl = (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b110) | (~ (VEC_LOOP_j_sva_11_0[0]))
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[9]) | (~ (fsm_output[8]))
      | (fsm_output[10]);
  assign or_1989_nl = (COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b1101) | (fsm_output[3])
      | (~ (fsm_output[6])) | (~ (fsm_output[9])) | (~ (fsm_output[8])) | (fsm_output[10]);
  assign mux_2013_nl = MUX_s_1_2_2(or_1990_nl, or_1989_nl, fsm_output[0]);
  assign nand_426_nl = ~((COMP_LOOP_acc_1_cse_sva[3:0]==4'b1101) & (fsm_output[0])
      & (fsm_output[3]) & (fsm_output[6]) & (fsm_output[9]) & (~ (fsm_output[8]))
      & (fsm_output[10]));
  assign mux_2014_nl = MUX_s_1_2_2(mux_2013_nl, nand_426_nl, fsm_output[5]);
  assign or_1986_nl = (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b110) | (~ (fsm_output[5]))
      | (fsm_output[0]) | (~ (VEC_LOOP_j_sva_11_0[0])) | (fsm_output[3]) | (~ (fsm_output[6]))
      | (fsm_output[9]) | (fsm_output[8]) | (~ (fsm_output[10]));
  assign mux_tmp_2015 = MUX_s_1_2_2(mux_2014_nl, or_1986_nl, fsm_output[4]);
  assign nand_414_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]==4'b1101) & (fsm_output[0])
      & (fsm_output[3]) & (fsm_output[6]) & (~ (fsm_output[9])) & (~ (fsm_output[8]))
      & (fsm_output[10]));
  assign or_1991_nl = (~ (fsm_output[0])) | (fsm_output[3]) | (fsm_output[6]) | (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b1101)
      | (fsm_output[10:8]!=3'b001);
  assign mux_tmp_2017 = MUX_s_1_2_2(nand_414_nl, or_1991_nl, fsm_output[5]);
  assign or_tmp_2009 = (COMP_LOOP_acc_19_psp_sva[1:0]!=2'b11) | (fsm_output[0]) |
      (VEC_LOOP_j_sva_11_0[1:0]!=2'b10) | (~ (fsm_output[3])) | (fsm_output[6]) |
      (fsm_output[9]) | not_tmp_51;
  assign or_tmp_2012 = (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b1110) | (fsm_output[5])
      | (~ (fsm_output[0])) | (~ (fsm_output[3])) | (fsm_output[6]) | (fsm_output[9])
      | (fsm_output[8]) | (~ (fsm_output[10]));
  assign or_2073_nl = (~ (VEC_LOOP_j_sva_11_0[3])) | (fsm_output[0]) | (VEC_LOOP_j_sva_11_0[2:0]!=3'b110)
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[9]) | (fsm_output[8]) | (fsm_output[10]);
  assign or_2072_nl = (~ (COMP_LOOP_acc_16_psp_sva[0])) | (VEC_LOOP_j_sva_11_0[2:0]!=3'b110)
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[9])) | (~ (fsm_output[8]))
      | (fsm_output[10]);
  assign or_2071_nl = (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b1110) | (fsm_output[3])
      | (fsm_output[6]) | (fsm_output[9]) | not_tmp_51;
  assign mux_2070_nl = MUX_s_1_2_2(or_2072_nl, or_2071_nl, fsm_output[0]);
  assign mux_tmp_2071 = MUX_s_1_2_2(or_2073_nl, mux_2070_nl, fsm_output[5]);
  assign or_2081_nl = (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b111) | (VEC_LOOP_j_sva_11_0[0])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[9]) | (~ (fsm_output[8]))
      | (fsm_output[10]);
  assign or_2080_nl = (COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b1110) | (fsm_output[3])
      | (~ (fsm_output[6])) | (~ (fsm_output[9])) | (~ (fsm_output[8])) | (fsm_output[10]);
  assign mux_2074_nl = MUX_s_1_2_2(or_2081_nl, or_2080_nl, fsm_output[0]);
  assign nand_425_nl = ~((COMP_LOOP_acc_1_cse_sva[3:0]==4'b1110) & (fsm_output[0])
      & (fsm_output[3]) & (fsm_output[6]) & (fsm_output[9]) & (~ (fsm_output[8]))
      & (fsm_output[10]));
  assign mux_2075_nl = MUX_s_1_2_2(mux_2074_nl, nand_425_nl, fsm_output[5]);
  assign or_2077_nl = (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b111) | (~ (fsm_output[5]))
      | (fsm_output[0]) | (VEC_LOOP_j_sva_11_0[0]) | (fsm_output[3]) | (~ (fsm_output[6]))
      | (fsm_output[9]) | (fsm_output[8]) | (~ (fsm_output[10]));
  assign mux_tmp_2076 = MUX_s_1_2_2(mux_2075_nl, or_2077_nl, fsm_output[4]);
  assign nand_412_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]==4'b1110) & (fsm_output[0])
      & (fsm_output[3]) & (fsm_output[6]) & (~ (fsm_output[9])) & (~ (fsm_output[8]))
      & (fsm_output[10]));
  assign or_2083_nl = (~ (fsm_output[0])) | (fsm_output[3]) | (fsm_output[6]) | (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b1110)
      | (fsm_output[10:8]!=3'b001);
  assign mux_tmp_2077 = MUX_s_1_2_2(nand_412_nl, or_2083_nl, fsm_output[5]);
  assign or_tmp_2120 = (COMP_LOOP_acc_19_psp_sva[1:0]!=2'b11) | (fsm_output[0]) |
      (VEC_LOOP_j_sva_11_0[1:0]!=2'b11) | (~ (fsm_output[3])) | (fsm_output[6]) |
      (fsm_output[9]) | not_tmp_51;
  assign or_tmp_2124 = (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b1111) | (fsm_output[5])
      | (~ (fsm_output[0])) | (~ (fsm_output[3])) | (fsm_output[6]) | (fsm_output[9])
      | (fsm_output[8]) | (~ (fsm_output[10]));
  assign or_2187_nl = (~ (VEC_LOOP_j_sva_11_0[3])) | (fsm_output[0]) | (VEC_LOOP_j_sva_11_0[2:0]!=3'b111)
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[9]) | (fsm_output[8]) | (fsm_output[10]);
  assign nand_291_nl = ~((COMP_LOOP_acc_16_psp_sva[0]) & (VEC_LOOP_j_sva_11_0[2:0]==3'b111)
      & (fsm_output[3]) & (~ (fsm_output[6])) & (fsm_output[9]) & (fsm_output[8])
      & (~ (fsm_output[10])));
  assign or_2185_nl = (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b1111) | (fsm_output[3])
      | (fsm_output[6]) | (fsm_output[9]) | not_tmp_51;
  assign mux_2147_nl = MUX_s_1_2_2(nand_291_nl, or_2185_nl, fsm_output[0]);
  assign mux_tmp_2148 = MUX_s_1_2_2(or_2187_nl, mux_2147_nl, fsm_output[5]);
  assign nand_288_nl = ~((COMP_LOOP_acc_11_psp_sva[2:0]==3'b111) & (VEC_LOOP_j_sva_11_0[0])
      & (fsm_output[3]) & (fsm_output[6]) & (~ (fsm_output[9])) & (fsm_output[8])
      & (~ (fsm_output[10])));
  assign nand_289_nl = ~((~ (fsm_output[3])) & (COMP_LOOP_acc_1_cse_8_sva[3:0]==4'b1111)
      & (fsm_output[6]) & (fsm_output[9]) & (fsm_output[8]) & (~ (fsm_output[10])));
  assign mux_2157_nl = MUX_s_1_2_2(nand_288_nl, nand_289_nl, fsm_output[0]);
  assign nand_424_nl = ~((COMP_LOOP_acc_1_cse_sva[3:0]==4'b1111) & (fsm_output[0])
      & (fsm_output[3]) & (fsm_output[6]) & (fsm_output[9]) & (~ (fsm_output[8]))
      & (fsm_output[10]));
  assign mux_2158_nl = MUX_s_1_2_2(mux_2157_nl, nand_424_nl, fsm_output[5]);
  assign or_2199_nl = (~ (fsm_output[5])) | (fsm_output[0]) | (~ (VEC_LOOP_j_sva_11_0[0]))
      | (fsm_output[3]) | (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b111) | (~ (fsm_output[6]))
      | (fsm_output[9]) | (fsm_output[8]) | (~ (fsm_output[10]));
  assign mux_tmp_2159 = MUX_s_1_2_2(mux_2158_nl, or_2199_nl, fsm_output[4]);
  assign nand_410_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]==4'b1111) & (fsm_output[0])
      & (fsm_output[3]) & (fsm_output[6]) & (~ (fsm_output[9])) & (~ (fsm_output[8]))
      & (fsm_output[10]));
  assign or_2204_nl = (~ (fsm_output[0])) | (fsm_output[3]) | (fsm_output[6]) | (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b1111)
      | (fsm_output[10:8]!=3'b001);
  assign mux_tmp_2161 = MUX_s_1_2_2(nand_410_nl, or_2204_nl, fsm_output[5]);
  assign and_dcpl_260 = and_dcpl_124 & and_dcpl_100 & and_dcpl_98;
  assign nor_784_cse = ~((fsm_output[1:0]!=2'b00));
  assign or_tmp_2220 = nor_784_cse | (~ (fsm_output[3])) | (fsm_output[10]);
  assign or_tmp_2223 = (fsm_output[6]) | (fsm_output[3]) | (fsm_output[10]);
  assign or_tmp_2225 = (~(and_573_cse | (fsm_output[3]))) | (fsm_output[10]);
  assign or_tmp_2230 = and_573_cse | (fsm_output[3]) | (fsm_output[10]);
  assign or_tmp_2233 = ((fsm_output[3]) & (fsm_output[0]) & (fsm_output[1])) | (fsm_output[10]);
  assign mux_tmp_2218 = MUX_s_1_2_2((~ or_tmp_2233), or_tmp_21, fsm_output[6]);
  assign mux_tmp_2220 = MUX_s_1_2_2(and_dcpl_102, nor_tmp_6, fsm_output[6]);
  assign mux_tmp_2223 = MUX_s_1_2_2((~ nor_tmp_9), or_tmp_2233, fsm_output[6]);
  assign or_tmp_2237 = ~((fsm_output[6]) & (fsm_output[1]) & (fsm_output[3]) & (~
      (fsm_output[10])));
  assign or_tmp_2238 = (fsm_output[0]) | (fsm_output[1]) | (fsm_output[3]) | (fsm_output[10]);
  assign mux_tmp_2239 = MUX_s_1_2_2((~ (fsm_output[10])), (fsm_output[10]), fsm_output[3]);
  assign mux_2240_nl = MUX_s_1_2_2(and_dcpl_101, mux_tmp_2239, or_2348_cse);
  assign nand_tmp_92 = ~((fsm_output[6]) & (~ mux_2240_nl));
  assign nor_tmp_286 = or_2898_cse & (fsm_output[10]);
  assign or_tmp_2246 = (fsm_output[6]) | (~ (fsm_output[3])) | (fsm_output[10]);
  assign or_tmp_2248 = (or_2348_cse & (fsm_output[3])) | (fsm_output[10]);
  assign not_tmp_426 = ~((fsm_output[6]) & or_tmp_2248);
  assign nor_tmp_288 = ((fsm_output[3]) | (fsm_output[1])) & (fsm_output[10]);
  assign and_tmp_10 = (fsm_output[6]) & nor_tmp_288;
  assign mux_tmp_2250 = MUX_s_1_2_2(mux_tmp_2239, nor_tmp_6, or_2348_cse);
  assign mux_tmp_2251 = MUX_s_1_2_2(and_dcpl_101, mux_tmp_2239, fsm_output[1]);
  assign mux_tmp_2254 = MUX_s_1_2_2(and_dcpl_101, mux_tmp_2239, and_573_cse);
  assign or_tmp_2253 = ((fsm_output[3]) & (fsm_output[1])) | (fsm_output[10]);
  assign or_tmp_2255 = (fsm_output[6]) | or_tmp_2253;
  assign mux_tmp_2265 = MUX_s_1_2_2(and_dcpl_109, (fsm_output[10]), fsm_output[6]);
  assign nor_tmp_291 = or_2348_cse & (fsm_output[3]) & (fsm_output[10]);
  assign or_tmp_2257 = (fsm_output[6]) | or_tmp_2248;
  assign nor_tmp_295 = or_2902_cse & (fsm_output[10]);
  assign mux_tmp_2285 = MUX_s_1_2_2((~ nor_tmp_288), (fsm_output[10]), fsm_output[6]);
  assign mux_2289_nl = MUX_s_1_2_2(and_dcpl_101, or_tmp_2230, fsm_output[6]);
  assign mux_tmp_2290 = MUX_s_1_2_2(not_tmp_378, mux_2289_nl, fsm_output[7]);
  assign or_tmp_2260 = (fsm_output[3]) | (~ (fsm_output[10]));
  assign or_tmp_2263 = (fsm_output[7]) | (~ (fsm_output[6])) | (fsm_output[10]);
  assign nand_tmp_93 = ~((fsm_output[6]) & (~ or_tmp_2230));
  assign or_tmp_2266 = (fsm_output[1]) | (~ mux_tmp_2239);
  assign mux_tmp_2309 = MUX_s_1_2_2(mux_tmp_2239, nor_tmp_6, fsm_output[1]);
  assign mux_2310_nl = MUX_s_1_2_2(mux_tmp_2309, (~ or_tmp_2266), fsm_output[0]);
  assign or_tmp_2267 = (fsm_output[6]) | mux_2310_nl;
  assign or_tmp_2269 = (~((~ (fsm_output[0])) | (~ (fsm_output[1])) | (fsm_output[3])))
      | (fsm_output[10]);
  assign nand_tmp_95 = ~((fsm_output[6]) & (~ or_tmp_2269));
  assign or_tmp_2271 = (~((fsm_output[1]) | (fsm_output[3]))) | (fsm_output[10]);
  assign nand_tmp_96 = ~((fsm_output[6]) & (~ or_tmp_2253));
  assign or_tmp_2275 = (~((fsm_output[3]) | (fsm_output[0]) | (fsm_output[1]))) |
      (fsm_output[10]);
  assign or_tmp_2276 = (fsm_output[6]) | (~ (fsm_output[1])) | (~ (fsm_output[3]))
      | (fsm_output[10]);
  assign or_tmp_2277 = (fsm_output[0]) | (fsm_output[1]) | (~ (fsm_output[3])) |
      (fsm_output[10]);
  assign mux_tmp_2327 = MUX_s_1_2_2(or_tmp_2277, nor_tmp_291, fsm_output[6]);
  assign or_tmp_2280 = (fsm_output[6]) | (~ or_tmp_2220);
  assign or_tmp_2281 = (fsm_output[6]) | and_dcpl_110;
  assign or_tmp_2282 = (~ (fsm_output[1])) | (~ (fsm_output[3])) | (fsm_output[10]);
  assign or_tmp_2289 = nor_784_cse | (fsm_output[3]) | (~ (fsm_output[10]));
  assign not_tmp_463 = ~((fsm_output[6]) & or_tmp_2289);
  assign mux_tmp_2349 = MUX_s_1_2_2((~ or_tmp_2248), or_tmp_21, fsm_output[6]);
  assign and_tmp_16 = (fsm_output[6]) & or_tmp_2282;
  assign or_tmp_2293 = (fsm_output[6]) | (~ nor_tmp_295);
  assign mux_tmp_2362 = MUX_s_1_2_2(mux_tmp_2239, nor_tmp_6, and_573_cse);
  assign nor_tmp_300 = (fsm_output[0]) & (fsm_output[1]) & (fsm_output[3]) & (fsm_output[10]);
  assign or_tmp_2327 = ~((fsm_output[5]) & (fsm_output[8]) & (fsm_output[6]) & (~
      (fsm_output[10])));
  assign or_tmp_2329 = (fsm_output[5]) | (fsm_output[8]) | (~ (fsm_output[6])) |
      (fsm_output[10]);
  assign or_tmp_2331 = (fsm_output[5]) | (fsm_output[8]) | (~ (fsm_output[6]));
  assign or_tmp_2333 = (~ (fsm_output[8])) | (~ (fsm_output[6])) | (fsm_output[10]);
  assign or_tmp_2334 = (~ (fsm_output[8])) | (fsm_output[6]) | (fsm_output[10]);
  assign mux_tmp_2400 = MUX_s_1_2_2(or_tmp_2334, or_tmp_2333, fsm_output[5]);
  assign mux_tmp_2401 = MUX_s_1_2_2(or_tmp_4, or_tmp_14, fsm_output[8]);
  assign mux_tmp_2402 = MUX_s_1_2_2(mux_tmp_2401, or_tmp_2333, fsm_output[5]);
  assign or_tmp_2335 = (fsm_output[5]) | mux_tmp_2401;
  assign or_2393_nl = (fsm_output[8]) | not_tmp_378;
  assign mux_tmp_2406 = MUX_s_1_2_2(or_2393_nl, or_tmp_2334, fsm_output[5]);
  assign or_tmp_2338 = (fsm_output[5]) | (fsm_output[8]) | not_tmp_378;
  assign nand_tmp_105 = ~((fsm_output[5]) & (~ mux_tmp_2401));
  assign mux_tmp_2423 = MUX_s_1_2_2(or_tmp_2334, mux_tmp_917, fsm_output[5]);
  assign nor_tmp_307 = (fsm_output[8]) & (fsm_output[6]) & (fsm_output[10]);
  assign mux_tmp_2425 = MUX_s_1_2_2((~ (fsm_output[6])), or_tmp_434, fsm_output[8]);
  assign mux_tmp_2426 = MUX_s_1_2_2((~ mux_tmp_2425), nor_tmp_307, fsm_output[5]);
  assign or_tmp_2342 = (fsm_output[5]) | mux_tmp_2425;
  assign mux_2427_nl = MUX_s_1_2_2(not_tmp_378, or_tmp_434, fsm_output[8]);
  assign or_tmp_2343 = (fsm_output[5]) | mux_2427_nl;
  assign mux_2433_itm = MUX_s_1_2_2(or_tmp_4, (fsm_output[6]), fsm_output[8]);
  assign mux_2435_itm = MUX_s_1_2_2(or_tmp_4, or_tmp_434, fsm_output[8]);
  assign mux_tmp_2436 = MUX_s_1_2_2((~ mux_2435_itm), nor_tmp_307, fsm_output[5]);
  assign nand_tmp_107 = ~((fsm_output[5]) & (~ mux_2433_itm));
  assign nand_tmp_108 = ~((fsm_output[5]) & (~ mux_2435_itm));
  assign or_2415_cse = (fsm_output[9]) | (fsm_output[4]) | (~ (fsm_output[10]));
  assign mux_tmp_2466 = MUX_s_1_2_2(or_tmp_195, or_2415_cse, fsm_output[1]);
  assign or_2409_nl = (~ (fsm_output[3])) | (~ (fsm_output[1])) | (fsm_output[9])
      | (~ (fsm_output[4])) | (fsm_output[10]);
  assign mux_2463_cse = MUX_s_1_2_2(or_2409_nl, or_2824_cse, fsm_output[0]);
  assign or_2425_nl = (fsm_output[5]) | (fsm_output[2]) | (~ (fsm_output[0])) | (fsm_output[3])
      | (~ (fsm_output[1])) | (~ (fsm_output[9])) | (fsm_output[4]) | (fsm_output[10]);
  assign or_2424_nl = (fsm_output[2]) | (fsm_output[0]) | nand_226_cse;
  assign mux_2470_nl = MUX_s_1_2_2(or_529_cse, or_2826_cse, fsm_output[0]);
  assign mux_2471_nl = MUX_s_1_2_2(mux_2470_nl, or_2839_cse, fsm_output[2]);
  assign mux_2472_nl = MUX_s_1_2_2(or_2424_nl, mux_2471_nl, fsm_output[5]);
  assign mux_2473_nl = MUX_s_1_2_2(or_2425_nl, mux_2472_nl, fsm_output[6]);
  assign or_2419_nl = (fsm_output[3]) | mux_tmp_2466;
  assign mux_2469_nl = MUX_s_1_2_2(or_2419_nl, or_529_cse, fsm_output[0]);
  assign or_3285_nl = (~ (fsm_output[6])) | (fsm_output[5]) | (~ (fsm_output[2]))
      | mux_2469_nl;
  assign mux_2474_nl = MUX_s_1_2_2(mux_2473_nl, or_3285_nl, fsm_output[7]);
  assign nand_111_nl = ~((fsm_output[3]) & (~ mux_tmp_2466));
  assign mux_2467_nl = MUX_s_1_2_2(or_2824_cse, nand_111_nl, fsm_output[0]);
  assign or_2417_nl = (fsm_output[6]) | (~ (fsm_output[5])) | (fsm_output[2]) | mux_2467_nl;
  assign mux_2464_nl = MUX_s_1_2_2(or_2819_cse, mux_2463_cse, fsm_output[2]);
  assign or_2412_nl = (fsm_output[5]) | mux_2464_nl;
  assign nor_756_nl = ~((~ (fsm_output[3])) | (fsm_output[1]) | (~ (fsm_output[9]))
      | (~ (fsm_output[4])) | (fsm_output[10]));
  assign nor_757_nl = ~((fsm_output[3]) | (fsm_output[1]) | (fsm_output[9]) | nand_398_cse);
  assign mux_2462_nl = MUX_s_1_2_2(nor_756_nl, nor_757_nl, fsm_output[0]);
  assign nand_110_nl = ~((fsm_output[5]) & (fsm_output[2]) & mux_2462_nl);
  assign mux_2465_nl = MUX_s_1_2_2(or_2412_nl, nand_110_nl, fsm_output[6]);
  assign mux_2468_nl = MUX_s_1_2_2(or_2417_nl, mux_2465_nl, fsm_output[7]);
  assign mux_2475_itm = MUX_s_1_2_2(mux_2474_nl, mux_2468_nl, fsm_output[8]);
  assign nor_743_nl = ~((fsm_output[2]) | (~ (fsm_output[7])) | (~ (fsm_output[3]))
      | (fsm_output[9]) | (fsm_output[8]) | (~ (fsm_output[4])) | (fsm_output[10]));
  assign nor_744_nl = ~((~ (fsm_output[2])) | (fsm_output[7]) | (~ (fsm_output[3]))
      | (~ (fsm_output[9])) | (fsm_output[8]) | (fsm_output[4]) | (fsm_output[10]));
  assign mux_2486_nl = MUX_s_1_2_2(nor_743_nl, nor_744_nl, fsm_output[5]);
  assign or_3233_nl = (~ (fsm_output[7])) | (fsm_output[3]) | (~ (fsm_output[9]))
      | (~ (fsm_output[8])) | (fsm_output[4]) | (fsm_output[10]);
  assign or_3232_nl = (fsm_output[7]) | (fsm_output[3]) | (fsm_output[9]) | not_tmp_34;
  assign mux_3706_nl = MUX_s_1_2_2(or_3233_nl, or_3232_nl, fsm_output[2]);
  assign nor_745_nl = ~((fsm_output[5]) | mux_3706_nl);
  assign mux_2487_nl = MUX_s_1_2_2(mux_2486_nl, nor_745_nl, fsm_output[6]);
  assign or_2441_nl = (~ (fsm_output[7])) | (~ (fsm_output[3])) | (fsm_output[9])
      | (fsm_output[8]) | (fsm_output[4]) | (~ (fsm_output[10]));
  assign or_2439_nl = (fsm_output[7]) | (~ (fsm_output[3])) | (~ (fsm_output[9]))
      | (fsm_output[8]) | nand_398_cse;
  assign mux_2483_nl = MUX_s_1_2_2(or_2441_nl, or_2439_nl, fsm_output[2]);
  assign nor_746_nl = ~((fsm_output[5]) | mux_2483_nl);
  assign nor_1285_nl = ~((fsm_output[7]) | (fsm_output[3]) | (~ (fsm_output[8]))
      | (fsm_output[4]) | (fsm_output[9]) | (fsm_output[10]));
  assign nor_1286_nl = ~((~ (fsm_output[7])) | (fsm_output[3]) | (fsm_output[8])
      | (~ (fsm_output[4])) | (~ (fsm_output[9])) | (fsm_output[10]));
  assign mux_89_nl = MUX_s_1_2_2(nor_1285_nl, nor_1286_nl, fsm_output[2]);
  assign and_558_nl = (fsm_output[5]) & mux_89_nl;
  assign mux_2484_nl = MUX_s_1_2_2(nor_746_nl, and_558_nl, fsm_output[6]);
  assign mux_2488_nl = MUX_s_1_2_2(mux_2487_nl, mux_2484_nl, fsm_output[1]);
  assign nor_750_nl = ~((~ (fsm_output[7])) | (~ (fsm_output[3])) | (fsm_output[9])
      | not_tmp_34);
  assign nor_1278_nl = ~((fsm_output[7]) | (fsm_output[3]) | (fsm_output[8]) | (fsm_output[4])
      | (fsm_output[9]) | (~ (fsm_output[10])));
  assign mux_2478_nl = MUX_s_1_2_2(nor_750_nl, nor_1278_nl, fsm_output[2]);
  assign mux_2479_nl = MUX_s_1_2_2(nor_1276_cse, mux_2478_nl, fsm_output[5]);
  assign mux_2480_nl = MUX_s_1_2_2(mux_2479_nl, nor_1279_cse, fsm_output[6]);
  assign nor_1280_nl = ~((fsm_output[7]) | (~ (fsm_output[3])) | (~ (fsm_output[8]))
      | (~ (fsm_output[4])) | (~ (fsm_output[9])) | (fsm_output[10]));
  assign nor_1281_nl = ~((~ (fsm_output[7])) | (fsm_output[3]) | (~ (fsm_output[8]))
      | (fsm_output[4]) | (fsm_output[9]) | (fsm_output[10]));
  assign mux_93_nl = MUX_s_1_2_2(nor_1280_nl, nor_1281_nl, fsm_output[2]);
  assign mux_94_nl = MUX_s_1_2_2(mux_93_nl, nor_544_cse, fsm_output[5]);
  assign and_796_nl = (fsm_output[6]) & mux_94_nl;
  assign mux_2481_nl = MUX_s_1_2_2(mux_2480_nl, and_796_nl, fsm_output[1]);
  assign not_tmp_519 = MUX_s_1_2_2(mux_2488_nl, mux_2481_nl, fsm_output[0]);
  assign and_dcpl_264 = ~((fsm_output[10]) | (fsm_output[6]));
  assign mux_2490_nl = MUX_s_1_2_2((~ (fsm_output[3])), (fsm_output[3]), fsm_output[1]);
  assign or_463_nl = (~ (fsm_output[1])) | (fsm_output[3]);
  assign mux_2491_nl = MUX_s_1_2_2(mux_2490_nl, or_463_nl, fsm_output[0]);
  assign mux_2492_nl = MUX_s_1_2_2(mux_2491_nl, (fsm_output[3]), fsm_output[2]);
  assign and_dcpl_266 = (~ mux_2492_nl) & and_dcpl_264 & (~ (fsm_output[7])) & (~
      (fsm_output[5])) & (~ (fsm_output[8])) & and_dcpl;
  assign and_dcpl_268 = ~((fsm_output[7:6]!=2'b00));
  assign nor_741_nl = ~((fsm_output[5]) | (~((fsm_output[0]) & (fsm_output[3]))));
  assign nor_742_nl = ~((~ (fsm_output[5])) | (fsm_output[0]) | (fsm_output[3]));
  assign mux_2496_nl = MUX_s_1_2_2(nor_741_nl, nor_742_nl, fsm_output[4]);
  assign and_dcpl_273 = mux_2496_nl & and_dcpl_26 & and_dcpl_268 & (~ (fsm_output[2]))
      & nor_610_cse;
  assign mux_tmp_2502 = MUX_s_1_2_2(and_dcpl_101, mux_tmp_2239, fsm_output[2]);
  assign not_tmp_529 = ~(and_459_cse | (fsm_output[10]));
  assign nor_tmp_330 = (and_573_cse | (fsm_output[3:2]!=2'b00)) & (fsm_output[10]);
  assign or_2468_nl = (or_2385_cse & (fsm_output[3])) | (fsm_output[10]);
  assign mux_tmp_2508 = MUX_s_1_2_2(nor_tmp_330, or_2468_nl, fsm_output[9]);
  assign or_tmp_2416 = and_458_cse | (fsm_output[10]);
  assign or_tmp_2419 = and_440_cse | (fsm_output[10]);
  assign mux_tmp_2519 = MUX_s_1_2_2(mux_tmp_2239, nor_tmp_6, fsm_output[2]);
  assign mux_tmp_2523 = MUX_s_1_2_2(and_dcpl_101, nor_tmp_6, fsm_output[2]);
  assign mux_tmp_2525 = MUX_s_1_2_2(mux_tmp_2502, mux_tmp_2519, fsm_output[1]);
  assign nor_tmp_338 = or_2894_cse & (fsm_output[10]);
  assign or_3280_cse = and_573_cse | (fsm_output[2]);
  assign or_tmp_2429 = (or_3280_cse & (fsm_output[3])) | (fsm_output[10]);
  assign or_3279_cse = (fsm_output[3:2]!=2'b00);
  assign nor_tmp_342 = or_3279_cse & (fsm_output[10]);
  assign or_2489_nl = (fsm_output[2]) | (fsm_output[3]) | (fsm_output[10]);
  assign mux_tmp_2549 = MUX_s_1_2_2(or_tmp_2429, or_2489_nl, fsm_output[9]);
  assign mux_tmp_2650 = MUX_s_1_2_2(nor_601_cse, and_816_cse, fsm_output[7]);
  assign and_dcpl_279 = and_dcpl_40 & and_dcpl_30;
  assign and_dcpl_281 = and_dcpl_103 & and_dcpl_116;
  assign mux_tmp_2687 = MUX_s_1_2_2((~ and_dcpl_240), nor_tmp_6, fsm_output[6]);
  assign or_tmp_2474 = (fsm_output[6]) | or_tmp_2275;
  assign mux_tmp_2696 = MUX_s_1_2_2(and_dcpl_101, or_tmp_21, fsm_output[6]);
  assign nand_117_nl = ~((fsm_output[6]) & (~ or_tmp_2248));
  assign mux_tmp_2698 = MUX_s_1_2_2((~ (fsm_output[6])), nand_117_nl, fsm_output[7]);
  assign nor_719_nl = ~((fsm_output[6]) | (~ or_tmp_2230));
  assign mux_tmp_2701 = MUX_s_1_2_2(nor_719_nl, or_tmp_4, fsm_output[7]);
  assign or_tmp_2479 = (fsm_output[6]) | and_dcpl_101;
  assign nand_tmp_119 = ~((fsm_output[6]) & (~ nor_tmp_300));
  assign or_tmp_2483 = (fsm_output[0]) | (fsm_output[1]) | (fsm_output[3]) | (~ (fsm_output[10]));
  assign and_dcpl_283 = and_dcpl_128 & and_dcpl_100 & and_dcpl_116;
  assign and_dcpl_305 = and_dcpl_2 & and_dcpl;
  assign or_2556_nl = (fsm_output[7]) | (fsm_output[9]) | (~ (fsm_output[8])) | (fsm_output[4])
      | (fsm_output[10]);
  assign or_2555_nl = (~ (fsm_output[7])) | (~ (fsm_output[9])) | (fsm_output[8])
      | (~ (fsm_output[4])) | (fsm_output[10]);
  assign mux_2746_cse = MUX_s_1_2_2(or_2556_nl, or_2555_nl, fsm_output[2]);
  assign nor_702_nl = ~((fsm_output[1]) | (fsm_output[2]) | (~ (fsm_output[7])) |
      (~ (fsm_output[9])) | (fsm_output[8]) | (~ (fsm_output[4])) | (fsm_output[10]));
  assign nor_704_nl = ~((fsm_output[2]) | (fsm_output[7]) | (fsm_output[9]) | (fsm_output[8])
      | (~ (fsm_output[4])) | (fsm_output[10]));
  assign mux_2753_nl = MUX_s_1_2_2(nor_539_cse, nor_704_nl, fsm_output[1]);
  assign mux_2754_nl = MUX_s_1_2_2(nor_702_nl, mux_2753_nl, fsm_output[5]);
  assign nor_705_nl = ~((fsm_output[5]) | (~ (fsm_output[1])) | (~ (fsm_output[2]))
      | (~ (fsm_output[7])) | (fsm_output[9]) | (~ (fsm_output[8])) | (fsm_output[4])
      | (fsm_output[10]));
  assign mux_2755_nl = MUX_s_1_2_2(mux_2754_nl, nor_705_nl, fsm_output[6]);
  assign nor_706_nl = ~((~ (fsm_output[5])) | (fsm_output[1]) | (fsm_output[2]) |
      (~ (fsm_output[7])) | (fsm_output[9]) | not_tmp_34);
  assign nor_707_nl = ~((~ (fsm_output[1])) | (fsm_output[2]) | (fsm_output[7]) |
      (~ (fsm_output[9])) | (~ (fsm_output[8])) | (~ (fsm_output[4])) | (fsm_output[10]));
  assign nor_708_nl = ~((~ (fsm_output[2])) | (~ (fsm_output[7])) | (fsm_output[9])
      | (fsm_output[8]) | (~ (fsm_output[4])) | (fsm_output[10]));
  assign nor_1296_nl = ~((~ (fsm_output[2])) | (~ (fsm_output[7])) | (fsm_output[9])
      | (fsm_output[8]) | (fsm_output[4]) | (~ (fsm_output[10])));
  assign mux_2750_nl = MUX_s_1_2_2(nor_708_nl, nor_1296_nl, fsm_output[1]);
  assign mux_2751_nl = MUX_s_1_2_2(nor_707_nl, mux_2750_nl, fsm_output[5]);
  assign mux_2752_nl = MUX_s_1_2_2(nor_706_nl, mux_2751_nl, fsm_output[6]);
  assign mux_2756_nl = MUX_s_1_2_2(mux_2755_nl, mux_2752_nl, fsm_output[3]);
  assign nor_710_nl = ~((fsm_output[5]) | (~ (fsm_output[1])) | (~ (fsm_output[2]))
      | (~ (fsm_output[7])) | (fsm_output[9]) | (fsm_output[8]) | (~ (fsm_output[4]))
      | (fsm_output[10]));
  assign nor_711_nl = ~((~ (fsm_output[1])) | (fsm_output[2]) | (fsm_output[7]) |
      (fsm_output[9]) | not_tmp_34);
  assign nor_712_nl = ~((fsm_output[1]) | mux_2746_cse);
  assign mux_2747_nl = MUX_s_1_2_2(nor_711_nl, nor_712_nl, fsm_output[5]);
  assign mux_2748_nl = MUX_s_1_2_2(nor_710_nl, mux_2747_nl, fsm_output[6]);
  assign or_53_nl = (~ (fsm_output[7])) | (fsm_output[9]) | (fsm_output[8]) | (fsm_output[4])
      | (~ (fsm_output[10]));
  assign or_51_nl = (fsm_output[9:7]!=3'b100) | nand_398_cse;
  assign mux_74_nl = MUX_s_1_2_2(or_53_nl, or_51_nl, fsm_output[2]);
  assign or_2553_nl = (fsm_output[1]) | mux_74_nl;
  assign nand_120_nl = ~((fsm_output[1]) & mux_71_cse);
  assign mux_2745_nl = MUX_s_1_2_2(or_2553_nl, nand_120_nl, fsm_output[5]);
  assign nor_713_nl = ~((fsm_output[6]) | mux_2745_nl);
  assign mux_2749_nl = MUX_s_1_2_2(mux_2748_nl, nor_713_nl, fsm_output[3]);
  assign not_tmp_596 = MUX_s_1_2_2(mux_2756_nl, mux_2749_nl, fsm_output[0]);
  assign or_tmp_2516 = (fsm_output[2]) | (~ (fsm_output[7])) | (fsm_output[4]) |
      (fsm_output[10]);
  assign or_2578_nl = (~ (fsm_output[2])) | (fsm_output[7]) | nand_398_cse;
  assign mux_tmp_2758 = MUX_s_1_2_2(or_2578_nl, or_tmp_2516, fsm_output[9]);
  assign mux_tmp_2788 = MUX_s_1_2_2(or_tmp_2238, (fsm_output[10]), fsm_output[6]);
  assign mux_tmp_2790 = MUX_s_1_2_2(or_tmp_21, or_tmp_237, fsm_output[6]);
  assign or_2621_nl = (fsm_output[0]) | (~ and_dcpl_240);
  assign mux_tmp_2796 = MUX_s_1_2_2(or_2621_nl, mux_tmp_2309, fsm_output[6]);
  assign mux_2799_nl = MUX_s_1_2_2(nor_tmp_6, mux_tmp_2239, fsm_output[1]);
  assign mux_tmp_2800 = MUX_s_1_2_2(and_dcpl_240, mux_2799_nl, fsm_output[0]);
  assign mux_tmp_2813 = MUX_s_1_2_2(or_tmp_2277, or_tmp_2230, fsm_output[6]);
  assign or_207_nl = (fsm_output[4]) | (~ (fsm_output[10]));
  assign mux_2871_nl = MUX_s_1_2_2(or_tmp_178, or_207_nl, fsm_output[1]);
  assign or_tmp_2594 = (fsm_output[3]) | (fsm_output[9]) | mux_2871_nl;
  assign nor_672_nl = ~((~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[1]) |
      nand_398_cse);
  assign nor_673_nl = ~((fsm_output[3]) | (~ (fsm_output[9])) | (fsm_output[1]) |
      nand_398_cse);
  assign mux_2878_nl = MUX_s_1_2_2(nor_672_nl, nor_673_nl, fsm_output[0]);
  assign mux_2879_nl = MUX_s_1_2_2(mux_2878_nl, and_464_cse, fsm_output[2]);
  assign and_503_nl = (~((fsm_output[6:5]!=2'b01))) & mux_2879_nl;
  assign or_2662_nl = (~ (fsm_output[2])) | (~ (fsm_output[0])) | (~ (fsm_output[3]))
      | (fsm_output[9]) | (fsm_output[1]) | nand_398_cse;
  assign or_2659_nl = (fsm_output[0]) | (fsm_output[3]) | (~ (fsm_output[9])) | (fsm_output[1])
      | (fsm_output[4]) | (fsm_output[10]);
  assign mux_2876_nl = MUX_s_1_2_2(or_2839_cse, or_2659_nl, fsm_output[2]);
  assign mux_2877_nl = MUX_s_1_2_2(or_2662_nl, mux_2876_nl, fsm_output[5]);
  assign nor_674_nl = ~((fsm_output[6]) | mux_2877_nl);
  assign mux_2880_nl = MUX_s_1_2_2(and_503_nl, nor_674_nl, fsm_output[7]);
  assign mux_2873_nl = MUX_s_1_2_2(or_tmp_2594, or_529_cse, fsm_output[0]);
  assign nor_675_nl = ~((fsm_output[5]) | (fsm_output[2]) | mux_2873_nl);
  assign mux_2872_nl = MUX_s_1_2_2(or_525_cse, or_tmp_2594, fsm_output[0]);
  assign and_505_nl = (fsm_output[5]) & (fsm_output[2]) & (~ mux_2872_nl);
  assign mux_2874_nl = MUX_s_1_2_2(nor_675_nl, and_505_nl, fsm_output[6]);
  assign or_2647_nl = (fsm_output[0]) | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[1])
      | (fsm_output[4]) | (~ (fsm_output[10]));
  assign mux_2870_nl = MUX_s_1_2_2(mux_2463_cse, or_2647_nl, fsm_output[2]);
  assign nor_676_nl = ~((fsm_output[6:5]!=2'b10) | mux_2870_nl);
  assign mux_2875_nl = MUX_s_1_2_2(mux_2874_nl, nor_676_nl, fsm_output[7]);
  assign not_tmp_634 = MUX_s_1_2_2(mux_2880_nl, mux_2875_nl, fsm_output[8]);
  assign or_tmp_2631 = (fsm_output[2]) | (~ (fsm_output[8])) | (~ (fsm_output[7]))
      | (fsm_output[4]) | (fsm_output[10]);
  assign nor_654_nl = ~((~ (fsm_output[9])) | (~ (fsm_output[2])) | (fsm_output[8])
      | (fsm_output[7]) | (fsm_output[4]) | (~ (fsm_output[10])));
  assign nor_655_nl = ~((~ (fsm_output[2])) | (fsm_output[8]) | (fsm_output[7]) |
      (fsm_output[4]) | (fsm_output[10]));
  assign nor_656_nl = ~((fsm_output[2]) | (fsm_output[8]) | (fsm_output[7]) | (~
      (fsm_output[4])) | (fsm_output[10]));
  assign mux_2899_nl = MUX_s_1_2_2(nor_655_nl, nor_656_nl, fsm_output[9]);
  assign mux_2900_nl = MUX_s_1_2_2(nor_654_nl, mux_2899_nl, fsm_output[1]);
  assign and_498_nl = (fsm_output[6]) & mux_2900_nl;
  assign nor_657_nl = ~((fsm_output[1]) | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[8])
      | nand_240_cse);
  assign and_499_nl = (fsm_output[1]) & (fsm_output[9]) & (fsm_output[2]) & (fsm_output[8])
      & (fsm_output[7]) & (~ (fsm_output[4])) & (~ (fsm_output[10]));
  assign mux_2898_nl = MUX_s_1_2_2(nor_657_nl, and_499_nl, fsm_output[6]);
  assign mux_2901_nl = MUX_s_1_2_2(and_498_nl, mux_2898_nl, fsm_output[5]);
  assign or_2699_nl = (~ (fsm_output[2])) | (~ (fsm_output[8])) | (fsm_output[7])
      | (~ (fsm_output[4])) | (fsm_output[10]);
  assign mux_2896_nl = MUX_s_1_2_2(or_tmp_2631, or_2699_nl, fsm_output[9]);
  assign nor_658_nl = ~((fsm_output[6]) | (fsm_output[1]) | mux_2896_nl);
  assign nor_659_nl = ~((~ (fsm_output[1])) | (fsm_output[9]) | (~ (fsm_output[2]))
      | (fsm_output[8]) | (~ (fsm_output[7])) | (~ (fsm_output[4])) | (fsm_output[10]));
  assign nor_660_nl = ~((~ (fsm_output[1])) | (fsm_output[9]) | (fsm_output[2]) |
      (~ (fsm_output[8])) | (fsm_output[7]) | nand_398_cse);
  assign mux_2895_nl = MUX_s_1_2_2(nor_659_nl, nor_660_nl, fsm_output[6]);
  assign mux_2897_nl = MUX_s_1_2_2(nor_658_nl, mux_2895_nl, fsm_output[5]);
  assign mux_2902_nl = MUX_s_1_2_2(mux_2901_nl, mux_2897_nl, fsm_output[3]);
  assign or_2693_nl = (~ (fsm_output[2])) | (~ (fsm_output[8])) | (fsm_output[7])
      | nand_398_cse;
  assign mux_2892_nl = MUX_s_1_2_2(or_2693_nl, or_tmp_2631, fsm_output[9]);
  assign nor_661_nl = ~((fsm_output[6]) | (fsm_output[1]) | mux_2892_nl);
  assign nor_662_nl = ~((fsm_output[2]) | (~ (fsm_output[8])) | (fsm_output[7]) |
      (fsm_output[4]) | (fsm_output[10]));
  assign nor_663_nl = ~((~ (fsm_output[2])) | (fsm_output[8]) | (~ (fsm_output[7]))
      | (~ (fsm_output[4])) | (fsm_output[10]));
  assign mux_2891_nl = MUX_s_1_2_2(nor_662_nl, nor_663_nl, fsm_output[9]);
  assign and_500_nl = (~((fsm_output[6]) | (~ (fsm_output[1])))) & mux_2891_nl;
  assign mux_2893_nl = MUX_s_1_2_2(nor_661_nl, and_500_nl, fsm_output[5]);
  assign nor_664_nl = ~((~ (fsm_output[6])) | (~ (fsm_output[1])) | (fsm_output[9])
      | mux_3498_cse);
  assign nor_665_nl = ~((~ (fsm_output[6])) | (fsm_output[1]) | (fsm_output[9]) |
      (~ (fsm_output[2])) | (~ (fsm_output[8])) | (~ (fsm_output[7])) | (fsm_output[4])
      | (fsm_output[10]));
  assign mux_2890_nl = MUX_s_1_2_2(nor_664_nl, nor_665_nl, fsm_output[5]);
  assign mux_2894_nl = MUX_s_1_2_2(mux_2893_nl, mux_2890_nl, fsm_output[3]);
  assign not_tmp_646 = MUX_s_1_2_2(mux_2902_nl, mux_2894_nl, fsm_output[0]);
  assign or_248_nl = (fsm_output[10:9]!=2'b10);
  assign mux_523_nl = MUX_s_1_2_2(or_248_nl, and_816_cse, fsm_output[4]);
  assign or_tmp_2649 = (fsm_output[8]) | mux_523_nl;
  assign nand_tmp_136 = (fsm_output[8]) | (~ (fsm_output[4])) | and_816_cse;
  assign mux_tmp_2905 = MUX_s_1_2_2(nand_tmp_136, or_tmp_2649, fsm_output[1]);
  assign nand_tmp_137 = ~((fsm_output[4]) & (~ mux_726_cse));
  assign mux_tmp_2907 = MUX_s_1_2_2(nand_tmp_137, or_tmp_182, fsm_output[8]);
  assign or_tmp_2652 = (~ (fsm_output[4])) | (fsm_output[9]) | (~ (fsm_output[10]));
  assign or_tmp_2653 = (fsm_output[4]) | and_816_cse;
  assign mux_tmp_2911 = MUX_s_1_2_2(and_816_cse, or_tmp_187, fsm_output[4]);
  assign mux_tmp_2912 = MUX_s_1_2_2(mux_tmp_2911, or_tmp_2652, fsm_output[8]);
  assign mux_2910_nl = MUX_s_1_2_2(or_tmp_2653, or_tmp_2652, fsm_output[8]);
  assign mux_tmp_2913 = MUX_s_1_2_2(mux_tmp_2912, mux_2910_nl, fsm_output[1]);
  assign mux_tmp_2919 = MUX_s_1_2_2(or_tmp_179, nand_tmp_137, fsm_output[8]);
  assign mux_2920_nl = MUX_s_1_2_2(or_tmp_187, (~ and_816_cse), fsm_output[4]);
  assign mux_tmp_2921 = MUX_s_1_2_2(mux_2920_nl, mux_tmp_2911, fsm_output[8]);
  assign mux_tmp_2930 = MUX_s_1_2_2(or_tmp_2652, or_tmp_179, fsm_output[8]);
  assign or_tmp_2659 = (fsm_output[8]) | mux_tmp_2911;
  assign or_tmp_2663 = (fsm_output[8]) | (~ or_tmp_2653);
  assign mux_520_nl = MUX_s_1_2_2(mux_726_cse, and_816_cse, fsm_output[4]);
  assign nand_tmp_140 = ~((fsm_output[8]) & (~ mux_520_nl));
  assign or_tmp_2707 = (fsm_output[7]) | (~((fsm_output[2]) & (fsm_output[4]) & (fsm_output[10])));
  assign and_dcpl_332 = and_dcpl_128 & and_dcpl_117 & and_dcpl_116;
  assign nor_627_nl = ~((fsm_output[9]) | (~ (fsm_output[4])) | (fsm_output[10]));
  assign nor_628_nl = ~((fsm_output[9]) | (fsm_output[4]) | (~ (fsm_output[10])));
  assign mux_3168_nl = MUX_s_1_2_2(nor_627_nl, nor_628_nl, fsm_output[1]);
  assign nand_tmp_148 = ~((fsm_output[3]) & mux_3168_nl);
  assign or_2886_nl = (or_2894_cse & (fsm_output[4])) | (fsm_output[8:6]!=3'b000);
  assign mux_3213_nl = MUX_s_1_2_2(or_2951_cse, or_2886_nl, fsm_output[5]);
  assign or_3260_nl = (fsm_output[10]) | mux_3213_nl;
  assign or_2882_nl = (or_2348_cse & (fsm_output[4])) | (fsm_output[8:6]!=3'b000);
  assign mux_3212_nl = MUX_s_1_2_2(or_2951_cse, or_2882_nl, and_459_cse);
  assign nand_220_nl = ~((fsm_output[10]) & ((fsm_output[5]) | mux_3212_nl));
  assign not_tmp_708 = MUX_s_1_2_2(or_3260_nl, nand_220_nl, fsm_output[9]);
  assign nor_tmp_445 = or_2935_cse & (fsm_output[9]);
  assign mux_tmp_3219 = MUX_s_1_2_2((~ (fsm_output[9])), (fsm_output[9]), or_2935_cse);
  assign or_2905_nl = (fsm_output[7]) | (fsm_output[6]) | (fsm_output[1]) | (fsm_output[3]);
  assign mux_3235_nl = MUX_s_1_2_2(or_2520_cse, or_2905_nl, fsm_output[5]);
  assign or_2904_nl = (fsm_output[7:5]!=3'b000);
  assign mux_tmp_3236 = MUX_s_1_2_2(mux_3235_nl, or_2904_nl, fsm_output[2]);
  assign or_tmp_2849 = nor_1316_cse | (fsm_output[9]);
  assign mux_tmp_3244 = MUX_s_1_2_2((~ (fsm_output[9])), (fsm_output[9]), or_2951_cse);
  assign nor_tmp_456 = (fsm_output[9:7]==3'b111);
  assign mux_tmp_3256 = MUX_s_1_2_2(nor_610_cse, nor_tmp_116, fsm_output[7]);
  assign not_tmp_728 = ~((fsm_output[9:7]!=3'b000));
  assign or_tmp_2864 = (~((fsm_output[9:6]!=4'b0000))) | (fsm_output[10]);
  assign mux_tmp_3269 = MUX_s_1_2_2(and_dcpl_264, (fsm_output[10]), fsm_output[7]);
  assign nor_tmp_461 = (and_450_cse | (fsm_output[9:8]!=2'b00)) & (fsm_output[10]);
  assign mux_3279_nl = MUX_s_1_2_2(mux_tmp_741, and_754_cse, fsm_output[7]);
  assign and_436_nl = ((fsm_output[9:7]!=3'b000)) & (fsm_output[10]);
  assign mux_tmp_3280 = MUX_s_1_2_2(mux_3279_nl, and_436_nl, fsm_output[6]);
  assign mux_tmp_3281 = MUX_s_1_2_2(mux_tmp_741, and_754_cse, or_2520_cse);
  assign nand_tmp_157 = ~((fsm_output[8]) & nand_376_cse);
  assign mux_tmp_3323 = MUX_s_1_2_2(or_tmp_179, mux_tmp_374, fsm_output[8]);
  assign mux_3350_nl = MUX_s_1_2_2(mux_tmp_381, mux_tmp_3323, fsm_output[1]);
  assign mux_3351_nl = MUX_s_1_2_2(mux_382_cse, mux_3350_nl, fsm_output[0]);
  assign mux_3352_nl = MUX_s_1_2_2(nand_tmp_12, mux_3351_nl, fsm_output[6]);
  assign mux_3353_nl = MUX_s_1_2_2(mux_3352_nl, mux_3557_cse, fsm_output[5]);
  assign mux_3354_nl = MUX_s_1_2_2(mux_3353_nl, mux_3555_cse, fsm_output[7]);
  assign mux_3368_nl = MUX_s_1_2_2(mux_3575_cse, mux_3354_nl, fsm_output[3]);
  assign mux_3369_itm = MUX_s_1_2_2(mux_3368_nl, mux_3551_cse, fsm_output[2]);
  assign mux_3380_nl = MUX_s_1_2_2(nor_1276_cse, mux_3603_cse, fsm_output[5]);
  assign mux_3381_nl = MUX_s_1_2_2(mux_3380_nl, nor_1279_cse, fsm_output[6]);
  assign nor_591_nl = ~((~ (fsm_output[2])) | (~ (fsm_output[7])) | (fsm_output[9])
      | (~ (fsm_output[8])) | (fsm_output[4]) | (fsm_output[10]));
  assign nor_1295_nl = ~((fsm_output[2]) | (fsm_output[7]) | (~ (fsm_output[9]))
      | (~ (fsm_output[8])) | (~ (fsm_output[4])) | (fsm_output[10]));
  assign mux_3377_nl = MUX_s_1_2_2(nor_591_nl, nor_1295_nl, fsm_output[3]);
  assign mux_3378_nl = MUX_s_1_2_2(mux_3377_nl, nor_544_cse, fsm_output[5]);
  assign and_417_nl = (fsm_output[6]) & mux_3378_nl;
  assign mux_3382_nl = MUX_s_1_2_2(mux_3381_nl, and_417_nl, fsm_output[1]);
  assign nor_594_nl = ~((~ (fsm_output[7])) | (fsm_output[9]) | (fsm_output[8]) |
      (fsm_output[4]) | (~ (fsm_output[10])));
  assign nor_595_nl = ~((fsm_output[9:7]!=3'b100) | nand_398_cse);
  assign mux_3374_nl = MUX_s_1_2_2(nor_594_nl, nor_595_nl, fsm_output[2]);
  assign and_418_nl = nor_515_cse & mux_3374_nl;
  assign nor_596_nl = ~((~ (fsm_output[5])) | (fsm_output[3]) | mux_2746_cse);
  assign mux_3375_nl = MUX_s_1_2_2(and_418_nl, nor_596_nl, fsm_output[6]);
  assign nor_1287_nl = ~((~ (fsm_output[2])) | (~ (fsm_output[7])) | (fsm_output[3])
      | (fsm_output[8]) | (~ (fsm_output[4])) | (fsm_output[9]) | (fsm_output[10]));
  assign and_419_nl = (fsm_output[3]) & mux_71_cse;
  assign mux_3371_nl = MUX_s_1_2_2(nor_1287_nl, and_419_nl, fsm_output[5]);
  assign mux_3372_nl = MUX_s_1_2_2(mux_3371_nl, nor_545_cse, fsm_output[6]);
  assign mux_3376_nl = MUX_s_1_2_2(mux_3375_nl, mux_3372_nl, fsm_output[1]);
  assign not_tmp_762 = MUX_s_1_2_2(mux_3382_nl, mux_3376_nl, fsm_output[0]);
  assign or_3007_nl = (fsm_output[1]) | (fsm_output[2]) | (~ (fsm_output[7])) | (~
      (fsm_output[8])) | (fsm_output[4]) | (fsm_output[10]);
  assign or_3006_nl = (~ (fsm_output[1])) | (~ (fsm_output[2])) | (~ (fsm_output[7]))
      | (fsm_output[8]) | (~ (fsm_output[4])) | (fsm_output[10]);
  assign mux_tmp_3386 = MUX_s_1_2_2(or_3007_nl, or_3006_nl, fsm_output[5]);
  assign mux_3406_nl = MUX_s_1_2_2(or_tmp_178, or_tmp_179, fsm_output[8]);
  assign or_3037_nl = (~ (fsm_output[1])) | (fsm_output[2]) | (fsm_output[7]) | mux_3406_nl;
  assign mux_3407_nl = MUX_s_1_2_2(or_3016_cse, or_3037_nl, fsm_output[5]);
  assign mux_3408_nl = MUX_s_1_2_2(or_3018_cse, mux_3407_nl, fsm_output[0]);
  assign nor_573_nl = ~((fsm_output[6]) | mux_3408_nl);
  assign mux_3409_nl = MUX_s_1_2_2(nor_573_nl, mux_3392_cse, fsm_output[3]);
  assign not_tmp_776 = MUX_s_1_2_2(mux_3409_nl, mux_3388_cse, fsm_output[9]);
  assign mux_tmp_3418 = MUX_s_1_2_2(or_tmp_118, or_154_cse, fsm_output[5]);
  assign mux_3421_nl = MUX_s_1_2_2(or_tmp_179, or_tmp_178, fsm_output[8]);
  assign mux_tmp_3422 = MUX_s_1_2_2(mux_3421_nl, or_tmp_118, fsm_output[5]);
  assign mux_tmp_3426 = MUX_s_1_2_2((~ and_491_cse), or_tmp_179, fsm_output[8]);
  assign mux_tmp_3430 = MUX_s_1_2_2(or_tmp_118, or_tmp_191, fsm_output[5]);
  assign mux_tmp_3436 = MUX_s_1_2_2(or_154_cse, or_tmp_110, fsm_output[5]);
  assign nand_tmp_167 = ~((fsm_output[8]) & (~ and_491_cse));
  assign mux_tmp_3449 = MUX_s_1_2_2(nand_tmp_167, or_tmp_191, fsm_output[5]);
  assign mux_tmp_3450 = MUX_s_1_2_2((~ (fsm_output[8])), or_tmp_150, fsm_output[5]);
  assign mux_tmp_3452 = MUX_s_1_2_2((~ (fsm_output[8])), mux_tmp_3426, fsm_output[5]);
  assign mux_tmp_3456 = MUX_s_1_2_2((~ (fsm_output[4])), and_491_cse, fsm_output[8]);
  assign mux_tmp_3458 = MUX_s_1_2_2((~ and_491_cse), and_491_cse, fsm_output[8]);
  assign mux_tmp_3459 = MUX_s_1_2_2((~ or_tmp_191), mux_tmp_3458, fsm_output[5]);
  assign mux_tmp_3467 = MUX_s_1_2_2(not_tmp_34, nand_tmp_167, fsm_output[5]);
  assign nor_568_nl = ~((fsm_output[4]) | (~ (fsm_output[10])));
  assign mux_tmp_3468 = MUX_s_1_2_2(nor_568_nl, and_491_cse, fsm_output[8]);
  assign mux_tmp_3471 = MUX_s_1_2_2(mux_tmp_3468, (fsm_output[8]), fsm_output[5]);
  assign and_tmp_36 = (fsm_output[8]) & or_tmp_179;
  assign or_tmp_3025 = (fsm_output[6]) | (fsm_output[5]) | (~ (fsm_output[3])) |
      (fsm_output[8]) | (~ (fsm_output[10]));
  assign mux_3613_nl = MUX_s_1_2_2(and_dcpl_109, (fsm_output[10]), fsm_output[1]);
  assign or_tmp_3107 = (fsm_output[6]) | (~ mux_3613_nl);
  assign STAGE_LOOP_i_3_0_sva_mx0c1 = and_dcpl_111 & and_dcpl_106;
  assign and_540_cse = or_2348_cse & (fsm_output[2]);
  assign nor_738_cse = ~((fsm_output[3:1]!=3'b000));
  assign VEC_LOOP_j_sva_11_0_mx0c1 = and_dcpl_110 & and_dcpl_127 & and_dcpl_106;
  assign nor_724_nl = ~((fsm_output[2]) | (fsm_output[1]) | (fsm_output[9]) | (fsm_output[10]));
  assign mux_2662_nl = MUX_s_1_2_2(nor_601_cse, nor_724_nl, fsm_output[3]);
  assign and_521_nl = (fsm_output[0]) & (fsm_output[1]) & (fsm_output[9]) & (fsm_output[10]);
  assign mux_2661_nl = MUX_s_1_2_2(and_521_nl, and_816_cse, or_3279_cse);
  assign mux_2663_nl = MUX_s_1_2_2(mux_2662_nl, mux_2661_nl, fsm_output[7]);
  assign or_2522_nl = (fsm_output[6:4]!=3'b000);
  assign mux_2664_nl = MUX_s_1_2_2(mux_2663_nl, and_815_cse, or_2522_nl);
  assign modExp_result_sva_mx0c0 = MUX_s_1_2_2(mux_2664_nl, and_816_cse, fsm_output[8]);
  assign nl_STAGE_LOOP_acc_nl = (STAGE_LOOP_i_3_0_sva_2[3:1]) + 3'b011;
  assign STAGE_LOOP_acc_nl = nl_STAGE_LOOP_acc_nl[2:0];
  assign STAGE_LOOP_acc_itm_2_1 = readslicef_3_1_2(STAGE_LOOP_acc_nl);
  assign and_305_m1c = and_dcpl_128 & and_dcpl_108 & and_dcpl_279;
  assign and_307_m1c = and_dcpl_156 & and_dcpl_162 & and_dcpl_139;
  assign and_309_m1c = and_dcpl_102 & and_dcpl_173 & and_dcpl_245;
  assign and_312_m1c = and_dcpl_128 & and_dcpl_162 & and_dcpl_22 & and_dcpl;
  assign and_315_m1c = and_dcpl_124 & and_dcpl_117 & and_dcpl_46 & and_dcpl_50;
  assign and_317_m1c = and_dcpl_102 & and_dcpl_127 & and_dcpl_172;
  assign and_320_m1c = and_dcpl_102 & and_dcpl_204 & and_dcpl_2 & and_472_cse;
  assign and_322_m1c = and_dcpl_125 & and_dcpl_154 & and_472_cse;
  assign and_324_m1c = and_dcpl_140 & and_dcpl_145 & and_472_cse;
  assign and_327_m1c = and_dcpl_223 & and_dcpl_100 & and_dcpl_305;
  assign and_329_m1c = and_dcpl_215 & and_dcpl_108 & and_dcpl_98;
  assign and_331_m1c = and_dcpl_240 & and_dcpl_162 & and_dcpl_305;
  assign and_334_m1c = and_dcpl_110 & and_dcpl_173 & and_dcpl_154 & and_dcpl_30;
  assign and_336_m1c = and_dcpl_215 & and_dcpl_127 & and_dcpl_239;
  assign and_339_m1c = and_dcpl_215 & and_dcpl_117 & and_dcpl_40 & and_472_cse;
  assign and_139_nl = and_dcpl_129 & and_dcpl_98;
  assign or_533_nl = (fsm_output[2]) | (~((fsm_output[0]) & (fsm_output[1]) & (fsm_output[9])
      & (fsm_output[3]) & (fsm_output[4]) & (fsm_output[10])));
  assign or_531_nl = (~ (fsm_output[1])) | (fsm_output[9]) | (fsm_output[3]) | (fsm_output[4])
      | (~ (fsm_output[10]));
  assign mux_1041_nl = MUX_s_1_2_2(or_531_nl, or_529_cse, fsm_output[0]);
  assign or_532_nl = (fsm_output[2]) | mux_1041_nl;
  assign mux_1042_nl = MUX_s_1_2_2(or_533_nl, or_532_nl, fsm_output[5]);
  assign nor_1194_nl = ~((fsm_output[6]) | mux_1042_nl);
  assign or_527_nl = (fsm_output[0]) | (fsm_output[1]) | (~ (fsm_output[9])) | (fsm_output[3])
      | (fsm_output[4]) | (~ (fsm_output[10]));
  assign or_524_nl = (fsm_output[9]) | (fsm_output[3]) | (~ (fsm_output[4])) | (fsm_output[10]);
  assign or_523_nl = (fsm_output[9]) | (fsm_output[3]) | (fsm_output[4]) | (~ (fsm_output[10]));
  assign mux_1037_nl = MUX_s_1_2_2(or_524_nl, or_523_nl, fsm_output[1]);
  assign mux_1038_nl = MUX_s_1_2_2(or_525_cse, mux_1037_nl, fsm_output[0]);
  assign mux_1039_nl = MUX_s_1_2_2(or_527_nl, mux_1038_nl, fsm_output[2]);
  assign nor_1195_nl = ~((fsm_output[5]) | mux_1039_nl);
  assign nor_1196_nl = ~((~ (fsm_output[1])) | (fsm_output[9]) | (~ (fsm_output[3]))
      | (~ (fsm_output[4])) | (fsm_output[10]));
  assign nor_1197_nl = ~((~ (fsm_output[1])) | (~ (fsm_output[9])) | (fsm_output[3])
      | (~ (fsm_output[4])) | (fsm_output[10]));
  assign mux_1035_nl = MUX_s_1_2_2(nor_1196_nl, nor_1197_nl, fsm_output[0]);
  assign nor_1198_nl = ~((fsm_output[0]) | (fsm_output[1]) | (fsm_output[9]) | (~
      (fsm_output[3])) | (fsm_output[4]) | (~ (fsm_output[10])));
  assign mux_1036_nl = MUX_s_1_2_2(mux_1035_nl, nor_1198_nl, fsm_output[2]);
  assign and_660_nl = (fsm_output[5]) & mux_1036_nl;
  assign mux_1040_nl = MUX_s_1_2_2(nor_1195_nl, and_660_nl, fsm_output[6]);
  assign mux_1043_nl = MUX_s_1_2_2(nor_1194_nl, mux_1040_nl, fsm_output[7]);
  assign or_516_nl = (fsm_output[1]) | (fsm_output[9]) | (fsm_output[3]) | nand_398_cse;
  assign mux_1032_nl = MUX_s_1_2_2(or_tmp_453, or_516_nl, fsm_output[0]);
  assign or_514_nl = (~ (fsm_output[0])) | (~ (fsm_output[1])) | (fsm_output[9])
      | (~ (fsm_output[3])) | (~ (fsm_output[4])) | (fsm_output[10]);
  assign mux_1033_nl = MUX_s_1_2_2(mux_1032_nl, or_514_nl, fsm_output[2]);
  assign nor_1199_nl = ~((fsm_output[6:5]!=2'b10) | mux_1033_nl);
  assign or_512_nl = (~ (fsm_output[1])) | (fsm_output[9]) | (fsm_output[3]) | nand_398_cse;
  assign mux_1030_nl = MUX_s_1_2_2(or_512_nl, or_tmp_453, fsm_output[0]);
  assign and_661_nl = (fsm_output[5]) & (fsm_output[2]) & (~ mux_1030_nl);
  assign nor_1200_nl = ~((fsm_output[5]) | (~ (fsm_output[2])) | (fsm_output[0])
      | (fsm_output[1]) | (fsm_output[9]) | (fsm_output[3]) | (fsm_output[4]) | (fsm_output[10]));
  assign mux_1031_nl = MUX_s_1_2_2(and_661_nl, nor_1200_nl, fsm_output[6]);
  assign mux_1034_nl = MUX_s_1_2_2(nor_1199_nl, mux_1031_nl, fsm_output[7]);
  assign mux_1044_nl = MUX_s_1_2_2(mux_1043_nl, mux_1034_nl, fsm_output[8]);
  assign and_145_nl = not_tmp_240 & and_dcpl_101 & (fsm_output[1]) & (fsm_output[7])
      & (fsm_output[2]) & nor_610_cse;
  assign nor_1191_nl = ~((~ (fsm_output[8])) | (~ (fsm_output[2])) | (fsm_output[5])
      | (fsm_output[7]) | (fsm_output[0]) | (fsm_output[1]));
  assign nor_1192_nl = ~((fsm_output[8]) | (fsm_output[2]) | (~((fsm_output[5]) &
      (fsm_output[7]) & (fsm_output[0]) & (fsm_output[1]))));
  assign mux_1046_nl = MUX_s_1_2_2(nor_1191_nl, nor_1192_nl, fsm_output[4]);
  assign and_153_nl = mux_1046_nl & and_dcpl_123 & (fsm_output[6]) & (~ (fsm_output[9]));
  assign nor_1189_nl = ~((fsm_output[7]) | (~ (fsm_output[6])) | (fsm_output[0]));
  assign nor_1190_nl = ~((~ (fsm_output[7])) | (fsm_output[6]) | (~ (fsm_output[0])));
  assign mux_1047_nl = MUX_s_1_2_2(nor_1189_nl, nor_1190_nl, fsm_output[4]);
  assign and_162_nl = mux_1047_nl & and_dcpl_101 & (~ (fsm_output[1])) & (fsm_output[5])
      & (~ (fsm_output[2])) & and_dcpl_148;
  assign nor_1187_nl = ~((fsm_output[4]) | (~ (fsm_output[8])) | (~ (fsm_output[7]))
      | (~ (fsm_output[6])) | (~ (fsm_output[0])) | (fsm_output[1]));
  assign nor_1188_nl = ~((~ (fsm_output[4])) | (fsm_output[8]) | (fsm_output[7])
      | (fsm_output[6]) | (fsm_output[0]) | (~ (fsm_output[1])));
  assign mux_1048_nl = MUX_s_1_2_2(nor_1187_nl, nor_1188_nl, fsm_output[9]);
  assign and_170_nl = mux_1048_nl & and_dcpl_101 & and_dcpl_21;
  assign and_179_nl = mux_tmp_1049 & and_dcpl_124 & (~ (fsm_output[7])) & (fsm_output[5])
      & (~ (fsm_output[2])) & and_dcpl_165;
  assign nor_1185_nl = ~((~ (fsm_output[5])) | (~ (fsm_output[6])) | (fsm_output[0])
      | (fsm_output[1]) | (fsm_output[3]));
  assign nor_1186_nl = ~((fsm_output[5]) | (fsm_output[6]) | (~((fsm_output[0]) &
      (fsm_output[1]) & (fsm_output[3]))));
  assign mux_1050_nl = MUX_s_1_2_2(nor_1185_nl, nor_1186_nl, fsm_output[2]);
  assign and_188_nl = mux_1050_nl & (~ (fsm_output[10])) & (fsm_output[7]) & (~ (fsm_output[8]))
      & and_dcpl_50;
  assign nor_1183_nl = ~((~ (fsm_output[8])) | (fsm_output[5]) | (fsm_output[7])
      | (~ (fsm_output[0])));
  assign nor_1184_nl = ~((fsm_output[8]) | (~ (fsm_output[5])) | (~ (fsm_output[7]))
      | (fsm_output[0]));
  assign mux_1051_nl = MUX_s_1_2_2(nor_1183_nl, nor_1184_nl, fsm_output[4]);
  assign and_197_nl = mux_1051_nl & (~ (fsm_output[10])) & (~ (fsm_output[3])) &
      (~ (fsm_output[1])) & (fsm_output[6]) & (fsm_output[2]) & (fsm_output[9]);
  assign nor_1181_nl = ~((~ (fsm_output[5])) | (~ (fsm_output[7])) | (fsm_output[6])
      | (fsm_output[0]) | (~ (fsm_output[1])));
  assign nor_1182_nl = ~((fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[6]))
      | (~ (fsm_output[0])) | (fsm_output[1]));
  assign mux_1052_nl = MUX_s_1_2_2(nor_1181_nl, nor_1182_nl, fsm_output[4]);
  assign and_205_nl = mux_1052_nl & and_dcpl_123 & (~ (fsm_output[2])) & (fsm_output[8])
      & (fsm_output[9]);
  assign nor_1179_nl = ~((fsm_output[4]) | (fsm_output[8]) | (fsm_output[5]) | (fsm_output[7])
      | (~((fsm_output[0]) & (fsm_output[10]))));
  assign nor_1180_nl = ~((~ (fsm_output[4])) | (~ (fsm_output[8])) | (~ (fsm_output[5]))
      | (~ (fsm_output[7])) | (fsm_output[0]) | (fsm_output[10]));
  assign mux_1053_nl = MUX_s_1_2_2(nor_1179_nl, nor_1180_nl, fsm_output[9]);
  assign and_211_nl = mux_1053_nl & (fsm_output[3]) & (fsm_output[1]) & (~ (fsm_output[6]))
      & (fsm_output[2]);
  assign nor_1177_nl = ~((fsm_output[2]) | (fsm_output[6]) | nand_237_cse);
  assign nor_1178_nl = ~((~ (fsm_output[2])) | (~ (fsm_output[6])) | (fsm_output[0])
      | (fsm_output[1]));
  assign mux_1054_nl = MUX_s_1_2_2(nor_1177_nl, nor_1178_nl, fsm_output[4]);
  assign and_220_nl = mux_1054_nl & (fsm_output[10]) & (~ (fsm_output[3])) & (~ (fsm_output[7]))
      & (fsm_output[5]) & nor_610_cse;
  assign and_231_nl = mux_tmp_1049 & and_dcpl_215 & (fsm_output[7]) & (~ (fsm_output[5]))
      & (~ (fsm_output[2])) & nor_610_cse;
  assign nor_1175_nl = ~((fsm_output[8]) | (~ (fsm_output[7])) | (~ (fsm_output[6]))
      | (~ (fsm_output[0])) | (fsm_output[1]));
  assign nor_1176_nl = ~((~ (fsm_output[8])) | (fsm_output[7]) | (fsm_output[6])
      | (fsm_output[0]) | (~ (fsm_output[1])));
  assign mux_1055_nl = MUX_s_1_2_2(nor_1175_nl, nor_1176_nl, fsm_output[4]);
  assign and_238_nl = mux_1055_nl & nor_tmp_6 & (fsm_output[5]) & (fsm_output[2])
      & (~ (fsm_output[9]));
  assign and_817_nl = (fsm_output[5]) & (fsm_output[7]) & (~ (fsm_output[6])) & (fsm_output[0]);
  assign nor_1174_nl = ~((fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[6]))
      | (fsm_output[0]));
  assign mux_1056_nl = MUX_s_1_2_2(and_817_nl, nor_1174_nl, fsm_output[4]);
  assign and_246_nl = mux_1056_nl & (fsm_output[10]) & (~ (fsm_output[3])) & (fsm_output[1])
      & (~ (fsm_output[2])) & and_dcpl_148;
  assign and_657_nl = (fsm_output[4]) & (fsm_output[8]) & (fsm_output[2]) & (fsm_output[5])
      & (fsm_output[7]) & (fsm_output[0]) & (fsm_output[1]) & (~ (fsm_output[3]));
  assign nor_1172_nl = ~((fsm_output[4]) | (fsm_output[8]) | (fsm_output[2]) | (fsm_output[5])
      | (fsm_output[7]) | (fsm_output[0]) | (fsm_output[1]) | (~ (fsm_output[3])));
  assign mux_1057_nl = MUX_s_1_2_2(and_657_nl, nor_1172_nl, fsm_output[9]);
  assign and_253_nl = mux_1057_nl & and_dcpl_243;
  assign and_261_nl = not_tmp_240 & nor_tmp_6 & (~ (fsm_output[1])) & (~ (fsm_output[7]))
      & (fsm_output[2]) & and_dcpl_165;
  assign vec_rsc_0_0_i_adra_d_pff = MUX1HOT_v_8_19_2(COMP_LOOP_acc_psp_sva_1, (z_out_7[12:5]),
      COMP_LOOP_acc_psp_sva, (COMP_LOOP_acc_10_cse_12_1_1_sva[11:4]), (COMP_LOOP_acc_1_cse_2_sva[11:4]),
      (COMP_LOOP_acc_11_psp_sva[10:3]), (COMP_LOOP_acc_1_cse_4_sva[11:4]), (COMP_LOOP_acc_13_psp_sva[9:2]),
      (COMP_LOOP_acc_1_cse_6_sva[11:4]), (COMP_LOOP_acc_14_psp_sva[10:3]), (COMP_LOOP_acc_1_cse_8_sva[11:4]),
      (COMP_LOOP_acc_16_psp_sva[8:1]), (COMP_LOOP_acc_1_cse_10_sva[11:4]), (COMP_LOOP_acc_17_psp_sva[10:3]),
      (COMP_LOOP_acc_1_cse_12_sva[11:4]), (COMP_LOOP_acc_19_psp_sva[9:2]), (COMP_LOOP_acc_1_cse_14_sva[11:4]),
      (COMP_LOOP_acc_20_psp_sva[10:3]), (COMP_LOOP_acc_1_cse_sva[11:4]), {and_dcpl_119
      , COMP_LOOP_or_32_cse , and_139_nl , mux_1044_nl , and_145_nl , and_153_nl
      , and_162_nl , and_170_nl , and_179_nl , and_188_nl , and_197_nl , and_205_nl
      , and_211_nl , and_220_nl , and_231_nl , and_238_nl , and_246_nl , and_253_nl
      , and_261_nl});
  assign vec_rsc_0_0_i_da_d_pff = modulo_result_mux_1_cse;
  assign or_624_nl = (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b000) | (fsm_output[0]) |
      (VEC_LOOP_j_sva_11_0[0]) | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[9]))
      | (fsm_output[8]) | (~ (fsm_output[10]));
  assign mux_1093_nl = MUX_s_1_2_2(or_624_nl, or_622_cse, fsm_output[5]);
  assign mux_1094_nl = MUX_s_1_2_2(mux_1093_nl, or_621_cse, fsm_output[4]);
  assign or_615_nl = (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b000) | (fsm_output[0]) |
      (VEC_LOOP_j_sva_11_0[0]) | (fsm_output[3]) | (~ (fsm_output[6])) | (~ (fsm_output[9]))
      | (fsm_output[8]) | (fsm_output[10]);
  assign mux_1090_nl = MUX_s_1_2_2(or_617_cse, or_615_nl, fsm_output[5]);
  assign mux_1091_nl = MUX_s_1_2_2(mux_1090_nl, mux_tmp_1068, fsm_output[4]);
  assign mux_1095_nl = MUX_s_1_2_2(mux_1094_nl, mux_1091_nl, fsm_output[7]);
  assign mux_1089_nl = MUX_s_1_2_2(mux_tmp_1067, mux_1088_cse, fsm_output[7]);
  assign mux_1096_nl = MUX_s_1_2_2(mux_1095_nl, mux_1089_nl, fsm_output[2]);
  assign or_605_nl = (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0000) | (~ (fsm_output[0]))
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (~ (fsm_output[9])) | (fsm_output[8])
      | (fsm_output[10]);
  assign mux_1082_nl = MUX_s_1_2_2(or_607_cse, or_605_nl, fsm_output[5]);
  assign mux_1083_nl = MUX_s_1_2_2(or_609_cse, mux_1082_nl, fsm_output[4]);
  assign mux_1081_nl = MUX_s_1_2_2(mux_tmp_1062, nand_25_cse, fsm_output[4]);
  assign mux_1084_nl = MUX_s_1_2_2(mux_1083_nl, mux_1081_nl, fsm_output[7]);
  assign or_602_nl = (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b00) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b00)
      | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[9])) | (fsm_output[8])
      | (fsm_output[10]);
  assign mux_1076_nl = MUX_s_1_2_2(or_602_nl, or_601_cse, fsm_output[0]);
  assign mux_1077_nl = MUX_s_1_2_2(mux_1076_nl, or_tmp_515, fsm_output[5]);
  assign mux_1078_nl = MUX_s_1_2_2(or_tmp_518, mux_1077_nl, fsm_output[4]);
  assign or_597_nl = (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0000) | (~ (fsm_output[0]))
      | (fsm_output[3]) | (~ (fsm_output[6])) | (fsm_output[9]) | (fsm_output[8])
      | (fsm_output[10]);
  assign mux_1074_nl = MUX_s_1_2_2(mux_1073_cse, or_597_nl, fsm_output[5]);
  assign mux_1075_nl = MUX_s_1_2_2(mux_1074_nl, or_596_cse, fsm_output[4]);
  assign mux_1079_nl = MUX_s_1_2_2(mux_1078_nl, mux_1075_nl, fsm_output[7]);
  assign mux_1085_nl = MUX_s_1_2_2(mux_1084_nl, mux_1079_nl, fsm_output[2]);
  assign mux_1097_nl = MUX_s_1_2_2(mux_1096_nl, mux_1085_nl, fsm_output[1]);
  assign or_594_nl = (fsm_output[5:4]!=2'b00) | (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b000)
      | (fsm_output[0]) | (VEC_LOOP_j_sva_11_0[0]) | (~ (fsm_output[3])) | (fsm_output[6])
      | (~ (fsm_output[9])) | (fsm_output[8]) | (~ (fsm_output[10]));
  assign or_592_nl = (~ (fsm_output[5])) | (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b000)
      | (fsm_output[0]) | (VEC_LOOP_j_sva_11_0[0]) | (fsm_output[3]) | (~ (fsm_output[6]))
      | (~ (fsm_output[9])) | (fsm_output[8]) | (fsm_output[10]);
  assign mux_1069_nl = MUX_s_1_2_2(or_592_nl, mux_tmp_1068, fsm_output[4]);
  assign mux_1070_nl = MUX_s_1_2_2(or_594_nl, mux_1069_nl, fsm_output[7]);
  assign or_588_nl = (fsm_output[7]) | mux_tmp_1067;
  assign mux_1071_nl = MUX_s_1_2_2(mux_1070_nl, or_588_nl, fsm_output[2]);
  assign or_581_nl = (fsm_output[5:4]!=2'b11) | (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0000)
      | (~ (fsm_output[0])) | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (~ (fsm_output[9]))
      | (fsm_output[8]) | (fsm_output[10]);
  assign or_580_nl = (fsm_output[4]) | mux_tmp_1062;
  assign mux_1063_nl = MUX_s_1_2_2(or_581_nl, or_580_nl, fsm_output[7]);
  assign or_573_nl = (fsm_output[0]) | (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b00) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b00)
      | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[9])) | (fsm_output[8])
      | (fsm_output[10]);
  assign mux_1058_nl = MUX_s_1_2_2(or_573_nl, or_tmp_515, fsm_output[5]);
  assign mux_1059_nl = MUX_s_1_2_2(or_tmp_518, mux_1058_nl, fsm_output[4]);
  assign or_570_nl = (fsm_output[5:4]!=2'b10) | (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0000)
      | (~ (fsm_output[0])) | (fsm_output[3]) | (~ (fsm_output[6])) | (fsm_output[9])
      | (fsm_output[8]) | (fsm_output[10]);
  assign mux_1060_nl = MUX_s_1_2_2(mux_1059_nl, or_570_nl, fsm_output[7]);
  assign mux_1064_nl = MUX_s_1_2_2(mux_1063_nl, mux_1060_nl, fsm_output[2]);
  assign mux_1072_nl = MUX_s_1_2_2(mux_1071_nl, mux_1064_nl, fsm_output[1]);
  assign or_569_nl = (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0000);
  assign mux_1098_nl = MUX_s_1_2_2(mux_1097_nl, mux_1072_nl, or_569_nl);
  assign vec_rsc_0_0_i_wea_d_pff = ~ mux_1098_nl;
  assign nor_1148_cse = ~((z_out_7[4:1]!=4'b0000) | (fsm_output[3]) | (~ (fsm_output[9]))
      | (~ (fsm_output[1])) | (fsm_output[10]));
  assign or_642_cse = (z_out_7[4:1]!=4'b0000) | (~ (fsm_output[3])) | (~ (fsm_output[9]))
      | (fsm_output[1]) | (fsm_output[10]);
  assign nor_1147_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b0000) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[0]) | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[1])
      | (~ (fsm_output[10])));
  assign nor_1149_nl = ~((~ (fsm_output[3])) | (z_out_7[4:1]!=4'b0000) | (fsm_output[9])
      | (fsm_output[1]) | (fsm_output[10]));
  assign mux_1125_nl = MUX_s_1_2_2(nor_1148_cse, nor_1149_nl, fsm_output[0]);
  assign mux_1126_nl = MUX_s_1_2_2(nor_1147_nl, mux_1125_nl, fsm_output[8]);
  assign and_654_nl = nor_223_cse & mux_1126_nl;
  assign or_670_nl = (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0000) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (~ (fsm_output[1])) | (fsm_output[10]);
  assign or_669_nl = (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b000) | (VEC_LOOP_j_sva_11_0[0])
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[3]) | (fsm_output[9])
      | not_tmp_260;
  assign mux_1123_nl = MUX_s_1_2_2(or_670_nl, or_669_nl, fsm_output[0]);
  assign nor_1150_nl = ~((fsm_output[8:7]!=2'b00) | mux_1123_nl);
  assign nor_1151_nl = ~((~ (fsm_output[8])) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b0000) | (fsm_output[0]) | (fsm_output[3])
      | (fsm_output[9]) | (fsm_output[1]) | (fsm_output[10]));
  assign nor_1152_nl = ~((~ (fsm_output[8])) | (fsm_output[0]) | (z_out_7[4:1]!=4'b0000)
      | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[1]) | (~ (fsm_output[10])));
  assign mux_1122_nl = MUX_s_1_2_2(nor_1151_nl, nor_1152_nl, fsm_output[7]);
  assign mux_1124_nl = MUX_s_1_2_2(nor_1150_nl, mux_1122_nl, fsm_output[6]);
  assign mux_1127_nl = MUX_s_1_2_2(and_654_nl, mux_1124_nl, fsm_output[5]);
  assign nor_1153_nl = ~((~ (fsm_output[7])) | (fsm_output[8]) | (~ (fsm_output[0]))
      | (VEC_LOOP_j_sva_11_0[0]) | (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b000) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (~ (fsm_output[1])) | (fsm_output[10]));
  assign or_661_nl = (z_out_7[4:1]!=4'b0000) | (~ (fsm_output[3])) | (fsm_output[9])
      | (fsm_output[1]) | (~ (fsm_output[10]));
  assign or_659_nl = (fsm_output[3]) | (z_out_7[4:1]!=4'b0000) | (~ (fsm_output[9]))
      | (fsm_output[1]) | (~ (fsm_output[10]));
  assign mux_1118_nl = MUX_s_1_2_2(or_661_nl, or_659_nl, fsm_output[0]);
  assign nor_1154_nl = ~((fsm_output[8]) | mux_1118_nl);
  assign nor_1155_nl = ~((COMP_LOOP_acc_13_psp_sva[1:0]!=2'b00) | (~ (fsm_output[8]))
      | (~ (fsm_output[0])) | (VEC_LOOP_j_sva_11_0[0]) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (VEC_LOOP_j_sva_11_0[1]) | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[1])
      | (fsm_output[10]));
  assign mux_1119_nl = MUX_s_1_2_2(nor_1154_nl, nor_1155_nl, fsm_output[7]);
  assign mux_1120_nl = MUX_s_1_2_2(nor_1153_nl, mux_1119_nl, fsm_output[6]);
  assign nor_1156_nl = ~((fsm_output[8:7]!=2'b10) | (z_out_7[4:1]!=4'b0000) | (fsm_output[0])
      | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[1]) | (fsm_output[10]));
  assign nor_1157_nl = ~((COMP_LOOP_acc_19_psp_sva[1:0]!=2'b00) | (~ (fsm_output[0]))
      | (VEC_LOOP_j_sva_11_0[0]) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (VEC_LOOP_j_sva_11_0[1])
      | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[1]) | (~ (fsm_output[10])));
  assign nor_1158_nl = ~((z_out_7[4:1]!=4'b0000) | (~ (fsm_output[3])) | (fsm_output[9])
      | (~ (fsm_output[1])) | (fsm_output[10]));
  assign mux_1115_nl = MUX_s_1_2_2(nor_1158_nl, nor_1148_cse, fsm_output[0]);
  assign mux_1116_nl = MUX_s_1_2_2(nor_1157_nl, mux_1115_nl, fsm_output[8]);
  assign and_655_nl = (fsm_output[7]) & mux_1116_nl;
  assign mux_1117_nl = MUX_s_1_2_2(nor_1156_nl, and_655_nl, fsm_output[6]);
  assign mux_1121_nl = MUX_s_1_2_2(mux_1120_nl, mux_1117_nl, fsm_output[5]);
  assign mux_1128_nl = MUX_s_1_2_2(mux_1127_nl, mux_1121_nl, fsm_output[2]);
  assign or_650_nl = (z_out_7[4:1]!=4'b0000) | (~ (fsm_output[3])) | (fsm_output[9])
      | (~ (fsm_output[1])) | (fsm_output[10]);
  assign or_649_nl = (z_out_7[4:1]!=4'b0000) | (fsm_output[3]) | (~ (fsm_output[9]))
      | (~ (fsm_output[1])) | (fsm_output[10]);
  assign mux_1111_nl = MUX_s_1_2_2(or_650_nl, or_649_nl, fsm_output[0]);
  assign or_648_nl = (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b0000) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (fsm_output[3]) | (fsm_output[9]) | not_tmp_260;
  assign or_646_nl = (COMP_LOOP_acc_16_psp_sva[0]) | (VEC_LOOP_j_sva_11_0[2]) | (VEC_LOOP_j_sva_11_0[0])
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (VEC_LOOP_j_sva_11_0[1]) | (~
      (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[1]) | (fsm_output[10]);
  assign mux_1110_nl = MUX_s_1_2_2(or_648_nl, or_646_nl, fsm_output[0]);
  assign mux_1112_nl = MUX_s_1_2_2(mux_1111_nl, mux_1110_nl, fsm_output[8]);
  assign nor_1160_nl = ~((fsm_output[7:6]!=2'b01) | mux_1112_nl);
  assign nor_1161_nl = ~((fsm_output[8]) | (VEC_LOOP_j_sva_11_0[3]) | (~ (fsm_output[0]))
      | (VEC_LOOP_j_sva_11_0[2:0]!=3'b000) | (fsm_output[3]) | (fsm_output[9]) |
      (fsm_output[1]) | (fsm_output[10]));
  assign or_641_nl = (z_out_7[4:1]!=4'b0000) | (fsm_output[3]) | (fsm_output[9])
      | (fsm_output[1]) | (~ (fsm_output[10]));
  assign mux_1107_nl = MUX_s_1_2_2(or_642_cse, or_641_nl, fsm_output[0]);
  assign nor_1162_nl = ~((fsm_output[8]) | mux_1107_nl);
  assign mux_1108_nl = MUX_s_1_2_2(nor_1161_nl, nor_1162_nl, fsm_output[7]);
  assign nor_1163_nl = ~((~ (fsm_output[8])) | (~ (fsm_output[0])) | (~ (fsm_output[3]))
      | (z_out_7[4:1]!=4'b0000) | (fsm_output[9]) | not_tmp_260);
  assign nor_1164_nl = ~((fsm_output[8]) | (~ (fsm_output[0])) | (VEC_LOOP_j_sva_11_0[0])
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b000)
      | (~ (fsm_output[3])) | (fsm_output[9]) | (~ (fsm_output[1])) | (fsm_output[10]));
  assign mux_1106_nl = MUX_s_1_2_2(nor_1163_nl, nor_1164_nl, fsm_output[7]);
  assign mux_1109_nl = MUX_s_1_2_2(mux_1108_nl, mux_1106_nl, fsm_output[6]);
  assign mux_1113_nl = MUX_s_1_2_2(nor_1160_nl, mux_1109_nl, fsm_output[5]);
  assign or_635_nl = (COMP_LOOP_acc_1_cse_sva[3:0]!=4'b0000) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[0]) | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[1])
      | (~ (fsm_output[10]));
  assign or_633_nl = (z_out_7[4:1]!=4'b0000) | (fsm_output[3]) | (fsm_output[9])
      | not_tmp_260;
  assign mux_1102_nl = MUX_s_1_2_2(or_633_nl, or_642_cse, fsm_output[0]);
  assign mux_1103_nl = MUX_s_1_2_2(or_635_nl, mux_1102_nl, fsm_output[8]);
  assign or_630_nl = (fsm_output[8]) | (fsm_output[0]) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (fsm_output[3]) | (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0000) | (fsm_output[9])
      | (~ (fsm_output[1])) | (fsm_output[10]);
  assign mux_1104_nl = MUX_s_1_2_2(mux_1103_nl, or_630_nl, fsm_output[7]);
  assign nor_1165_nl = ~((fsm_output[6]) | mux_1104_nl);
  assign nor_1166_nl = ~((~ (fsm_output[0])) | (z_out_7[4:1]!=4'b0000) | (~ (fsm_output[3]))
      | (fsm_output[9]) | (~ (fsm_output[1])) | (fsm_output[10]));
  assign nor_1167_nl = ~((COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b0000) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (~ (fsm_output[1])) | (fsm_output[10]));
  assign nor_1168_nl = ~((COMP_LOOP_acc_20_psp_sva[2:0]!=3'b000) | (VEC_LOOP_j_sva_11_0[0])
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[3]) | (fsm_output[9])
      | not_tmp_260);
  assign mux_1099_nl = MUX_s_1_2_2(nor_1167_nl, nor_1168_nl, fsm_output[0]);
  assign mux_1100_nl = MUX_s_1_2_2(nor_1166_nl, mux_1099_nl, fsm_output[8]);
  assign and_656_nl = (fsm_output[7]) & mux_1100_nl;
  assign nor_1169_nl = ~((fsm_output[8:7]!=2'b01) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[0]) | (fsm_output[3]) | (COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b0000)
      | (~ (fsm_output[9])) | (fsm_output[1]) | (fsm_output[10]));
  assign mux_1101_nl = MUX_s_1_2_2(and_656_nl, nor_1169_nl, fsm_output[6]);
  assign mux_1105_nl = MUX_s_1_2_2(nor_1165_nl, mux_1101_nl, fsm_output[5]);
  assign mux_1114_nl = MUX_s_1_2_2(mux_1113_nl, mux_1105_nl, fsm_output[2]);
  assign vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_1128_nl,
      mux_1114_nl, fsm_output[4]);
  assign or_730_nl = (fsm_output[5:4]!=2'b00) | (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b000)
      | (fsm_output[0]) | (~ (VEC_LOOP_j_sva_11_0[0])) | (~ (fsm_output[3])) | (fsm_output[6])
      | (~ (fsm_output[9])) | (fsm_output[8]) | (~ (fsm_output[10]));
  assign or_728_nl = (~ (fsm_output[5])) | (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b000)
      | (fsm_output[0]) | (~ (VEC_LOOP_j_sva_11_0[0])) | (fsm_output[3]) | (~ (fsm_output[6]))
      | (~ (fsm_output[9])) | (fsm_output[8]) | (fsm_output[10]);
  assign mux_1166_nl = MUX_s_1_2_2(or_728_nl, mux_tmp_1152, fsm_output[4]);
  assign mux_1167_nl = MUX_s_1_2_2(or_730_nl, mux_1166_nl, fsm_output[7]);
  assign or_727_nl = (fsm_output[7]) | mux_tmp_1150;
  assign mux_1168_nl = MUX_s_1_2_2(mux_1167_nl, or_727_nl, fsm_output[2]);
  assign or_726_nl = (fsm_output[5:4]!=2'b11) | (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0001)
      | (~ (fsm_output[0])) | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (~ (fsm_output[9]))
      | (fsm_output[8]) | (fsm_output[10]);
  assign or_725_nl = (fsm_output[4]) | mux_tmp_1139;
  assign mux_1164_nl = MUX_s_1_2_2(or_726_nl, or_725_nl, fsm_output[7]);
  assign or_724_nl = (fsm_output[0]) | (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b00) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b01)
      | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[9])) | (fsm_output[8])
      | (fsm_output[10]);
  assign mux_1161_nl = MUX_s_1_2_2(or_724_nl, or_tmp_626, fsm_output[5]);
  assign mux_1162_nl = MUX_s_1_2_2(or_tmp_630, mux_1161_nl, fsm_output[4]);
  assign or_723_nl = (fsm_output[5:4]!=2'b10) | (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0001)
      | (~ (fsm_output[0])) | (fsm_output[3]) | (~ (fsm_output[6])) | (fsm_output[9])
      | (fsm_output[8]) | (fsm_output[10]);
  assign mux_1163_nl = MUX_s_1_2_2(mux_1162_nl, or_723_nl, fsm_output[7]);
  assign mux_1165_nl = MUX_s_1_2_2(mux_1164_nl, mux_1163_nl, fsm_output[2]);
  assign mux_1169_nl = MUX_s_1_2_2(mux_1168_nl, mux_1165_nl, fsm_output[1]);
  assign or_722_nl = (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b000) | (fsm_output[0]) |
      (~ (VEC_LOOP_j_sva_11_0[0])) | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[9]))
      | (fsm_output[8]) | (~ (fsm_output[10]));
  assign mux_1156_nl = MUX_s_1_2_2(or_722_nl, or_622_cse, fsm_output[5]);
  assign mux_1157_nl = MUX_s_1_2_2(mux_1156_nl, or_621_cse, fsm_output[4]);
  assign or_713_nl = (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b000) | (fsm_output[0]) |
      (~ (VEC_LOOP_j_sva_11_0[0])) | (fsm_output[3]) | (~ (fsm_output[6])) | (~ (fsm_output[9]))
      | (fsm_output[8]) | (fsm_output[10]);
  assign mux_1153_nl = MUX_s_1_2_2(or_617_cse, or_713_nl, fsm_output[5]);
  assign mux_1154_nl = MUX_s_1_2_2(mux_1153_nl, mux_tmp_1152, fsm_output[4]);
  assign mux_1158_nl = MUX_s_1_2_2(mux_1157_nl, mux_1154_nl, fsm_output[7]);
  assign mux_1151_nl = MUX_s_1_2_2(mux_tmp_1150, mux_1088_cse, fsm_output[7]);
  assign mux_1159_nl = MUX_s_1_2_2(mux_1158_nl, mux_1151_nl, fsm_output[2]);
  assign or_694_nl = (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0001) | (~ (fsm_output[0]))
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (~ (fsm_output[9])) | (fsm_output[8])
      | (fsm_output[10]);
  assign mux_1141_nl = MUX_s_1_2_2(or_607_cse, or_694_nl, fsm_output[5]);
  assign mux_1142_nl = MUX_s_1_2_2(or_609_cse, mux_1141_nl, fsm_output[4]);
  assign mux_1140_nl = MUX_s_1_2_2(mux_tmp_1139, nand_25_cse, fsm_output[4]);
  assign mux_1143_nl = MUX_s_1_2_2(mux_1142_nl, mux_1140_nl, fsm_output[7]);
  assign or_685_nl = (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b00) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b01)
      | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[9])) | (fsm_output[8])
      | (fsm_output[10]);
  assign mux_1133_nl = MUX_s_1_2_2(or_685_nl, or_601_cse, fsm_output[0]);
  assign mux_1134_nl = MUX_s_1_2_2(mux_1133_nl, or_tmp_626, fsm_output[5]);
  assign mux_1135_nl = MUX_s_1_2_2(or_tmp_630, mux_1134_nl, fsm_output[4]);
  assign or_678_nl = (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0001) | (~ (fsm_output[0]))
      | (fsm_output[3]) | (~ (fsm_output[6])) | (fsm_output[9]) | (fsm_output[8])
      | (fsm_output[10]);
  assign mux_1131_nl = MUX_s_1_2_2(mux_1073_cse, or_678_nl, fsm_output[5]);
  assign mux_1132_nl = MUX_s_1_2_2(mux_1131_nl, or_596_cse, fsm_output[4]);
  assign mux_1136_nl = MUX_s_1_2_2(mux_1135_nl, mux_1132_nl, fsm_output[7]);
  assign mux_1144_nl = MUX_s_1_2_2(mux_1143_nl, mux_1136_nl, fsm_output[2]);
  assign mux_1160_nl = MUX_s_1_2_2(mux_1159_nl, mux_1144_nl, fsm_output[1]);
  assign nor_224_nl = ~((COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0001));
  assign mux_1170_nl = MUX_s_1_2_2(mux_1169_nl, mux_1160_nl, nor_224_nl);
  assign vec_rsc_0_1_i_wea_d_pff = ~ mux_1170_nl;
  assign nor_1123_cse = ~((z_out_7[4:1]!=4'b0001) | (fsm_output[3]) | (~ (fsm_output[9]))
      | (~ (fsm_output[1])) | (fsm_output[10]));
  assign or_748_cse = (z_out_7[4:1]!=4'b0001) | (~ (fsm_output[3])) | (~ (fsm_output[9]))
      | (fsm_output[1]) | (fsm_output[10]);
  assign nor_1122_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b0001) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[0]) | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[1])
      | (~ (fsm_output[10])));
  assign nor_1124_nl = ~((~ (fsm_output[3])) | (z_out_7[4:1]!=4'b0001) | (fsm_output[9])
      | (fsm_output[1]) | (fsm_output[10]));
  assign mux_1197_nl = MUX_s_1_2_2(nor_1123_cse, nor_1124_nl, fsm_output[0]);
  assign mux_1198_nl = MUX_s_1_2_2(nor_1122_nl, mux_1197_nl, fsm_output[8]);
  assign and_651_nl = nor_223_cse & mux_1198_nl;
  assign or_776_nl = (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0001) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (~ (fsm_output[1])) | (fsm_output[10]);
  assign or_775_nl = (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b000) | (~ (VEC_LOOP_j_sva_11_0[0]))
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[3]) | (fsm_output[9])
      | not_tmp_260;
  assign mux_1195_nl = MUX_s_1_2_2(or_776_nl, or_775_nl, fsm_output[0]);
  assign nor_1125_nl = ~((fsm_output[8:7]!=2'b00) | mux_1195_nl);
  assign nor_1126_nl = ~((~ (fsm_output[8])) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b0001) | (fsm_output[0]) | (fsm_output[3])
      | (fsm_output[9]) | (fsm_output[1]) | (fsm_output[10]));
  assign nor_1127_nl = ~((~ (fsm_output[8])) | (fsm_output[0]) | (z_out_7[4:1]!=4'b0001)
      | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[1]) | (~ (fsm_output[10])));
  assign mux_1194_nl = MUX_s_1_2_2(nor_1126_nl, nor_1127_nl, fsm_output[7]);
  assign mux_1196_nl = MUX_s_1_2_2(nor_1125_nl, mux_1194_nl, fsm_output[6]);
  assign mux_1199_nl = MUX_s_1_2_2(and_651_nl, mux_1196_nl, fsm_output[5]);
  assign nor_1128_nl = ~((~ (fsm_output[7])) | (fsm_output[8]) | (~ (fsm_output[0]))
      | (~ (VEC_LOOP_j_sva_11_0[0])) | (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b000) |
      (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (~ (fsm_output[3])) | (~ (fsm_output[9]))
      | (~ (fsm_output[1])) | (fsm_output[10]));
  assign or_767_nl = (z_out_7[4:1]!=4'b0001) | (~ (fsm_output[3])) | (fsm_output[9])
      | (fsm_output[1]) | (~ (fsm_output[10]));
  assign or_765_nl = (fsm_output[3]) | (z_out_7[4:1]!=4'b0001) | (~ (fsm_output[9]))
      | (fsm_output[1]) | (~ (fsm_output[10]));
  assign mux_1190_nl = MUX_s_1_2_2(or_767_nl, or_765_nl, fsm_output[0]);
  assign nor_1129_nl = ~((fsm_output[8]) | mux_1190_nl);
  assign nor_1130_nl = ~((COMP_LOOP_acc_13_psp_sva[1:0]!=2'b00) | (~ (fsm_output[8]))
      | (~ (fsm_output[0])) | (~ (VEC_LOOP_j_sva_11_0[0])) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (VEC_LOOP_j_sva_11_0[1]) | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[1])
      | (fsm_output[10]));
  assign mux_1191_nl = MUX_s_1_2_2(nor_1129_nl, nor_1130_nl, fsm_output[7]);
  assign mux_1192_nl = MUX_s_1_2_2(nor_1128_nl, mux_1191_nl, fsm_output[6]);
  assign nor_1131_nl = ~((fsm_output[8:7]!=2'b10) | (z_out_7[4:1]!=4'b0001) | (fsm_output[0])
      | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[1]) | (fsm_output[10]));
  assign nor_1132_nl = ~((COMP_LOOP_acc_19_psp_sva[1:0]!=2'b00) | (~ (fsm_output[0]))
      | (~ (VEC_LOOP_j_sva_11_0[0])) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) |
      (VEC_LOOP_j_sva_11_0[1]) | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[1])
      | (~ (fsm_output[10])));
  assign nor_1133_nl = ~((z_out_7[4:1]!=4'b0001) | (~ (fsm_output[3])) | (fsm_output[9])
      | (~ (fsm_output[1])) | (fsm_output[10]));
  assign mux_1187_nl = MUX_s_1_2_2(nor_1133_nl, nor_1123_cse, fsm_output[0]);
  assign mux_1188_nl = MUX_s_1_2_2(nor_1132_nl, mux_1187_nl, fsm_output[8]);
  assign and_652_nl = (fsm_output[7]) & mux_1188_nl;
  assign mux_1189_nl = MUX_s_1_2_2(nor_1131_nl, and_652_nl, fsm_output[6]);
  assign mux_1193_nl = MUX_s_1_2_2(mux_1192_nl, mux_1189_nl, fsm_output[5]);
  assign mux_1200_nl = MUX_s_1_2_2(mux_1199_nl, mux_1193_nl, fsm_output[2]);
  assign or_756_nl = (z_out_7[4:1]!=4'b0001) | (~ (fsm_output[3])) | (fsm_output[9])
      | (~ (fsm_output[1])) | (fsm_output[10]);
  assign or_755_nl = (z_out_7[4:1]!=4'b0001) | (fsm_output[3]) | (~ (fsm_output[9]))
      | (~ (fsm_output[1])) | (fsm_output[10]);
  assign mux_1183_nl = MUX_s_1_2_2(or_756_nl, or_755_nl, fsm_output[0]);
  assign or_754_nl = (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b0001) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (fsm_output[3]) | (fsm_output[9]) | not_tmp_260;
  assign or_752_nl = (COMP_LOOP_acc_16_psp_sva[0]) | (VEC_LOOP_j_sva_11_0[2]) | (~
      (VEC_LOOP_j_sva_11_0[0])) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (VEC_LOOP_j_sva_11_0[1])
      | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[1]) | (fsm_output[10]);
  assign mux_1182_nl = MUX_s_1_2_2(or_754_nl, or_752_nl, fsm_output[0]);
  assign mux_1184_nl = MUX_s_1_2_2(mux_1183_nl, mux_1182_nl, fsm_output[8]);
  assign nor_1135_nl = ~((fsm_output[7:6]!=2'b01) | mux_1184_nl);
  assign nor_1136_nl = ~((fsm_output[8]) | (VEC_LOOP_j_sva_11_0[3]) | (~ (fsm_output[0]))
      | (VEC_LOOP_j_sva_11_0[2:0]!=3'b001) | (fsm_output[3]) | (fsm_output[9]) |
      (fsm_output[1]) | (fsm_output[10]));
  assign or_747_nl = (z_out_7[4:1]!=4'b0001) | (fsm_output[3]) | (fsm_output[9])
      | (fsm_output[1]) | (~ (fsm_output[10]));
  assign mux_1179_nl = MUX_s_1_2_2(or_748_cse, or_747_nl, fsm_output[0]);
  assign nor_1137_nl = ~((fsm_output[8]) | mux_1179_nl);
  assign mux_1180_nl = MUX_s_1_2_2(nor_1136_nl, nor_1137_nl, fsm_output[7]);
  assign nor_1138_nl = ~((~ (fsm_output[8])) | (~ (fsm_output[0])) | (~ (fsm_output[3]))
      | (z_out_7[4:1]!=4'b0001) | (fsm_output[9]) | not_tmp_260);
  assign nor_1139_nl = ~((fsm_output[8]) | (~ (fsm_output[0])) | (~ (VEC_LOOP_j_sva_11_0[0]))
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b000)
      | (~ (fsm_output[3])) | (fsm_output[9]) | (~ (fsm_output[1])) | (fsm_output[10]));
  assign mux_1178_nl = MUX_s_1_2_2(nor_1138_nl, nor_1139_nl, fsm_output[7]);
  assign mux_1181_nl = MUX_s_1_2_2(mux_1180_nl, mux_1178_nl, fsm_output[6]);
  assign mux_1185_nl = MUX_s_1_2_2(nor_1135_nl, mux_1181_nl, fsm_output[5]);
  assign or_741_nl = (COMP_LOOP_acc_1_cse_sva[3:0]!=4'b0001) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[0]) | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[1])
      | (~ (fsm_output[10]));
  assign or_739_nl = (z_out_7[4:1]!=4'b0001) | (fsm_output[3]) | (fsm_output[9])
      | not_tmp_260;
  assign mux_1174_nl = MUX_s_1_2_2(or_739_nl, or_748_cse, fsm_output[0]);
  assign mux_1175_nl = MUX_s_1_2_2(or_741_nl, mux_1174_nl, fsm_output[8]);
  assign or_736_nl = (fsm_output[8]) | (fsm_output[0]) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (fsm_output[3]) | (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0001) | (fsm_output[9])
      | (~ (fsm_output[1])) | (fsm_output[10]);
  assign mux_1176_nl = MUX_s_1_2_2(mux_1175_nl, or_736_nl, fsm_output[7]);
  assign nor_1140_nl = ~((fsm_output[6]) | mux_1176_nl);
  assign nor_1141_nl = ~((~ (fsm_output[0])) | (z_out_7[4:1]!=4'b0001) | (~ (fsm_output[3]))
      | (fsm_output[9]) | (~ (fsm_output[1])) | (fsm_output[10]));
  assign nor_1142_nl = ~((COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b0001) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (~ (fsm_output[1])) | (fsm_output[10]));
  assign nor_1143_nl = ~((COMP_LOOP_acc_20_psp_sva[2:0]!=3'b000) | (~ (VEC_LOOP_j_sva_11_0[0]))
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[3]) | (fsm_output[9])
      | not_tmp_260);
  assign mux_1171_nl = MUX_s_1_2_2(nor_1142_nl, nor_1143_nl, fsm_output[0]);
  assign mux_1172_nl = MUX_s_1_2_2(nor_1141_nl, mux_1171_nl, fsm_output[8]);
  assign and_653_nl = (fsm_output[7]) & mux_1172_nl;
  assign nor_1144_nl = ~((fsm_output[8:7]!=2'b01) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[0]) | (fsm_output[3]) | (COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b0001)
      | (~ (fsm_output[9])) | (fsm_output[1]) | (fsm_output[10]));
  assign mux_1173_nl = MUX_s_1_2_2(and_653_nl, nor_1144_nl, fsm_output[6]);
  assign mux_1177_nl = MUX_s_1_2_2(nor_1140_nl, mux_1173_nl, fsm_output[5]);
  assign mux_1186_nl = MUX_s_1_2_2(mux_1185_nl, mux_1177_nl, fsm_output[2]);
  assign vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_1200_nl,
      mux_1186_nl, fsm_output[4]);
  assign or_837_nl = (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b001) | (fsm_output[0]) |
      (VEC_LOOP_j_sva_11_0[0]) | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[9]))
      | (fsm_output[8]) | (~ (fsm_output[10]));
  assign mux_1237_nl = MUX_s_1_2_2(or_837_nl, or_622_cse, fsm_output[5]);
  assign mux_1238_nl = MUX_s_1_2_2(mux_1237_nl, or_621_cse, fsm_output[4]);
  assign or_828_nl = (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b001) | (fsm_output[0]) |
      (VEC_LOOP_j_sva_11_0[0]) | (fsm_output[3]) | (~ (fsm_output[6])) | (~ (fsm_output[9]))
      | (fsm_output[8]) | (fsm_output[10]);
  assign mux_1234_nl = MUX_s_1_2_2(or_617_cse, or_828_nl, fsm_output[5]);
  assign mux_1235_nl = MUX_s_1_2_2(mux_1234_nl, mux_tmp_1212, fsm_output[4]);
  assign mux_1239_nl = MUX_s_1_2_2(mux_1238_nl, mux_1235_nl, fsm_output[7]);
  assign mux_1233_nl = MUX_s_1_2_2(mux_tmp_1211, mux_1088_cse, fsm_output[7]);
  assign mux_1240_nl = MUX_s_1_2_2(mux_1239_nl, mux_1233_nl, fsm_output[2]);
  assign or_818_nl = (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0010) | (~ (fsm_output[0]))
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (~ (fsm_output[9])) | (fsm_output[8])
      | (fsm_output[10]);
  assign mux_1226_nl = MUX_s_1_2_2(or_607_cse, or_818_nl, fsm_output[5]);
  assign mux_1227_nl = MUX_s_1_2_2(or_609_cse, mux_1226_nl, fsm_output[4]);
  assign mux_1225_nl = MUX_s_1_2_2(mux_tmp_1206, nand_25_cse, fsm_output[4]);
  assign mux_1228_nl = MUX_s_1_2_2(mux_1227_nl, mux_1225_nl, fsm_output[7]);
  assign or_815_nl = (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b00) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b10)
      | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[9])) | (fsm_output[8])
      | (fsm_output[10]);
  assign mux_1220_nl = MUX_s_1_2_2(or_815_nl, or_601_cse, fsm_output[0]);
  assign mux_1221_nl = MUX_s_1_2_2(mux_1220_nl, or_tmp_728, fsm_output[5]);
  assign mux_1222_nl = MUX_s_1_2_2(or_tmp_731, mux_1221_nl, fsm_output[4]);
  assign or_810_nl = (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0010) | (~ (fsm_output[0]))
      | (fsm_output[3]) | (~ (fsm_output[6])) | (fsm_output[9]) | (fsm_output[8])
      | (fsm_output[10]);
  assign mux_1218_nl = MUX_s_1_2_2(mux_1073_cse, or_810_nl, fsm_output[5]);
  assign mux_1219_nl = MUX_s_1_2_2(mux_1218_nl, or_596_cse, fsm_output[4]);
  assign mux_1223_nl = MUX_s_1_2_2(mux_1222_nl, mux_1219_nl, fsm_output[7]);
  assign mux_1229_nl = MUX_s_1_2_2(mux_1228_nl, mux_1223_nl, fsm_output[2]);
  assign mux_1241_nl = MUX_s_1_2_2(mux_1240_nl, mux_1229_nl, fsm_output[1]);
  assign or_807_nl = (fsm_output[5:4]!=2'b00) | (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b001)
      | (fsm_output[0]) | (VEC_LOOP_j_sva_11_0[0]) | (~ (fsm_output[3])) | (fsm_output[6])
      | (~ (fsm_output[9])) | (fsm_output[8]) | (~ (fsm_output[10]));
  assign or_805_nl = (~ (fsm_output[5])) | (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b001)
      | (fsm_output[0]) | (VEC_LOOP_j_sva_11_0[0]) | (fsm_output[3]) | (~ (fsm_output[6]))
      | (~ (fsm_output[9])) | (fsm_output[8]) | (fsm_output[10]);
  assign mux_1213_nl = MUX_s_1_2_2(or_805_nl, mux_tmp_1212, fsm_output[4]);
  assign mux_1214_nl = MUX_s_1_2_2(or_807_nl, mux_1213_nl, fsm_output[7]);
  assign or_801_nl = (fsm_output[7]) | mux_tmp_1211;
  assign mux_1215_nl = MUX_s_1_2_2(mux_1214_nl, or_801_nl, fsm_output[2]);
  assign or_794_nl = (fsm_output[5:4]!=2'b11) | (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0010)
      | (~ (fsm_output[0])) | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (~ (fsm_output[9]))
      | (fsm_output[8]) | (fsm_output[10]);
  assign or_793_nl = (fsm_output[4]) | mux_tmp_1206;
  assign mux_1207_nl = MUX_s_1_2_2(or_794_nl, or_793_nl, fsm_output[7]);
  assign or_786_nl = (fsm_output[0]) | (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b00) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b10)
      | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[9])) | (fsm_output[8])
      | (fsm_output[10]);
  assign mux_1202_nl = MUX_s_1_2_2(or_786_nl, or_tmp_728, fsm_output[5]);
  assign mux_1203_nl = MUX_s_1_2_2(or_tmp_731, mux_1202_nl, fsm_output[4]);
  assign or_783_nl = (fsm_output[5:4]!=2'b10) | (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0010)
      | (~ (fsm_output[0])) | (fsm_output[3]) | (~ (fsm_output[6])) | (fsm_output[9])
      | (fsm_output[8]) | (fsm_output[10]);
  assign mux_1204_nl = MUX_s_1_2_2(mux_1203_nl, or_783_nl, fsm_output[7]);
  assign mux_1208_nl = MUX_s_1_2_2(mux_1207_nl, mux_1204_nl, fsm_output[2]);
  assign mux_1216_nl = MUX_s_1_2_2(mux_1215_nl, mux_1208_nl, fsm_output[1]);
  assign or_782_nl = (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0010);
  assign mux_1242_nl = MUX_s_1_2_2(mux_1241_nl, mux_1216_nl, or_782_nl);
  assign vec_rsc_0_2_i_wea_d_pff = ~ mux_1242_nl;
  assign nor_1098_cse = ~((z_out_7[4:1]!=4'b0010) | (fsm_output[3]) | (~ (fsm_output[9]))
      | (~ (fsm_output[1])) | (fsm_output[10]));
  assign or_855_cse = (z_out_7[4:1]!=4'b0010) | (~ (fsm_output[3])) | (~ (fsm_output[9]))
      | (fsm_output[1]) | (fsm_output[10]);
  assign nor_1097_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b0010) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[0]) | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[1])
      | (~ (fsm_output[10])));
  assign nor_1099_nl = ~((~ (fsm_output[3])) | (z_out_7[4:1]!=4'b0010) | (fsm_output[9])
      | (fsm_output[1]) | (fsm_output[10]));
  assign mux_1269_nl = MUX_s_1_2_2(nor_1098_cse, nor_1099_nl, fsm_output[0]);
  assign mux_1270_nl = MUX_s_1_2_2(nor_1097_nl, mux_1269_nl, fsm_output[8]);
  assign and_648_nl = nor_223_cse & mux_1270_nl;
  assign or_883_nl = (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0010) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (~ (fsm_output[1])) | (fsm_output[10]);
  assign or_882_nl = (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b001) | (VEC_LOOP_j_sva_11_0[0])
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[3]) | (fsm_output[9])
      | not_tmp_260;
  assign mux_1267_nl = MUX_s_1_2_2(or_883_nl, or_882_nl, fsm_output[0]);
  assign nor_1100_nl = ~((fsm_output[8:7]!=2'b00) | mux_1267_nl);
  assign nor_1101_nl = ~((~ (fsm_output[8])) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b0010) | (fsm_output[0]) | (fsm_output[3])
      | (fsm_output[9]) | (fsm_output[1]) | (fsm_output[10]));
  assign nor_1102_nl = ~((~ (fsm_output[8])) | (fsm_output[0]) | (z_out_7[4:1]!=4'b0010)
      | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[1]) | (~ (fsm_output[10])));
  assign mux_1266_nl = MUX_s_1_2_2(nor_1101_nl, nor_1102_nl, fsm_output[7]);
  assign mux_1268_nl = MUX_s_1_2_2(nor_1100_nl, mux_1266_nl, fsm_output[6]);
  assign mux_1271_nl = MUX_s_1_2_2(and_648_nl, mux_1268_nl, fsm_output[5]);
  assign nor_1103_nl = ~((~ (fsm_output[7])) | (fsm_output[8]) | (~ (fsm_output[0]))
      | (VEC_LOOP_j_sva_11_0[0]) | (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b001) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (~ (fsm_output[1])) | (fsm_output[10]));
  assign or_874_nl = (z_out_7[4:1]!=4'b0010) | (~ (fsm_output[3])) | (fsm_output[9])
      | (fsm_output[1]) | (~ (fsm_output[10]));
  assign or_872_nl = (fsm_output[3]) | (z_out_7[4:1]!=4'b0010) | (~ (fsm_output[9]))
      | (fsm_output[1]) | (~ (fsm_output[10]));
  assign mux_1262_nl = MUX_s_1_2_2(or_874_nl, or_872_nl, fsm_output[0]);
  assign nor_1104_nl = ~((fsm_output[8]) | mux_1262_nl);
  assign nor_1105_nl = ~((COMP_LOOP_acc_13_psp_sva[1:0]!=2'b00) | (~ (fsm_output[8]))
      | (~ (fsm_output[0])) | (VEC_LOOP_j_sva_11_0[0]) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (~ (VEC_LOOP_j_sva_11_0[1])) | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[1])
      | (fsm_output[10]));
  assign mux_1263_nl = MUX_s_1_2_2(nor_1104_nl, nor_1105_nl, fsm_output[7]);
  assign mux_1264_nl = MUX_s_1_2_2(nor_1103_nl, mux_1263_nl, fsm_output[6]);
  assign nor_1106_nl = ~((fsm_output[8:7]!=2'b10) | (z_out_7[4:1]!=4'b0010) | (fsm_output[0])
      | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[1]) | (fsm_output[10]));
  assign nor_1107_nl = ~((COMP_LOOP_acc_19_psp_sva[1:0]!=2'b00) | (~ (fsm_output[0]))
      | (VEC_LOOP_j_sva_11_0[0]) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (~
      (VEC_LOOP_j_sva_11_0[1])) | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[1])
      | (~ (fsm_output[10])));
  assign nor_1108_nl = ~((z_out_7[4:1]!=4'b0010) | (~ (fsm_output[3])) | (fsm_output[9])
      | (~ (fsm_output[1])) | (fsm_output[10]));
  assign mux_1259_nl = MUX_s_1_2_2(nor_1108_nl, nor_1098_cse, fsm_output[0]);
  assign mux_1260_nl = MUX_s_1_2_2(nor_1107_nl, mux_1259_nl, fsm_output[8]);
  assign and_649_nl = (fsm_output[7]) & mux_1260_nl;
  assign mux_1261_nl = MUX_s_1_2_2(nor_1106_nl, and_649_nl, fsm_output[6]);
  assign mux_1265_nl = MUX_s_1_2_2(mux_1264_nl, mux_1261_nl, fsm_output[5]);
  assign mux_1272_nl = MUX_s_1_2_2(mux_1271_nl, mux_1265_nl, fsm_output[2]);
  assign or_863_nl = (z_out_7[4:1]!=4'b0010) | (~ (fsm_output[3])) | (fsm_output[9])
      | (~ (fsm_output[1])) | (fsm_output[10]);
  assign or_862_nl = (z_out_7[4:1]!=4'b0010) | (fsm_output[3]) | (~ (fsm_output[9]))
      | (~ (fsm_output[1])) | (fsm_output[10]);
  assign mux_1255_nl = MUX_s_1_2_2(or_863_nl, or_862_nl, fsm_output[0]);
  assign or_861_nl = (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b0010) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (fsm_output[3]) | (fsm_output[9]) | not_tmp_260;
  assign or_859_nl = (COMP_LOOP_acc_16_psp_sva[0]) | (VEC_LOOP_j_sva_11_0[2]) | (VEC_LOOP_j_sva_11_0[0])
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (~ (VEC_LOOP_j_sva_11_0[1])) |
      (~ (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[1]) | (fsm_output[10]);
  assign mux_1254_nl = MUX_s_1_2_2(or_861_nl, or_859_nl, fsm_output[0]);
  assign mux_1256_nl = MUX_s_1_2_2(mux_1255_nl, mux_1254_nl, fsm_output[8]);
  assign nor_1110_nl = ~((fsm_output[7:6]!=2'b01) | mux_1256_nl);
  assign nor_1111_nl = ~((fsm_output[8]) | (VEC_LOOP_j_sva_11_0[3]) | (~ (fsm_output[0]))
      | (VEC_LOOP_j_sva_11_0[2:0]!=3'b010) | (fsm_output[3]) | (fsm_output[9]) |
      (fsm_output[1]) | (fsm_output[10]));
  assign or_854_nl = (z_out_7[4:1]!=4'b0010) | (fsm_output[3]) | (fsm_output[9])
      | (fsm_output[1]) | (~ (fsm_output[10]));
  assign mux_1251_nl = MUX_s_1_2_2(or_855_cse, or_854_nl, fsm_output[0]);
  assign nor_1112_nl = ~((fsm_output[8]) | mux_1251_nl);
  assign mux_1252_nl = MUX_s_1_2_2(nor_1111_nl, nor_1112_nl, fsm_output[7]);
  assign nor_1113_nl = ~((~ (fsm_output[8])) | (~ (fsm_output[0])) | (~ (fsm_output[3]))
      | (z_out_7[4:1]!=4'b0010) | (fsm_output[9]) | not_tmp_260);
  assign nor_1114_nl = ~((fsm_output[8]) | (~ (fsm_output[0])) | (VEC_LOOP_j_sva_11_0[0])
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b001)
      | (~ (fsm_output[3])) | (fsm_output[9]) | (~ (fsm_output[1])) | (fsm_output[10]));
  assign mux_1250_nl = MUX_s_1_2_2(nor_1113_nl, nor_1114_nl, fsm_output[7]);
  assign mux_1253_nl = MUX_s_1_2_2(mux_1252_nl, mux_1250_nl, fsm_output[6]);
  assign mux_1257_nl = MUX_s_1_2_2(nor_1110_nl, mux_1253_nl, fsm_output[5]);
  assign or_848_nl = (COMP_LOOP_acc_1_cse_sva[3:0]!=4'b0010) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[0]) | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[1])
      | (~ (fsm_output[10]));
  assign or_846_nl = (z_out_7[4:1]!=4'b0010) | (fsm_output[3]) | (fsm_output[9])
      | not_tmp_260;
  assign mux_1246_nl = MUX_s_1_2_2(or_846_nl, or_855_cse, fsm_output[0]);
  assign mux_1247_nl = MUX_s_1_2_2(or_848_nl, mux_1246_nl, fsm_output[8]);
  assign or_843_nl = (fsm_output[8]) | (fsm_output[0]) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (fsm_output[3]) | (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0010) | (fsm_output[9])
      | (~ (fsm_output[1])) | (fsm_output[10]);
  assign mux_1248_nl = MUX_s_1_2_2(mux_1247_nl, or_843_nl, fsm_output[7]);
  assign nor_1115_nl = ~((fsm_output[6]) | mux_1248_nl);
  assign nor_1116_nl = ~((~ (fsm_output[0])) | (z_out_7[4:1]!=4'b0010) | (~ (fsm_output[3]))
      | (fsm_output[9]) | (~ (fsm_output[1])) | (fsm_output[10]));
  assign nor_1117_nl = ~((COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b0010) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (~ (fsm_output[1])) | (fsm_output[10]));
  assign nor_1118_nl = ~((COMP_LOOP_acc_20_psp_sva[2:0]!=3'b001) | (VEC_LOOP_j_sva_11_0[0])
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[3]) | (fsm_output[9])
      | not_tmp_260);
  assign mux_1243_nl = MUX_s_1_2_2(nor_1117_nl, nor_1118_nl, fsm_output[0]);
  assign mux_1244_nl = MUX_s_1_2_2(nor_1116_nl, mux_1243_nl, fsm_output[8]);
  assign and_650_nl = (fsm_output[7]) & mux_1244_nl;
  assign nor_1119_nl = ~((fsm_output[8:7]!=2'b01) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[0]) | (fsm_output[3]) | (COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b0010)
      | (~ (fsm_output[9])) | (fsm_output[1]) | (fsm_output[10]));
  assign mux_1245_nl = MUX_s_1_2_2(and_650_nl, nor_1119_nl, fsm_output[6]);
  assign mux_1249_nl = MUX_s_1_2_2(nor_1115_nl, mux_1245_nl, fsm_output[5]);
  assign mux_1258_nl = MUX_s_1_2_2(mux_1257_nl, mux_1249_nl, fsm_output[2]);
  assign vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_1272_nl,
      mux_1258_nl, fsm_output[4]);
  assign or_943_nl = (fsm_output[5:4]!=2'b00) | (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b001)
      | (fsm_output[0]) | (~ (VEC_LOOP_j_sva_11_0[0])) | (~ (fsm_output[3])) | (fsm_output[6])
      | (~ (fsm_output[9])) | (fsm_output[8]) | (~ (fsm_output[10]));
  assign or_941_nl = (~ (fsm_output[5])) | (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b001)
      | (fsm_output[0]) | (~ (VEC_LOOP_j_sva_11_0[0])) | (fsm_output[3]) | (~ (fsm_output[6]))
      | (~ (fsm_output[9])) | (fsm_output[8]) | (fsm_output[10]);
  assign mux_1310_nl = MUX_s_1_2_2(or_941_nl, mux_tmp_1296, fsm_output[4]);
  assign mux_1311_nl = MUX_s_1_2_2(or_943_nl, mux_1310_nl, fsm_output[7]);
  assign or_940_nl = (fsm_output[7]) | mux_tmp_1294;
  assign mux_1312_nl = MUX_s_1_2_2(mux_1311_nl, or_940_nl, fsm_output[2]);
  assign or_939_nl = (fsm_output[5:4]!=2'b11) | (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0011)
      | (~ (fsm_output[0])) | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (~ (fsm_output[9]))
      | (fsm_output[8]) | (fsm_output[10]);
  assign or_938_nl = (fsm_output[4]) | mux_tmp_1283;
  assign mux_1308_nl = MUX_s_1_2_2(or_939_nl, or_938_nl, fsm_output[7]);
  assign or_937_nl = (fsm_output[0]) | (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b00) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b11)
      | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[9])) | (fsm_output[8])
      | (fsm_output[10]);
  assign mux_1305_nl = MUX_s_1_2_2(or_937_nl, or_tmp_839, fsm_output[5]);
  assign mux_1306_nl = MUX_s_1_2_2(or_tmp_843, mux_1305_nl, fsm_output[4]);
  assign or_936_nl = (fsm_output[5:4]!=2'b10) | (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0011)
      | (~ (fsm_output[0])) | (fsm_output[3]) | (~ (fsm_output[6])) | (fsm_output[9])
      | (fsm_output[8]) | (fsm_output[10]);
  assign mux_1307_nl = MUX_s_1_2_2(mux_1306_nl, or_936_nl, fsm_output[7]);
  assign mux_1309_nl = MUX_s_1_2_2(mux_1308_nl, mux_1307_nl, fsm_output[2]);
  assign mux_1313_nl = MUX_s_1_2_2(mux_1312_nl, mux_1309_nl, fsm_output[1]);
  assign or_935_nl = (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b001) | (fsm_output[0]) |
      (~ (VEC_LOOP_j_sva_11_0[0])) | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[9]))
      | (fsm_output[8]) | (~ (fsm_output[10]));
  assign mux_1300_nl = MUX_s_1_2_2(or_935_nl, or_622_cse, fsm_output[5]);
  assign mux_1301_nl = MUX_s_1_2_2(mux_1300_nl, or_621_cse, fsm_output[4]);
  assign or_926_nl = (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b001) | (fsm_output[0]) |
      (~ (VEC_LOOP_j_sva_11_0[0])) | (fsm_output[3]) | (~ (fsm_output[6])) | (~ (fsm_output[9]))
      | (fsm_output[8]) | (fsm_output[10]);
  assign mux_1297_nl = MUX_s_1_2_2(or_617_cse, or_926_nl, fsm_output[5]);
  assign mux_1298_nl = MUX_s_1_2_2(mux_1297_nl, mux_tmp_1296, fsm_output[4]);
  assign mux_1302_nl = MUX_s_1_2_2(mux_1301_nl, mux_1298_nl, fsm_output[7]);
  assign mux_1295_nl = MUX_s_1_2_2(mux_tmp_1294, mux_1088_cse, fsm_output[7]);
  assign mux_1303_nl = MUX_s_1_2_2(mux_1302_nl, mux_1295_nl, fsm_output[2]);
  assign or_907_nl = (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0011) | (~ (fsm_output[0]))
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (~ (fsm_output[9])) | (fsm_output[8])
      | (fsm_output[10]);
  assign mux_1285_nl = MUX_s_1_2_2(or_607_cse, or_907_nl, fsm_output[5]);
  assign mux_1286_nl = MUX_s_1_2_2(or_609_cse, mux_1285_nl, fsm_output[4]);
  assign mux_1284_nl = MUX_s_1_2_2(mux_tmp_1283, nand_25_cse, fsm_output[4]);
  assign mux_1287_nl = MUX_s_1_2_2(mux_1286_nl, mux_1284_nl, fsm_output[7]);
  assign or_898_nl = (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b00) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b11)
      | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[9])) | (fsm_output[8])
      | (fsm_output[10]);
  assign mux_1277_nl = MUX_s_1_2_2(or_898_nl, or_601_cse, fsm_output[0]);
  assign mux_1278_nl = MUX_s_1_2_2(mux_1277_nl, or_tmp_839, fsm_output[5]);
  assign mux_1279_nl = MUX_s_1_2_2(or_tmp_843, mux_1278_nl, fsm_output[4]);
  assign or_891_nl = (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0011) | (~ (fsm_output[0]))
      | (fsm_output[3]) | (~ (fsm_output[6])) | (fsm_output[9]) | (fsm_output[8])
      | (fsm_output[10]);
  assign mux_1275_nl = MUX_s_1_2_2(mux_1073_cse, or_891_nl, fsm_output[5]);
  assign mux_1276_nl = MUX_s_1_2_2(mux_1275_nl, or_596_cse, fsm_output[4]);
  assign mux_1280_nl = MUX_s_1_2_2(mux_1279_nl, mux_1276_nl, fsm_output[7]);
  assign mux_1288_nl = MUX_s_1_2_2(mux_1287_nl, mux_1280_nl, fsm_output[2]);
  assign mux_1304_nl = MUX_s_1_2_2(mux_1303_nl, mux_1288_nl, fsm_output[1]);
  assign nor_231_nl = ~((COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0011));
  assign mux_1314_nl = MUX_s_1_2_2(mux_1313_nl, mux_1304_nl, nor_231_nl);
  assign vec_rsc_0_3_i_wea_d_pff = ~ mux_1314_nl;
  assign nor_1073_cse = ~((z_out_7[4:1]!=4'b0011) | (fsm_output[3]) | (~ (fsm_output[9]))
      | (~ (fsm_output[1])) | (fsm_output[10]));
  assign or_961_cse = (z_out_7[4:1]!=4'b0011) | (~ (fsm_output[3])) | (~ (fsm_output[9]))
      | (fsm_output[1]) | (fsm_output[10]);
  assign nor_1072_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b0011) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[0]) | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[1])
      | (~ (fsm_output[10])));
  assign nor_1074_nl = ~((~ (fsm_output[3])) | (z_out_7[4:1]!=4'b0011) | (fsm_output[9])
      | (fsm_output[1]) | (fsm_output[10]));
  assign mux_1341_nl = MUX_s_1_2_2(nor_1073_cse, nor_1074_nl, fsm_output[0]);
  assign mux_1342_nl = MUX_s_1_2_2(nor_1072_nl, mux_1341_nl, fsm_output[8]);
  assign and_645_nl = nor_223_cse & mux_1342_nl;
  assign or_989_nl = (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0011) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (~ (fsm_output[1])) | (fsm_output[10]);
  assign or_988_nl = (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b001) | (~ (VEC_LOOP_j_sva_11_0[0]))
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[3]) | (fsm_output[9])
      | not_tmp_260;
  assign mux_1339_nl = MUX_s_1_2_2(or_989_nl, or_988_nl, fsm_output[0]);
  assign nor_1075_nl = ~((fsm_output[8:7]!=2'b00) | mux_1339_nl);
  assign nor_1076_nl = ~((~ (fsm_output[8])) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b0011) | (fsm_output[0]) | (fsm_output[3])
      | (fsm_output[9]) | (fsm_output[1]) | (fsm_output[10]));
  assign nor_1077_nl = ~((~ (fsm_output[8])) | (fsm_output[0]) | (z_out_7[4:1]!=4'b0011)
      | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[1]) | (~ (fsm_output[10])));
  assign mux_1338_nl = MUX_s_1_2_2(nor_1076_nl, nor_1077_nl, fsm_output[7]);
  assign mux_1340_nl = MUX_s_1_2_2(nor_1075_nl, mux_1338_nl, fsm_output[6]);
  assign mux_1343_nl = MUX_s_1_2_2(and_645_nl, mux_1340_nl, fsm_output[5]);
  assign nor_1078_nl = ~((~ (fsm_output[7])) | (fsm_output[8]) | (~ (fsm_output[0]))
      | (~ (VEC_LOOP_j_sva_11_0[0])) | (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b001) |
      (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (~ (fsm_output[3])) | (~ (fsm_output[9]))
      | (~ (fsm_output[1])) | (fsm_output[10]));
  assign or_980_nl = (z_out_7[4:1]!=4'b0011) | (~ (fsm_output[3])) | (fsm_output[9])
      | (fsm_output[1]) | (~ (fsm_output[10]));
  assign or_978_nl = (fsm_output[3]) | (z_out_7[4:1]!=4'b0011) | (~ (fsm_output[9]))
      | (fsm_output[1]) | (~ (fsm_output[10]));
  assign mux_1334_nl = MUX_s_1_2_2(or_980_nl, or_978_nl, fsm_output[0]);
  assign nor_1079_nl = ~((fsm_output[8]) | mux_1334_nl);
  assign nor_1080_nl = ~((COMP_LOOP_acc_13_psp_sva[1:0]!=2'b00) | (~ (fsm_output[8]))
      | (~ (fsm_output[0])) | (~ (VEC_LOOP_j_sva_11_0[0])) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (~ (VEC_LOOP_j_sva_11_0[1])) | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[1])
      | (fsm_output[10]));
  assign mux_1335_nl = MUX_s_1_2_2(nor_1079_nl, nor_1080_nl, fsm_output[7]);
  assign mux_1336_nl = MUX_s_1_2_2(nor_1078_nl, mux_1335_nl, fsm_output[6]);
  assign nor_1081_nl = ~((fsm_output[8:7]!=2'b10) | (z_out_7[4:1]!=4'b0011) | (fsm_output[0])
      | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[1]) | (fsm_output[10]));
  assign nor_1082_nl = ~((COMP_LOOP_acc_19_psp_sva[1:0]!=2'b00) | (~ (fsm_output[0]))
      | (~ (VEC_LOOP_j_sva_11_0[0])) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) |
      (~ (VEC_LOOP_j_sva_11_0[1])) | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[1])
      | (~ (fsm_output[10])));
  assign nor_1083_nl = ~((z_out_7[4:1]!=4'b0011) | (~ (fsm_output[3])) | (fsm_output[9])
      | (~ (fsm_output[1])) | (fsm_output[10]));
  assign mux_1331_nl = MUX_s_1_2_2(nor_1083_nl, nor_1073_cse, fsm_output[0]);
  assign mux_1332_nl = MUX_s_1_2_2(nor_1082_nl, mux_1331_nl, fsm_output[8]);
  assign and_646_nl = (fsm_output[7]) & mux_1332_nl;
  assign mux_1333_nl = MUX_s_1_2_2(nor_1081_nl, and_646_nl, fsm_output[6]);
  assign mux_1337_nl = MUX_s_1_2_2(mux_1336_nl, mux_1333_nl, fsm_output[5]);
  assign mux_1344_nl = MUX_s_1_2_2(mux_1343_nl, mux_1337_nl, fsm_output[2]);
  assign or_969_nl = (z_out_7[4:1]!=4'b0011) | (~ (fsm_output[3])) | (fsm_output[9])
      | (~ (fsm_output[1])) | (fsm_output[10]);
  assign or_968_nl = (z_out_7[4:1]!=4'b0011) | (fsm_output[3]) | (~ (fsm_output[9]))
      | (~ (fsm_output[1])) | (fsm_output[10]);
  assign mux_1327_nl = MUX_s_1_2_2(or_969_nl, or_968_nl, fsm_output[0]);
  assign or_967_nl = (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b0011) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (fsm_output[3]) | (fsm_output[9]) | not_tmp_260;
  assign or_965_nl = (COMP_LOOP_acc_16_psp_sva[0]) | (VEC_LOOP_j_sva_11_0[2]) | (~
      (VEC_LOOP_j_sva_11_0[0])) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (~ (VEC_LOOP_j_sva_11_0[1]))
      | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[1]) | (fsm_output[10]);
  assign mux_1326_nl = MUX_s_1_2_2(or_967_nl, or_965_nl, fsm_output[0]);
  assign mux_1328_nl = MUX_s_1_2_2(mux_1327_nl, mux_1326_nl, fsm_output[8]);
  assign nor_1085_nl = ~((fsm_output[7:6]!=2'b01) | mux_1328_nl);
  assign nor_1086_nl = ~((fsm_output[8]) | (VEC_LOOP_j_sva_11_0[3]) | (~ (fsm_output[0]))
      | (VEC_LOOP_j_sva_11_0[2:0]!=3'b011) | (fsm_output[3]) | (fsm_output[9]) |
      (fsm_output[1]) | (fsm_output[10]));
  assign or_960_nl = (z_out_7[4:1]!=4'b0011) | (fsm_output[3]) | (fsm_output[9])
      | (fsm_output[1]) | (~ (fsm_output[10]));
  assign mux_1323_nl = MUX_s_1_2_2(or_961_cse, or_960_nl, fsm_output[0]);
  assign nor_1087_nl = ~((fsm_output[8]) | mux_1323_nl);
  assign mux_1324_nl = MUX_s_1_2_2(nor_1086_nl, nor_1087_nl, fsm_output[7]);
  assign nor_1088_nl = ~((~ (fsm_output[8])) | (~ (fsm_output[0])) | (~ (fsm_output[3]))
      | (z_out_7[4:1]!=4'b0011) | (fsm_output[9]) | not_tmp_260);
  assign nor_1089_nl = ~((fsm_output[8]) | (~ (fsm_output[0])) | (~ (VEC_LOOP_j_sva_11_0[0]))
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b001)
      | (~ (fsm_output[3])) | (fsm_output[9]) | (~ (fsm_output[1])) | (fsm_output[10]));
  assign mux_1322_nl = MUX_s_1_2_2(nor_1088_nl, nor_1089_nl, fsm_output[7]);
  assign mux_1325_nl = MUX_s_1_2_2(mux_1324_nl, mux_1322_nl, fsm_output[6]);
  assign mux_1329_nl = MUX_s_1_2_2(nor_1085_nl, mux_1325_nl, fsm_output[5]);
  assign or_954_nl = (COMP_LOOP_acc_1_cse_sva[3:0]!=4'b0011) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[0]) | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[1])
      | (~ (fsm_output[10]));
  assign or_952_nl = (z_out_7[4:1]!=4'b0011) | (fsm_output[3]) | (fsm_output[9])
      | not_tmp_260;
  assign mux_1318_nl = MUX_s_1_2_2(or_952_nl, or_961_cse, fsm_output[0]);
  assign mux_1319_nl = MUX_s_1_2_2(or_954_nl, mux_1318_nl, fsm_output[8]);
  assign or_949_nl = (fsm_output[8]) | (fsm_output[0]) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (fsm_output[3]) | (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0011) | (fsm_output[9])
      | (~ (fsm_output[1])) | (fsm_output[10]);
  assign mux_1320_nl = MUX_s_1_2_2(mux_1319_nl, or_949_nl, fsm_output[7]);
  assign nor_1090_nl = ~((fsm_output[6]) | mux_1320_nl);
  assign nor_1091_nl = ~((~ (fsm_output[0])) | (z_out_7[4:1]!=4'b0011) | (~ (fsm_output[3]))
      | (fsm_output[9]) | (~ (fsm_output[1])) | (fsm_output[10]));
  assign nor_1092_nl = ~((COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b0011) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (~ (fsm_output[1])) | (fsm_output[10]));
  assign nor_1093_nl = ~((COMP_LOOP_acc_20_psp_sva[2:0]!=3'b001) | (~ (VEC_LOOP_j_sva_11_0[0]))
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[3]) | (fsm_output[9])
      | not_tmp_260);
  assign mux_1315_nl = MUX_s_1_2_2(nor_1092_nl, nor_1093_nl, fsm_output[0]);
  assign mux_1316_nl = MUX_s_1_2_2(nor_1091_nl, mux_1315_nl, fsm_output[8]);
  assign and_647_nl = (fsm_output[7]) & mux_1316_nl;
  assign nor_1094_nl = ~((fsm_output[8:7]!=2'b01) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[0]) | (fsm_output[3]) | (COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b0011)
      | (~ (fsm_output[9])) | (fsm_output[1]) | (fsm_output[10]));
  assign mux_1317_nl = MUX_s_1_2_2(and_647_nl, nor_1094_nl, fsm_output[6]);
  assign mux_1321_nl = MUX_s_1_2_2(nor_1090_nl, mux_1317_nl, fsm_output[5]);
  assign mux_1330_nl = MUX_s_1_2_2(mux_1329_nl, mux_1321_nl, fsm_output[2]);
  assign vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_1344_nl,
      mux_1330_nl, fsm_output[4]);
  assign or_1050_nl = (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b010) | (fsm_output[0]) |
      (VEC_LOOP_j_sva_11_0[0]) | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[9]))
      | (fsm_output[8]) | (~ (fsm_output[10]));
  assign mux_1381_nl = MUX_s_1_2_2(or_1050_nl, or_622_cse, fsm_output[5]);
  assign mux_1382_nl = MUX_s_1_2_2(mux_1381_nl, or_621_cse, fsm_output[4]);
  assign or_1041_nl = (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b010) | (fsm_output[0]) |
      (VEC_LOOP_j_sva_11_0[0]) | (fsm_output[3]) | (~ (fsm_output[6])) | (~ (fsm_output[9]))
      | (fsm_output[8]) | (fsm_output[10]);
  assign mux_1378_nl = MUX_s_1_2_2(or_617_cse, or_1041_nl, fsm_output[5]);
  assign mux_1379_nl = MUX_s_1_2_2(mux_1378_nl, mux_tmp_1356, fsm_output[4]);
  assign mux_1383_nl = MUX_s_1_2_2(mux_1382_nl, mux_1379_nl, fsm_output[7]);
  assign mux_1377_nl = MUX_s_1_2_2(mux_tmp_1355, mux_1088_cse, fsm_output[7]);
  assign mux_1384_nl = MUX_s_1_2_2(mux_1383_nl, mux_1377_nl, fsm_output[2]);
  assign or_1031_nl = (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0100) | (~ (fsm_output[0]))
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (~ (fsm_output[9])) | (fsm_output[8])
      | (fsm_output[10]);
  assign mux_1370_nl = MUX_s_1_2_2(or_607_cse, or_1031_nl, fsm_output[5]);
  assign mux_1371_nl = MUX_s_1_2_2(or_609_cse, mux_1370_nl, fsm_output[4]);
  assign mux_1369_nl = MUX_s_1_2_2(mux_tmp_1350, nand_25_cse, fsm_output[4]);
  assign mux_1372_nl = MUX_s_1_2_2(mux_1371_nl, mux_1369_nl, fsm_output[7]);
  assign or_1028_nl = (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b01) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b00)
      | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[9])) | (fsm_output[8])
      | (fsm_output[10]);
  assign mux_1364_nl = MUX_s_1_2_2(or_1028_nl, or_601_cse, fsm_output[0]);
  assign mux_1365_nl = MUX_s_1_2_2(mux_1364_nl, or_tmp_941, fsm_output[5]);
  assign mux_1366_nl = MUX_s_1_2_2(or_tmp_944, mux_1365_nl, fsm_output[4]);
  assign or_1023_nl = (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0100) | (~ (fsm_output[0]))
      | (fsm_output[3]) | (~ (fsm_output[6])) | (fsm_output[9]) | (fsm_output[8])
      | (fsm_output[10]);
  assign mux_1362_nl = MUX_s_1_2_2(mux_1073_cse, or_1023_nl, fsm_output[5]);
  assign mux_1363_nl = MUX_s_1_2_2(mux_1362_nl, or_596_cse, fsm_output[4]);
  assign mux_1367_nl = MUX_s_1_2_2(mux_1366_nl, mux_1363_nl, fsm_output[7]);
  assign mux_1373_nl = MUX_s_1_2_2(mux_1372_nl, mux_1367_nl, fsm_output[2]);
  assign mux_1385_nl = MUX_s_1_2_2(mux_1384_nl, mux_1373_nl, fsm_output[1]);
  assign or_1020_nl = (fsm_output[5:4]!=2'b00) | (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b010)
      | (fsm_output[0]) | (VEC_LOOP_j_sva_11_0[0]) | (~ (fsm_output[3])) | (fsm_output[6])
      | (~ (fsm_output[9])) | (fsm_output[8]) | (~ (fsm_output[10]));
  assign or_1018_nl = (~ (fsm_output[5])) | (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b010)
      | (fsm_output[0]) | (VEC_LOOP_j_sva_11_0[0]) | (fsm_output[3]) | (~ (fsm_output[6]))
      | (~ (fsm_output[9])) | (fsm_output[8]) | (fsm_output[10]);
  assign mux_1357_nl = MUX_s_1_2_2(or_1018_nl, mux_tmp_1356, fsm_output[4]);
  assign mux_1358_nl = MUX_s_1_2_2(or_1020_nl, mux_1357_nl, fsm_output[7]);
  assign or_1014_nl = (fsm_output[7]) | mux_tmp_1355;
  assign mux_1359_nl = MUX_s_1_2_2(mux_1358_nl, or_1014_nl, fsm_output[2]);
  assign or_1007_nl = (fsm_output[5:4]!=2'b11) | (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0100)
      | (~ (fsm_output[0])) | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (~ (fsm_output[9]))
      | (fsm_output[8]) | (fsm_output[10]);
  assign or_1006_nl = (fsm_output[4]) | mux_tmp_1350;
  assign mux_1351_nl = MUX_s_1_2_2(or_1007_nl, or_1006_nl, fsm_output[7]);
  assign or_999_nl = (fsm_output[0]) | (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b01) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b00)
      | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[9])) | (fsm_output[8])
      | (fsm_output[10]);
  assign mux_1346_nl = MUX_s_1_2_2(or_999_nl, or_tmp_941, fsm_output[5]);
  assign mux_1347_nl = MUX_s_1_2_2(or_tmp_944, mux_1346_nl, fsm_output[4]);
  assign or_996_nl = (fsm_output[5:4]!=2'b10) | (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0100)
      | (~ (fsm_output[0])) | (fsm_output[3]) | (~ (fsm_output[6])) | (fsm_output[9])
      | (fsm_output[8]) | (fsm_output[10]);
  assign mux_1348_nl = MUX_s_1_2_2(mux_1347_nl, or_996_nl, fsm_output[7]);
  assign mux_1352_nl = MUX_s_1_2_2(mux_1351_nl, mux_1348_nl, fsm_output[2]);
  assign mux_1360_nl = MUX_s_1_2_2(mux_1359_nl, mux_1352_nl, fsm_output[1]);
  assign or_995_nl = (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0100);
  assign mux_1386_nl = MUX_s_1_2_2(mux_1385_nl, mux_1360_nl, or_995_nl);
  assign vec_rsc_0_4_i_wea_d_pff = ~ mux_1386_nl;
  assign nor_1048_cse = ~((z_out_7[4:1]!=4'b0100) | (fsm_output[3]) | (~ (fsm_output[9]))
      | (~ (fsm_output[1])) | (fsm_output[10]));
  assign or_1068_cse = (z_out_7[4:1]!=4'b0100) | (~ (fsm_output[3])) | (~ (fsm_output[9]))
      | (fsm_output[1]) | (fsm_output[10]);
  assign nor_1047_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b0100) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[0]) | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[1])
      | (~ (fsm_output[10])));
  assign nor_1049_nl = ~((~ (fsm_output[3])) | (z_out_7[4:1]!=4'b0100) | (fsm_output[9])
      | (fsm_output[1]) | (fsm_output[10]));
  assign mux_1413_nl = MUX_s_1_2_2(nor_1048_cse, nor_1049_nl, fsm_output[0]);
  assign mux_1414_nl = MUX_s_1_2_2(nor_1047_nl, mux_1413_nl, fsm_output[8]);
  assign and_642_nl = nor_223_cse & mux_1414_nl;
  assign or_1096_nl = (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0100) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (~ (fsm_output[1])) | (fsm_output[10]);
  assign or_1095_nl = (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b010) | (VEC_LOOP_j_sva_11_0[0])
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[3]) | (fsm_output[9])
      | not_tmp_260;
  assign mux_1411_nl = MUX_s_1_2_2(or_1096_nl, or_1095_nl, fsm_output[0]);
  assign nor_1050_nl = ~((fsm_output[8:7]!=2'b00) | mux_1411_nl);
  assign nor_1051_nl = ~((~ (fsm_output[8])) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b0100) | (fsm_output[0]) | (fsm_output[3])
      | (fsm_output[9]) | (fsm_output[1]) | (fsm_output[10]));
  assign nor_1052_nl = ~((~ (fsm_output[8])) | (fsm_output[0]) | (z_out_7[4:1]!=4'b0100)
      | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[1]) | (~ (fsm_output[10])));
  assign mux_1410_nl = MUX_s_1_2_2(nor_1051_nl, nor_1052_nl, fsm_output[7]);
  assign mux_1412_nl = MUX_s_1_2_2(nor_1050_nl, mux_1410_nl, fsm_output[6]);
  assign mux_1415_nl = MUX_s_1_2_2(and_642_nl, mux_1412_nl, fsm_output[5]);
  assign nor_1053_nl = ~((~ (fsm_output[7])) | (fsm_output[8]) | (~ (fsm_output[0]))
      | (VEC_LOOP_j_sva_11_0[0]) | (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b010) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (~ (fsm_output[1])) | (fsm_output[10]));
  assign or_1087_nl = (z_out_7[4:1]!=4'b0100) | (~ (fsm_output[3])) | (fsm_output[9])
      | (fsm_output[1]) | (~ (fsm_output[10]));
  assign or_1085_nl = (fsm_output[3]) | (z_out_7[4:1]!=4'b0100) | (~ (fsm_output[9]))
      | (fsm_output[1]) | (~ (fsm_output[10]));
  assign mux_1406_nl = MUX_s_1_2_2(or_1087_nl, or_1085_nl, fsm_output[0]);
  assign nor_1054_nl = ~((fsm_output[8]) | mux_1406_nl);
  assign nor_1055_nl = ~((COMP_LOOP_acc_13_psp_sva[1:0]!=2'b01) | (~ (fsm_output[8]))
      | (~ (fsm_output[0])) | (VEC_LOOP_j_sva_11_0[0]) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (VEC_LOOP_j_sva_11_0[1]) | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[1])
      | (fsm_output[10]));
  assign mux_1407_nl = MUX_s_1_2_2(nor_1054_nl, nor_1055_nl, fsm_output[7]);
  assign mux_1408_nl = MUX_s_1_2_2(nor_1053_nl, mux_1407_nl, fsm_output[6]);
  assign nor_1056_nl = ~((fsm_output[8:7]!=2'b10) | (z_out_7[4:1]!=4'b0100) | (fsm_output[0])
      | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[1]) | (fsm_output[10]));
  assign nor_1057_nl = ~((COMP_LOOP_acc_19_psp_sva[1:0]!=2'b01) | (~ (fsm_output[0]))
      | (VEC_LOOP_j_sva_11_0[0]) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (VEC_LOOP_j_sva_11_0[1])
      | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[1]) | (~ (fsm_output[10])));
  assign nor_1058_nl = ~((z_out_7[4:1]!=4'b0100) | (~ (fsm_output[3])) | (fsm_output[9])
      | (~ (fsm_output[1])) | (fsm_output[10]));
  assign mux_1403_nl = MUX_s_1_2_2(nor_1058_nl, nor_1048_cse, fsm_output[0]);
  assign mux_1404_nl = MUX_s_1_2_2(nor_1057_nl, mux_1403_nl, fsm_output[8]);
  assign and_643_nl = (fsm_output[7]) & mux_1404_nl;
  assign mux_1405_nl = MUX_s_1_2_2(nor_1056_nl, and_643_nl, fsm_output[6]);
  assign mux_1409_nl = MUX_s_1_2_2(mux_1408_nl, mux_1405_nl, fsm_output[5]);
  assign mux_1416_nl = MUX_s_1_2_2(mux_1415_nl, mux_1409_nl, fsm_output[2]);
  assign or_1076_nl = (z_out_7[4:1]!=4'b0100) | (~ (fsm_output[3])) | (fsm_output[9])
      | (~ (fsm_output[1])) | (fsm_output[10]);
  assign or_1075_nl = (z_out_7[4:1]!=4'b0100) | (fsm_output[3]) | (~ (fsm_output[9]))
      | (~ (fsm_output[1])) | (fsm_output[10]);
  assign mux_1399_nl = MUX_s_1_2_2(or_1076_nl, or_1075_nl, fsm_output[0]);
  assign or_1074_nl = (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b0100) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (fsm_output[3]) | (fsm_output[9]) | not_tmp_260;
  assign or_1072_nl = (COMP_LOOP_acc_16_psp_sva[0]) | (~ (VEC_LOOP_j_sva_11_0[2]))
      | (VEC_LOOP_j_sva_11_0[0]) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (VEC_LOOP_j_sva_11_0[1])
      | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[1]) | (fsm_output[10]);
  assign mux_1398_nl = MUX_s_1_2_2(or_1074_nl, or_1072_nl, fsm_output[0]);
  assign mux_1400_nl = MUX_s_1_2_2(mux_1399_nl, mux_1398_nl, fsm_output[8]);
  assign nor_1060_nl = ~((fsm_output[7:6]!=2'b01) | mux_1400_nl);
  assign nor_1061_nl = ~((fsm_output[8]) | (VEC_LOOP_j_sva_11_0[3]) | (~ (fsm_output[0]))
      | (VEC_LOOP_j_sva_11_0[2:0]!=3'b100) | (fsm_output[3]) | (fsm_output[9]) |
      (fsm_output[1]) | (fsm_output[10]));
  assign or_1067_nl = (z_out_7[4:1]!=4'b0100) | (fsm_output[3]) | (fsm_output[9])
      | (fsm_output[1]) | (~ (fsm_output[10]));
  assign mux_1395_nl = MUX_s_1_2_2(or_1068_cse, or_1067_nl, fsm_output[0]);
  assign nor_1062_nl = ~((fsm_output[8]) | mux_1395_nl);
  assign mux_1396_nl = MUX_s_1_2_2(nor_1061_nl, nor_1062_nl, fsm_output[7]);
  assign nor_1063_nl = ~((~ (fsm_output[8])) | (~ (fsm_output[0])) | (~ (fsm_output[3]))
      | (z_out_7[4:1]!=4'b0100) | (fsm_output[9]) | not_tmp_260);
  assign nor_1064_nl = ~((fsm_output[8]) | (~ (fsm_output[0])) | (VEC_LOOP_j_sva_11_0[0])
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b010)
      | (~ (fsm_output[3])) | (fsm_output[9]) | (~ (fsm_output[1])) | (fsm_output[10]));
  assign mux_1394_nl = MUX_s_1_2_2(nor_1063_nl, nor_1064_nl, fsm_output[7]);
  assign mux_1397_nl = MUX_s_1_2_2(mux_1396_nl, mux_1394_nl, fsm_output[6]);
  assign mux_1401_nl = MUX_s_1_2_2(nor_1060_nl, mux_1397_nl, fsm_output[5]);
  assign or_1061_nl = (COMP_LOOP_acc_1_cse_sva[3:0]!=4'b0100) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[0]) | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[1])
      | (~ (fsm_output[10]));
  assign or_1059_nl = (z_out_7[4:1]!=4'b0100) | (fsm_output[3]) | (fsm_output[9])
      | not_tmp_260;
  assign mux_1390_nl = MUX_s_1_2_2(or_1059_nl, or_1068_cse, fsm_output[0]);
  assign mux_1391_nl = MUX_s_1_2_2(or_1061_nl, mux_1390_nl, fsm_output[8]);
  assign or_1056_nl = (fsm_output[8]) | (fsm_output[0]) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (fsm_output[3]) | (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0100) | (fsm_output[9])
      | (~ (fsm_output[1])) | (fsm_output[10]);
  assign mux_1392_nl = MUX_s_1_2_2(mux_1391_nl, or_1056_nl, fsm_output[7]);
  assign nor_1065_nl = ~((fsm_output[6]) | mux_1392_nl);
  assign nor_1066_nl = ~((~ (fsm_output[0])) | (z_out_7[4:1]!=4'b0100) | (~ (fsm_output[3]))
      | (fsm_output[9]) | (~ (fsm_output[1])) | (fsm_output[10]));
  assign nor_1067_nl = ~((COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b0100) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (~ (fsm_output[1])) | (fsm_output[10]));
  assign nor_1068_nl = ~((COMP_LOOP_acc_20_psp_sva[2:0]!=3'b010) | (VEC_LOOP_j_sva_11_0[0])
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[3]) | (fsm_output[9])
      | not_tmp_260);
  assign mux_1387_nl = MUX_s_1_2_2(nor_1067_nl, nor_1068_nl, fsm_output[0]);
  assign mux_1388_nl = MUX_s_1_2_2(nor_1066_nl, mux_1387_nl, fsm_output[8]);
  assign and_644_nl = (fsm_output[7]) & mux_1388_nl;
  assign nor_1069_nl = ~((fsm_output[8:7]!=2'b01) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[0]) | (fsm_output[3]) | (COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b0100)
      | (~ (fsm_output[9])) | (fsm_output[1]) | (fsm_output[10]));
  assign mux_1389_nl = MUX_s_1_2_2(and_644_nl, nor_1069_nl, fsm_output[6]);
  assign mux_1393_nl = MUX_s_1_2_2(nor_1065_nl, mux_1389_nl, fsm_output[5]);
  assign mux_1402_nl = MUX_s_1_2_2(mux_1401_nl, mux_1393_nl, fsm_output[2]);
  assign vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_1416_nl,
      mux_1402_nl, fsm_output[4]);
  assign or_1156_nl = (fsm_output[5:4]!=2'b00) | (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b010)
      | (fsm_output[0]) | (~ (VEC_LOOP_j_sva_11_0[0])) | (~ (fsm_output[3])) | (fsm_output[6])
      | (~ (fsm_output[9])) | (fsm_output[8]) | (~ (fsm_output[10]));
  assign or_1154_nl = (~ (fsm_output[5])) | (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b010)
      | (fsm_output[0]) | (~ (VEC_LOOP_j_sva_11_0[0])) | (fsm_output[3]) | (~ (fsm_output[6]))
      | (~ (fsm_output[9])) | (fsm_output[8]) | (fsm_output[10]);
  assign mux_1454_nl = MUX_s_1_2_2(or_1154_nl, mux_tmp_1440, fsm_output[4]);
  assign mux_1455_nl = MUX_s_1_2_2(or_1156_nl, mux_1454_nl, fsm_output[7]);
  assign or_1153_nl = (fsm_output[7]) | mux_tmp_1438;
  assign mux_1456_nl = MUX_s_1_2_2(mux_1455_nl, or_1153_nl, fsm_output[2]);
  assign or_1152_nl = (fsm_output[5:4]!=2'b11) | (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0101)
      | (~ (fsm_output[0])) | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (~ (fsm_output[9]))
      | (fsm_output[8]) | (fsm_output[10]);
  assign or_1151_nl = (fsm_output[4]) | mux_tmp_1427;
  assign mux_1452_nl = MUX_s_1_2_2(or_1152_nl, or_1151_nl, fsm_output[7]);
  assign or_1150_nl = (fsm_output[0]) | (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b01) |
      (VEC_LOOP_j_sva_11_0[1:0]!=2'b01) | (fsm_output[3]) | (fsm_output[6]) | (~
      (fsm_output[9])) | (fsm_output[8]) | (fsm_output[10]);
  assign mux_1449_nl = MUX_s_1_2_2(or_1150_nl, or_tmp_1052, fsm_output[5]);
  assign mux_1450_nl = MUX_s_1_2_2(or_tmp_1056, mux_1449_nl, fsm_output[4]);
  assign or_1149_nl = (fsm_output[5:4]!=2'b10) | (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0101)
      | (~ (fsm_output[0])) | (fsm_output[3]) | (~ (fsm_output[6])) | (fsm_output[9])
      | (fsm_output[8]) | (fsm_output[10]);
  assign mux_1451_nl = MUX_s_1_2_2(mux_1450_nl, or_1149_nl, fsm_output[7]);
  assign mux_1453_nl = MUX_s_1_2_2(mux_1452_nl, mux_1451_nl, fsm_output[2]);
  assign mux_1457_nl = MUX_s_1_2_2(mux_1456_nl, mux_1453_nl, fsm_output[1]);
  assign or_1148_nl = (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b010) | (fsm_output[0]) |
      (~ (VEC_LOOP_j_sva_11_0[0])) | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[9]))
      | (fsm_output[8]) | (~ (fsm_output[10]));
  assign mux_1444_nl = MUX_s_1_2_2(or_1148_nl, or_622_cse, fsm_output[5]);
  assign mux_1445_nl = MUX_s_1_2_2(mux_1444_nl, or_621_cse, fsm_output[4]);
  assign or_1139_nl = (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b010) | (fsm_output[0]) |
      (~ (VEC_LOOP_j_sva_11_0[0])) | (fsm_output[3]) | (~ (fsm_output[6])) | (~ (fsm_output[9]))
      | (fsm_output[8]) | (fsm_output[10]);
  assign mux_1441_nl = MUX_s_1_2_2(or_617_cse, or_1139_nl, fsm_output[5]);
  assign mux_1442_nl = MUX_s_1_2_2(mux_1441_nl, mux_tmp_1440, fsm_output[4]);
  assign mux_1446_nl = MUX_s_1_2_2(mux_1445_nl, mux_1442_nl, fsm_output[7]);
  assign mux_1439_nl = MUX_s_1_2_2(mux_tmp_1438, mux_1088_cse, fsm_output[7]);
  assign mux_1447_nl = MUX_s_1_2_2(mux_1446_nl, mux_1439_nl, fsm_output[2]);
  assign or_1120_nl = (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0101) | (~ (fsm_output[0]))
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (~ (fsm_output[9])) | (fsm_output[8])
      | (fsm_output[10]);
  assign mux_1429_nl = MUX_s_1_2_2(or_607_cse, or_1120_nl, fsm_output[5]);
  assign mux_1430_nl = MUX_s_1_2_2(or_609_cse, mux_1429_nl, fsm_output[4]);
  assign mux_1428_nl = MUX_s_1_2_2(mux_tmp_1427, nand_25_cse, fsm_output[4]);
  assign mux_1431_nl = MUX_s_1_2_2(mux_1430_nl, mux_1428_nl, fsm_output[7]);
  assign or_1111_nl = (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b01) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b01)
      | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[9])) | (fsm_output[8])
      | (fsm_output[10]);
  assign mux_1421_nl = MUX_s_1_2_2(or_1111_nl, or_601_cse, fsm_output[0]);
  assign mux_1422_nl = MUX_s_1_2_2(mux_1421_nl, or_tmp_1052, fsm_output[5]);
  assign mux_1423_nl = MUX_s_1_2_2(or_tmp_1056, mux_1422_nl, fsm_output[4]);
  assign or_1104_nl = (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0101) | (~ (fsm_output[0]))
      | (fsm_output[3]) | (~ (fsm_output[6])) | (fsm_output[9]) | (fsm_output[8])
      | (fsm_output[10]);
  assign mux_1419_nl = MUX_s_1_2_2(mux_1073_cse, or_1104_nl, fsm_output[5]);
  assign mux_1420_nl = MUX_s_1_2_2(mux_1419_nl, or_596_cse, fsm_output[4]);
  assign mux_1424_nl = MUX_s_1_2_2(mux_1423_nl, mux_1420_nl, fsm_output[7]);
  assign mux_1432_nl = MUX_s_1_2_2(mux_1431_nl, mux_1424_nl, fsm_output[2]);
  assign mux_1448_nl = MUX_s_1_2_2(mux_1447_nl, mux_1432_nl, fsm_output[1]);
  assign nor_238_nl = ~((COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0101));
  assign mux_1458_nl = MUX_s_1_2_2(mux_1457_nl, mux_1448_nl, nor_238_nl);
  assign vec_rsc_0_5_i_wea_d_pff = ~ mux_1458_nl;
  assign nor_1023_cse = ~((z_out_7[4:1]!=4'b0101) | (fsm_output[3]) | (~ (fsm_output[9]))
      | (~ (fsm_output[1])) | (fsm_output[10]));
  assign or_1174_cse = (z_out_7[4:1]!=4'b0101) | (~ (fsm_output[3])) | (~ (fsm_output[9]))
      | (fsm_output[1]) | (fsm_output[10]);
  assign nor_1022_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b0101) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[0]) | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[1])
      | (~ (fsm_output[10])));
  assign nor_1024_nl = ~((~ (fsm_output[3])) | (z_out_7[4:1]!=4'b0101) | (fsm_output[9])
      | (fsm_output[1]) | (fsm_output[10]));
  assign mux_1485_nl = MUX_s_1_2_2(nor_1023_cse, nor_1024_nl, fsm_output[0]);
  assign mux_1486_nl = MUX_s_1_2_2(nor_1022_nl, mux_1485_nl, fsm_output[8]);
  assign and_639_nl = nor_223_cse & mux_1486_nl;
  assign or_1202_nl = (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0101) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (~ (fsm_output[1])) | (fsm_output[10]);
  assign or_1201_nl = (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b010) | (~ (VEC_LOOP_j_sva_11_0[0]))
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[3]) | (fsm_output[9])
      | not_tmp_260;
  assign mux_1483_nl = MUX_s_1_2_2(or_1202_nl, or_1201_nl, fsm_output[0]);
  assign nor_1025_nl = ~((fsm_output[8:7]!=2'b00) | mux_1483_nl);
  assign nor_1026_nl = ~((~ (fsm_output[8])) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b0101) | (fsm_output[0]) | (fsm_output[3])
      | (fsm_output[9]) | (fsm_output[1]) | (fsm_output[10]));
  assign nor_1027_nl = ~((~ (fsm_output[8])) | (fsm_output[0]) | (z_out_7[4:1]!=4'b0101)
      | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[1]) | (~ (fsm_output[10])));
  assign mux_1482_nl = MUX_s_1_2_2(nor_1026_nl, nor_1027_nl, fsm_output[7]);
  assign mux_1484_nl = MUX_s_1_2_2(nor_1025_nl, mux_1482_nl, fsm_output[6]);
  assign mux_1487_nl = MUX_s_1_2_2(and_639_nl, mux_1484_nl, fsm_output[5]);
  assign nor_1028_nl = ~((~ (fsm_output[7])) | (fsm_output[8]) | (~ (fsm_output[0]))
      | (~ (VEC_LOOP_j_sva_11_0[0])) | (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b010) |
      (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (~ (fsm_output[3])) | (~ (fsm_output[9]))
      | (~ (fsm_output[1])) | (fsm_output[10]));
  assign or_1193_nl = (z_out_7[4:1]!=4'b0101) | (~ (fsm_output[3])) | (fsm_output[9])
      | (fsm_output[1]) | (~ (fsm_output[10]));
  assign or_1191_nl = (fsm_output[3]) | (z_out_7[4:1]!=4'b0101) | (~ (fsm_output[9]))
      | (fsm_output[1]) | (~ (fsm_output[10]));
  assign mux_1478_nl = MUX_s_1_2_2(or_1193_nl, or_1191_nl, fsm_output[0]);
  assign nor_1029_nl = ~((fsm_output[8]) | mux_1478_nl);
  assign nor_1030_nl = ~((COMP_LOOP_acc_13_psp_sva[1:0]!=2'b01) | (~ (fsm_output[8]))
      | (~ (fsm_output[0])) | (~ (VEC_LOOP_j_sva_11_0[0])) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (VEC_LOOP_j_sva_11_0[1]) | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[1])
      | (fsm_output[10]));
  assign mux_1479_nl = MUX_s_1_2_2(nor_1029_nl, nor_1030_nl, fsm_output[7]);
  assign mux_1480_nl = MUX_s_1_2_2(nor_1028_nl, mux_1479_nl, fsm_output[6]);
  assign nor_1031_nl = ~((fsm_output[8:7]!=2'b10) | (z_out_7[4:1]!=4'b0101) | (fsm_output[0])
      | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[1]) | (fsm_output[10]));
  assign nor_1032_nl = ~((COMP_LOOP_acc_19_psp_sva[1:0]!=2'b01) | (~ (fsm_output[0]))
      | (~ (VEC_LOOP_j_sva_11_0[0])) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) |
      (VEC_LOOP_j_sva_11_0[1]) | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[1])
      | (~ (fsm_output[10])));
  assign nor_1033_nl = ~((z_out_7[4:1]!=4'b0101) | (~ (fsm_output[3])) | (fsm_output[9])
      | (~ (fsm_output[1])) | (fsm_output[10]));
  assign mux_1475_nl = MUX_s_1_2_2(nor_1033_nl, nor_1023_cse, fsm_output[0]);
  assign mux_1476_nl = MUX_s_1_2_2(nor_1032_nl, mux_1475_nl, fsm_output[8]);
  assign and_640_nl = (fsm_output[7]) & mux_1476_nl;
  assign mux_1477_nl = MUX_s_1_2_2(nor_1031_nl, and_640_nl, fsm_output[6]);
  assign mux_1481_nl = MUX_s_1_2_2(mux_1480_nl, mux_1477_nl, fsm_output[5]);
  assign mux_1488_nl = MUX_s_1_2_2(mux_1487_nl, mux_1481_nl, fsm_output[2]);
  assign or_1182_nl = (z_out_7[4:1]!=4'b0101) | (~ (fsm_output[3])) | (fsm_output[9])
      | (~ (fsm_output[1])) | (fsm_output[10]);
  assign or_1181_nl = (z_out_7[4:1]!=4'b0101) | (fsm_output[3]) | (~ (fsm_output[9]))
      | (~ (fsm_output[1])) | (fsm_output[10]);
  assign mux_1471_nl = MUX_s_1_2_2(or_1182_nl, or_1181_nl, fsm_output[0]);
  assign or_1180_nl = (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b0101) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (fsm_output[3]) | (fsm_output[9]) | not_tmp_260;
  assign or_1178_nl = (COMP_LOOP_acc_16_psp_sva[0]) | (~ (VEC_LOOP_j_sva_11_0[2]))
      | (~ (VEC_LOOP_j_sva_11_0[0])) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) |
      (VEC_LOOP_j_sva_11_0[1]) | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[1])
      | (fsm_output[10]);
  assign mux_1470_nl = MUX_s_1_2_2(or_1180_nl, or_1178_nl, fsm_output[0]);
  assign mux_1472_nl = MUX_s_1_2_2(mux_1471_nl, mux_1470_nl, fsm_output[8]);
  assign nor_1035_nl = ~((fsm_output[7:6]!=2'b01) | mux_1472_nl);
  assign nor_1036_nl = ~((fsm_output[8]) | (VEC_LOOP_j_sva_11_0[3]) | (~ (fsm_output[0]))
      | (VEC_LOOP_j_sva_11_0[2:0]!=3'b101) | (fsm_output[3]) | (fsm_output[9]) |
      (fsm_output[1]) | (fsm_output[10]));
  assign or_1173_nl = (z_out_7[4:1]!=4'b0101) | (fsm_output[3]) | (fsm_output[9])
      | (fsm_output[1]) | (~ (fsm_output[10]));
  assign mux_1467_nl = MUX_s_1_2_2(or_1174_cse, or_1173_nl, fsm_output[0]);
  assign nor_1037_nl = ~((fsm_output[8]) | mux_1467_nl);
  assign mux_1468_nl = MUX_s_1_2_2(nor_1036_nl, nor_1037_nl, fsm_output[7]);
  assign nor_1038_nl = ~((~ (fsm_output[8])) | (~ (fsm_output[0])) | (~ (fsm_output[3]))
      | (z_out_7[4:1]!=4'b0101) | (fsm_output[9]) | not_tmp_260);
  assign nor_1039_nl = ~((fsm_output[8]) | (~ (fsm_output[0])) | (~ (VEC_LOOP_j_sva_11_0[0]))
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b010)
      | (~ (fsm_output[3])) | (fsm_output[9]) | (~ (fsm_output[1])) | (fsm_output[10]));
  assign mux_1466_nl = MUX_s_1_2_2(nor_1038_nl, nor_1039_nl, fsm_output[7]);
  assign mux_1469_nl = MUX_s_1_2_2(mux_1468_nl, mux_1466_nl, fsm_output[6]);
  assign mux_1473_nl = MUX_s_1_2_2(nor_1035_nl, mux_1469_nl, fsm_output[5]);
  assign or_1167_nl = (COMP_LOOP_acc_1_cse_sva[3:0]!=4'b0101) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[0]) | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[1])
      | (~ (fsm_output[10]));
  assign or_1165_nl = (z_out_7[4:1]!=4'b0101) | (fsm_output[3]) | (fsm_output[9])
      | not_tmp_260;
  assign mux_1462_nl = MUX_s_1_2_2(or_1165_nl, or_1174_cse, fsm_output[0]);
  assign mux_1463_nl = MUX_s_1_2_2(or_1167_nl, mux_1462_nl, fsm_output[8]);
  assign or_1162_nl = (fsm_output[8]) | (fsm_output[0]) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (fsm_output[3]) | (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0101) | (fsm_output[9])
      | (~ (fsm_output[1])) | (fsm_output[10]);
  assign mux_1464_nl = MUX_s_1_2_2(mux_1463_nl, or_1162_nl, fsm_output[7]);
  assign nor_1040_nl = ~((fsm_output[6]) | mux_1464_nl);
  assign nor_1041_nl = ~((~ (fsm_output[0])) | (z_out_7[4:1]!=4'b0101) | (~ (fsm_output[3]))
      | (fsm_output[9]) | (~ (fsm_output[1])) | (fsm_output[10]));
  assign nor_1042_nl = ~((COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b0101) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (~ (fsm_output[1])) | (fsm_output[10]));
  assign nor_1043_nl = ~((COMP_LOOP_acc_20_psp_sva[2:0]!=3'b010) | (~ (VEC_LOOP_j_sva_11_0[0]))
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[3]) | (fsm_output[9])
      | not_tmp_260);
  assign mux_1459_nl = MUX_s_1_2_2(nor_1042_nl, nor_1043_nl, fsm_output[0]);
  assign mux_1460_nl = MUX_s_1_2_2(nor_1041_nl, mux_1459_nl, fsm_output[8]);
  assign and_641_nl = (fsm_output[7]) & mux_1460_nl;
  assign nor_1044_nl = ~((fsm_output[8:7]!=2'b01) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[0]) | (fsm_output[3]) | (COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b0101)
      | (~ (fsm_output[9])) | (fsm_output[1]) | (fsm_output[10]));
  assign mux_1461_nl = MUX_s_1_2_2(and_641_nl, nor_1044_nl, fsm_output[6]);
  assign mux_1465_nl = MUX_s_1_2_2(nor_1040_nl, mux_1461_nl, fsm_output[5]);
  assign mux_1474_nl = MUX_s_1_2_2(mux_1473_nl, mux_1465_nl, fsm_output[2]);
  assign vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_1488_nl,
      mux_1474_nl, fsm_output[4]);
  assign or_1263_nl = (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b011) | (fsm_output[0]) |
      (VEC_LOOP_j_sva_11_0[0]) | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[9]))
      | (fsm_output[8]) | (~ (fsm_output[10]));
  assign mux_1525_nl = MUX_s_1_2_2(or_1263_nl, or_622_cse, fsm_output[5]);
  assign mux_1526_nl = MUX_s_1_2_2(mux_1525_nl, or_621_cse, fsm_output[4]);
  assign or_1254_nl = (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b011) | (fsm_output[0]) |
      (VEC_LOOP_j_sva_11_0[0]) | (fsm_output[3]) | (~ (fsm_output[6])) | (~ (fsm_output[9]))
      | (fsm_output[8]) | (fsm_output[10]);
  assign mux_1522_nl = MUX_s_1_2_2(or_617_cse, or_1254_nl, fsm_output[5]);
  assign mux_1523_nl = MUX_s_1_2_2(mux_1522_nl, mux_tmp_1500, fsm_output[4]);
  assign mux_1527_nl = MUX_s_1_2_2(mux_1526_nl, mux_1523_nl, fsm_output[7]);
  assign mux_1521_nl = MUX_s_1_2_2(mux_tmp_1499, mux_1088_cse, fsm_output[7]);
  assign mux_1528_nl = MUX_s_1_2_2(mux_1527_nl, mux_1521_nl, fsm_output[2]);
  assign or_1244_nl = (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0110) | (~ (fsm_output[0]))
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (~ (fsm_output[9])) | (fsm_output[8])
      | (fsm_output[10]);
  assign mux_1514_nl = MUX_s_1_2_2(or_607_cse, or_1244_nl, fsm_output[5]);
  assign mux_1515_nl = MUX_s_1_2_2(or_609_cse, mux_1514_nl, fsm_output[4]);
  assign mux_1513_nl = MUX_s_1_2_2(mux_tmp_1494, nand_25_cse, fsm_output[4]);
  assign mux_1516_nl = MUX_s_1_2_2(mux_1515_nl, mux_1513_nl, fsm_output[7]);
  assign or_1241_nl = (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b01) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b10)
      | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[9])) | (fsm_output[8])
      | (fsm_output[10]);
  assign mux_1508_nl = MUX_s_1_2_2(or_1241_nl, or_601_cse, fsm_output[0]);
  assign mux_1509_nl = MUX_s_1_2_2(mux_1508_nl, or_tmp_1154, fsm_output[5]);
  assign mux_1510_nl = MUX_s_1_2_2(or_tmp_1157, mux_1509_nl, fsm_output[4]);
  assign or_1236_nl = (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0110) | (~ (fsm_output[0]))
      | (fsm_output[3]) | (~ (fsm_output[6])) | (fsm_output[9]) | (fsm_output[8])
      | (fsm_output[10]);
  assign mux_1506_nl = MUX_s_1_2_2(mux_1073_cse, or_1236_nl, fsm_output[5]);
  assign mux_1507_nl = MUX_s_1_2_2(mux_1506_nl, or_596_cse, fsm_output[4]);
  assign mux_1511_nl = MUX_s_1_2_2(mux_1510_nl, mux_1507_nl, fsm_output[7]);
  assign mux_1517_nl = MUX_s_1_2_2(mux_1516_nl, mux_1511_nl, fsm_output[2]);
  assign mux_1529_nl = MUX_s_1_2_2(mux_1528_nl, mux_1517_nl, fsm_output[1]);
  assign or_1233_nl = (fsm_output[5:4]!=2'b00) | (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b011)
      | (fsm_output[0]) | (VEC_LOOP_j_sva_11_0[0]) | (~ (fsm_output[3])) | (fsm_output[6])
      | (~ (fsm_output[9])) | (fsm_output[8]) | (~ (fsm_output[10]));
  assign or_1231_nl = (~ (fsm_output[5])) | (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b011)
      | (fsm_output[0]) | (VEC_LOOP_j_sva_11_0[0]) | (fsm_output[3]) | (~ (fsm_output[6]))
      | (~ (fsm_output[9])) | (fsm_output[8]) | (fsm_output[10]);
  assign mux_1501_nl = MUX_s_1_2_2(or_1231_nl, mux_tmp_1500, fsm_output[4]);
  assign mux_1502_nl = MUX_s_1_2_2(or_1233_nl, mux_1501_nl, fsm_output[7]);
  assign or_1227_nl = (fsm_output[7]) | mux_tmp_1499;
  assign mux_1503_nl = MUX_s_1_2_2(mux_1502_nl, or_1227_nl, fsm_output[2]);
  assign or_1220_nl = (fsm_output[5:4]!=2'b11) | (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0110)
      | (~ (fsm_output[0])) | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (~ (fsm_output[9]))
      | (fsm_output[8]) | (fsm_output[10]);
  assign or_1219_nl = (fsm_output[4]) | mux_tmp_1494;
  assign mux_1495_nl = MUX_s_1_2_2(or_1220_nl, or_1219_nl, fsm_output[7]);
  assign or_1212_nl = (fsm_output[0]) | (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b01) |
      (VEC_LOOP_j_sva_11_0[1:0]!=2'b10) | (fsm_output[3]) | (fsm_output[6]) | (~
      (fsm_output[9])) | (fsm_output[8]) | (fsm_output[10]);
  assign mux_1490_nl = MUX_s_1_2_2(or_1212_nl, or_tmp_1154, fsm_output[5]);
  assign mux_1491_nl = MUX_s_1_2_2(or_tmp_1157, mux_1490_nl, fsm_output[4]);
  assign or_1209_nl = (fsm_output[5:4]!=2'b10) | (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0110)
      | (~ (fsm_output[0])) | (fsm_output[3]) | (~ (fsm_output[6])) | (fsm_output[9])
      | (fsm_output[8]) | (fsm_output[10]);
  assign mux_1492_nl = MUX_s_1_2_2(mux_1491_nl, or_1209_nl, fsm_output[7]);
  assign mux_1496_nl = MUX_s_1_2_2(mux_1495_nl, mux_1492_nl, fsm_output[2]);
  assign mux_1504_nl = MUX_s_1_2_2(mux_1503_nl, mux_1496_nl, fsm_output[1]);
  assign or_1208_nl = (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0110);
  assign mux_1530_nl = MUX_s_1_2_2(mux_1529_nl, mux_1504_nl, or_1208_nl);
  assign vec_rsc_0_6_i_wea_d_pff = ~ mux_1530_nl;
  assign nor_998_cse = ~((z_out_7[4:1]!=4'b0110) | (fsm_output[3]) | (~ (fsm_output[9]))
      | (~ (fsm_output[1])) | (fsm_output[10]));
  assign or_1281_cse = (z_out_7[4:1]!=4'b0110) | (~ (fsm_output[3])) | (~ (fsm_output[9]))
      | (fsm_output[1]) | (fsm_output[10]);
  assign nor_997_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b0110) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[0]) | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[1])
      | (~ (fsm_output[10])));
  assign nor_999_nl = ~((~ (fsm_output[3])) | (z_out_7[4:1]!=4'b0110) | (fsm_output[9])
      | (fsm_output[1]) | (fsm_output[10]));
  assign mux_1557_nl = MUX_s_1_2_2(nor_998_cse, nor_999_nl, fsm_output[0]);
  assign mux_1558_nl = MUX_s_1_2_2(nor_997_nl, mux_1557_nl, fsm_output[8]);
  assign and_636_nl = nor_223_cse & mux_1558_nl;
  assign or_1309_nl = (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0110) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (~ (fsm_output[1])) | (fsm_output[10]);
  assign or_1308_nl = (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b011) | (VEC_LOOP_j_sva_11_0[0])
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[3]) | (fsm_output[9])
      | not_tmp_260;
  assign mux_1555_nl = MUX_s_1_2_2(or_1309_nl, or_1308_nl, fsm_output[0]);
  assign nor_1000_nl = ~((fsm_output[8:7]!=2'b00) | mux_1555_nl);
  assign nor_1001_nl = ~((~ (fsm_output[8])) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b0110) | (fsm_output[0]) | (fsm_output[3])
      | (fsm_output[9]) | (fsm_output[1]) | (fsm_output[10]));
  assign nor_1002_nl = ~((~ (fsm_output[8])) | (fsm_output[0]) | (z_out_7[4:1]!=4'b0110)
      | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[1]) | (~ (fsm_output[10])));
  assign mux_1554_nl = MUX_s_1_2_2(nor_1001_nl, nor_1002_nl, fsm_output[7]);
  assign mux_1556_nl = MUX_s_1_2_2(nor_1000_nl, mux_1554_nl, fsm_output[6]);
  assign mux_1559_nl = MUX_s_1_2_2(and_636_nl, mux_1556_nl, fsm_output[5]);
  assign nor_1003_nl = ~((~ (fsm_output[7])) | (fsm_output[8]) | (~ (fsm_output[0]))
      | (VEC_LOOP_j_sva_11_0[0]) | (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b011) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (~ (fsm_output[1])) | (fsm_output[10]));
  assign or_1300_nl = (z_out_7[4:1]!=4'b0110) | (~ (fsm_output[3])) | (fsm_output[9])
      | (fsm_output[1]) | (~ (fsm_output[10]));
  assign or_1298_nl = (fsm_output[3]) | (z_out_7[4:1]!=4'b0110) | (~ (fsm_output[9]))
      | (fsm_output[1]) | (~ (fsm_output[10]));
  assign mux_1550_nl = MUX_s_1_2_2(or_1300_nl, or_1298_nl, fsm_output[0]);
  assign nor_1004_nl = ~((fsm_output[8]) | mux_1550_nl);
  assign nor_1005_nl = ~((COMP_LOOP_acc_13_psp_sva[1:0]!=2'b01) | (~ (fsm_output[8]))
      | (~ (fsm_output[0])) | (VEC_LOOP_j_sva_11_0[0]) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (~ (VEC_LOOP_j_sva_11_0[1])) | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[1])
      | (fsm_output[10]));
  assign mux_1551_nl = MUX_s_1_2_2(nor_1004_nl, nor_1005_nl, fsm_output[7]);
  assign mux_1552_nl = MUX_s_1_2_2(nor_1003_nl, mux_1551_nl, fsm_output[6]);
  assign nor_1006_nl = ~((fsm_output[8:7]!=2'b10) | (z_out_7[4:1]!=4'b0110) | (fsm_output[0])
      | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[1]) | (fsm_output[10]));
  assign nor_1007_nl = ~((COMP_LOOP_acc_19_psp_sva[1:0]!=2'b01) | (~ (fsm_output[0]))
      | (VEC_LOOP_j_sva_11_0[0]) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (~
      (VEC_LOOP_j_sva_11_0[1])) | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[1])
      | (~ (fsm_output[10])));
  assign nor_1008_nl = ~((z_out_7[4:1]!=4'b0110) | (~ (fsm_output[3])) | (fsm_output[9])
      | (~ (fsm_output[1])) | (fsm_output[10]));
  assign mux_1547_nl = MUX_s_1_2_2(nor_1008_nl, nor_998_cse, fsm_output[0]);
  assign mux_1548_nl = MUX_s_1_2_2(nor_1007_nl, mux_1547_nl, fsm_output[8]);
  assign and_637_nl = (fsm_output[7]) & mux_1548_nl;
  assign mux_1549_nl = MUX_s_1_2_2(nor_1006_nl, and_637_nl, fsm_output[6]);
  assign mux_1553_nl = MUX_s_1_2_2(mux_1552_nl, mux_1549_nl, fsm_output[5]);
  assign mux_1560_nl = MUX_s_1_2_2(mux_1559_nl, mux_1553_nl, fsm_output[2]);
  assign or_1289_nl = (z_out_7[4:1]!=4'b0110) | (~ (fsm_output[3])) | (fsm_output[9])
      | (~ (fsm_output[1])) | (fsm_output[10]);
  assign or_1288_nl = (z_out_7[4:1]!=4'b0110) | (fsm_output[3]) | (~ (fsm_output[9]))
      | (~ (fsm_output[1])) | (fsm_output[10]);
  assign mux_1543_nl = MUX_s_1_2_2(or_1289_nl, or_1288_nl, fsm_output[0]);
  assign or_1287_nl = (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b0110) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (fsm_output[3]) | (fsm_output[9]) | not_tmp_260;
  assign or_1285_nl = (COMP_LOOP_acc_16_psp_sva[0]) | (~ (VEC_LOOP_j_sva_11_0[2]))
      | (VEC_LOOP_j_sva_11_0[0]) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (~
      (VEC_LOOP_j_sva_11_0[1])) | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[1])
      | (fsm_output[10]);
  assign mux_1542_nl = MUX_s_1_2_2(or_1287_nl, or_1285_nl, fsm_output[0]);
  assign mux_1544_nl = MUX_s_1_2_2(mux_1543_nl, mux_1542_nl, fsm_output[8]);
  assign nor_1010_nl = ~((fsm_output[7:6]!=2'b01) | mux_1544_nl);
  assign nor_1011_nl = ~((fsm_output[8]) | (VEC_LOOP_j_sva_11_0[3]) | (~ (fsm_output[0]))
      | (VEC_LOOP_j_sva_11_0[2:0]!=3'b110) | (fsm_output[3]) | (fsm_output[9]) |
      (fsm_output[1]) | (fsm_output[10]));
  assign or_1280_nl = (z_out_7[4:1]!=4'b0110) | (fsm_output[3]) | (fsm_output[9])
      | (fsm_output[1]) | (~ (fsm_output[10]));
  assign mux_1539_nl = MUX_s_1_2_2(or_1281_cse, or_1280_nl, fsm_output[0]);
  assign nor_1012_nl = ~((fsm_output[8]) | mux_1539_nl);
  assign mux_1540_nl = MUX_s_1_2_2(nor_1011_nl, nor_1012_nl, fsm_output[7]);
  assign nor_1013_nl = ~((~ (fsm_output[8])) | (~ (fsm_output[0])) | (~ (fsm_output[3]))
      | (z_out_7[4:1]!=4'b0110) | (fsm_output[9]) | not_tmp_260);
  assign nor_1014_nl = ~((fsm_output[8]) | (~ (fsm_output[0])) | (VEC_LOOP_j_sva_11_0[0])
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b011)
      | (~ (fsm_output[3])) | (fsm_output[9]) | (~ (fsm_output[1])) | (fsm_output[10]));
  assign mux_1538_nl = MUX_s_1_2_2(nor_1013_nl, nor_1014_nl, fsm_output[7]);
  assign mux_1541_nl = MUX_s_1_2_2(mux_1540_nl, mux_1538_nl, fsm_output[6]);
  assign mux_1545_nl = MUX_s_1_2_2(nor_1010_nl, mux_1541_nl, fsm_output[5]);
  assign or_1274_nl = (COMP_LOOP_acc_1_cse_sva[3:0]!=4'b0110) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[0]) | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[1])
      | (~ (fsm_output[10]));
  assign or_1272_nl = (z_out_7[4:1]!=4'b0110) | (fsm_output[3]) | (fsm_output[9])
      | not_tmp_260;
  assign mux_1534_nl = MUX_s_1_2_2(or_1272_nl, or_1281_cse, fsm_output[0]);
  assign mux_1535_nl = MUX_s_1_2_2(or_1274_nl, mux_1534_nl, fsm_output[8]);
  assign or_1269_nl = (fsm_output[8]) | (fsm_output[0]) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (fsm_output[3]) | (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0110) | (fsm_output[9])
      | (~ (fsm_output[1])) | (fsm_output[10]);
  assign mux_1536_nl = MUX_s_1_2_2(mux_1535_nl, or_1269_nl, fsm_output[7]);
  assign nor_1015_nl = ~((fsm_output[6]) | mux_1536_nl);
  assign nor_1016_nl = ~((~ (fsm_output[0])) | (z_out_7[4:1]!=4'b0110) | (~ (fsm_output[3]))
      | (fsm_output[9]) | (~ (fsm_output[1])) | (fsm_output[10]));
  assign nor_1017_nl = ~((COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b0110) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (~ (fsm_output[1])) | (fsm_output[10]));
  assign nor_1018_nl = ~((COMP_LOOP_acc_20_psp_sva[2:0]!=3'b011) | (VEC_LOOP_j_sva_11_0[0])
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[3]) | (fsm_output[9])
      | not_tmp_260);
  assign mux_1531_nl = MUX_s_1_2_2(nor_1017_nl, nor_1018_nl, fsm_output[0]);
  assign mux_1532_nl = MUX_s_1_2_2(nor_1016_nl, mux_1531_nl, fsm_output[8]);
  assign and_638_nl = (fsm_output[7]) & mux_1532_nl;
  assign nor_1019_nl = ~((fsm_output[8:7]!=2'b01) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[0]) | (fsm_output[3]) | (COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b0110)
      | (~ (fsm_output[9])) | (fsm_output[1]) | (fsm_output[10]));
  assign mux_1533_nl = MUX_s_1_2_2(and_638_nl, nor_1019_nl, fsm_output[6]);
  assign mux_1537_nl = MUX_s_1_2_2(nor_1015_nl, mux_1533_nl, fsm_output[5]);
  assign mux_1546_nl = MUX_s_1_2_2(mux_1545_nl, mux_1537_nl, fsm_output[2]);
  assign vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_1560_nl,
      mux_1546_nl, fsm_output[4]);
  assign or_1369_nl = (fsm_output[5:4]!=2'b00) | (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b011)
      | (fsm_output[0]) | (~ (VEC_LOOP_j_sva_11_0[0])) | (~ (fsm_output[3])) | (fsm_output[6])
      | (~ (fsm_output[9])) | (fsm_output[8]) | (~ (fsm_output[10]));
  assign or_1367_nl = (~ (fsm_output[5])) | (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b011)
      | (fsm_output[0]) | (~ (VEC_LOOP_j_sva_11_0[0])) | (fsm_output[3]) | (~ (fsm_output[6]))
      | (~ (fsm_output[9])) | (fsm_output[8]) | (fsm_output[10]);
  assign mux_1598_nl = MUX_s_1_2_2(or_1367_nl, mux_tmp_1584, fsm_output[4]);
  assign mux_1599_nl = MUX_s_1_2_2(or_1369_nl, mux_1598_nl, fsm_output[7]);
  assign or_1366_nl = (fsm_output[7]) | mux_tmp_1582;
  assign mux_1600_nl = MUX_s_1_2_2(mux_1599_nl, or_1366_nl, fsm_output[2]);
  assign nand_336_nl = ~((fsm_output[5:4]==2'b11) & (COMP_LOOP_acc_1_cse_6_sva[3:0]==4'b0111)
      & (fsm_output[0]) & (fsm_output[3]) & (fsm_output[6]) & (fsm_output[9]) & (~
      (fsm_output[8])) & (~ (fsm_output[10])));
  assign or_1364_nl = (fsm_output[4]) | mux_tmp_1571;
  assign mux_1596_nl = MUX_s_1_2_2(nand_336_nl, or_1364_nl, fsm_output[7]);
  assign or_1363_nl = (fsm_output[0]) | (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b01) |
      (VEC_LOOP_j_sva_11_0[1:0]!=2'b11) | (fsm_output[3]) | (fsm_output[6]) | (~
      (fsm_output[9])) | (fsm_output[8]) | (fsm_output[10]);
  assign mux_1593_nl = MUX_s_1_2_2(or_1363_nl, or_tmp_1265, fsm_output[5]);
  assign mux_1594_nl = MUX_s_1_2_2(or_tmp_1269, mux_1593_nl, fsm_output[4]);
  assign or_1362_nl = (fsm_output[5:4]!=2'b10) | (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0111)
      | (~ (fsm_output[0])) | (fsm_output[3]) | (~ (fsm_output[6])) | (fsm_output[9])
      | (fsm_output[8]) | (fsm_output[10]);
  assign mux_1595_nl = MUX_s_1_2_2(mux_1594_nl, or_1362_nl, fsm_output[7]);
  assign mux_1597_nl = MUX_s_1_2_2(mux_1596_nl, mux_1595_nl, fsm_output[2]);
  assign mux_1601_nl = MUX_s_1_2_2(mux_1600_nl, mux_1597_nl, fsm_output[1]);
  assign or_1361_nl = (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b011) | (fsm_output[0]) |
      (~ (VEC_LOOP_j_sva_11_0[0])) | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[9]))
      | (fsm_output[8]) | (~ (fsm_output[10]));
  assign mux_1588_nl = MUX_s_1_2_2(or_1361_nl, or_622_cse, fsm_output[5]);
  assign mux_1589_nl = MUX_s_1_2_2(mux_1588_nl, or_621_cse, fsm_output[4]);
  assign or_1352_nl = (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b011) | (fsm_output[0]) |
      (~ (VEC_LOOP_j_sva_11_0[0])) | (fsm_output[3]) | (~ (fsm_output[6])) | (~ (fsm_output[9]))
      | (fsm_output[8]) | (fsm_output[10]);
  assign mux_1585_nl = MUX_s_1_2_2(or_617_cse, or_1352_nl, fsm_output[5]);
  assign mux_1586_nl = MUX_s_1_2_2(mux_1585_nl, mux_tmp_1584, fsm_output[4]);
  assign mux_1590_nl = MUX_s_1_2_2(mux_1589_nl, mux_1586_nl, fsm_output[7]);
  assign mux_1583_nl = MUX_s_1_2_2(mux_tmp_1582, mux_1088_cse, fsm_output[7]);
  assign mux_1591_nl = MUX_s_1_2_2(mux_1590_nl, mux_1583_nl, fsm_output[2]);
  assign nand_338_nl = ~((COMP_LOOP_acc_1_cse_6_sva[3:0]==4'b0111) & (fsm_output[0])
      & (fsm_output[3]) & (fsm_output[6]) & (fsm_output[9]) & (~ (fsm_output[8]))
      & (~ (fsm_output[10])));
  assign mux_1573_nl = MUX_s_1_2_2(or_607_cse, nand_338_nl, fsm_output[5]);
  assign mux_1574_nl = MUX_s_1_2_2(or_609_cse, mux_1573_nl, fsm_output[4]);
  assign mux_1572_nl = MUX_s_1_2_2(mux_tmp_1571, nand_25_cse, fsm_output[4]);
  assign mux_1575_nl = MUX_s_1_2_2(mux_1574_nl, mux_1572_nl, fsm_output[7]);
  assign or_1324_nl = (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b01) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b11)
      | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[9])) | (fsm_output[8])
      | (fsm_output[10]);
  assign mux_1565_nl = MUX_s_1_2_2(or_1324_nl, or_601_cse, fsm_output[0]);
  assign mux_1566_nl = MUX_s_1_2_2(mux_1565_nl, or_tmp_1265, fsm_output[5]);
  assign mux_1567_nl = MUX_s_1_2_2(or_tmp_1269, mux_1566_nl, fsm_output[4]);
  assign or_1317_nl = (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0111) | (~ (fsm_output[0]))
      | (fsm_output[3]) | (~ (fsm_output[6])) | (fsm_output[9]) | (fsm_output[8])
      | (fsm_output[10]);
  assign mux_1563_nl = MUX_s_1_2_2(mux_1073_cse, or_1317_nl, fsm_output[5]);
  assign mux_1564_nl = MUX_s_1_2_2(mux_1563_nl, or_596_cse, fsm_output[4]);
  assign mux_1568_nl = MUX_s_1_2_2(mux_1567_nl, mux_1564_nl, fsm_output[7]);
  assign mux_1576_nl = MUX_s_1_2_2(mux_1575_nl, mux_1568_nl, fsm_output[2]);
  assign mux_1592_nl = MUX_s_1_2_2(mux_1591_nl, mux_1576_nl, fsm_output[1]);
  assign and_635_nl = (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]==4'b0111);
  assign mux_1602_nl = MUX_s_1_2_2(mux_1601_nl, mux_1592_nl, and_635_nl);
  assign vec_rsc_0_7_i_wea_d_pff = ~ mux_1602_nl;
  assign nor_975_cse = ~((z_out_7[4:1]!=4'b0111) | (fsm_output[3]) | (~ (fsm_output[9]))
      | (~ (fsm_output[1])) | (fsm_output[10]));
  assign or_1387_cse = (z_out_7[4:1]!=4'b0111) | (~ (fsm_output[3])) | (~ (fsm_output[9]))
      | (fsm_output[1]) | (fsm_output[10]);
  assign nor_974_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b0111) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[0]) | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[1])
      | (~ (fsm_output[10])));
  assign nor_976_nl = ~((~ (fsm_output[3])) | (z_out_7[4:1]!=4'b0111) | (fsm_output[9])
      | (fsm_output[1]) | (fsm_output[10]));
  assign mux_1629_nl = MUX_s_1_2_2(nor_975_cse, nor_976_nl, fsm_output[0]);
  assign mux_1630_nl = MUX_s_1_2_2(nor_974_nl, mux_1629_nl, fsm_output[8]);
  assign and_630_nl = nor_223_cse & mux_1630_nl;
  assign nand_333_nl = ~((COMP_LOOP_acc_1_cse_6_sva[3:0]==4'b0111) & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm
      & (fsm_output[3]) & (fsm_output[9]) & (fsm_output[1]) & (~ (fsm_output[10])));
  assign or_1414_nl = (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b011) | (~ (VEC_LOOP_j_sva_11_0[0]))
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[3]) | (fsm_output[9])
      | not_tmp_260;
  assign mux_1627_nl = MUX_s_1_2_2(nand_333_nl, or_1414_nl, fsm_output[0]);
  assign nor_977_nl = ~((fsm_output[8:7]!=2'b00) | mux_1627_nl);
  assign nor_978_nl = ~((~ (fsm_output[8])) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b0111) | (fsm_output[0]) | (fsm_output[3])
      | (fsm_output[9]) | (fsm_output[1]) | (fsm_output[10]));
  assign nor_979_nl = ~((~ (fsm_output[8])) | (fsm_output[0]) | (z_out_7[4:1]!=4'b0111)
      | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[1]) | (~ (fsm_output[10])));
  assign mux_1626_nl = MUX_s_1_2_2(nor_978_nl, nor_979_nl, fsm_output[7]);
  assign mux_1628_nl = MUX_s_1_2_2(nor_977_nl, mux_1626_nl, fsm_output[6]);
  assign mux_1631_nl = MUX_s_1_2_2(and_630_nl, mux_1628_nl, fsm_output[5]);
  assign and_631_nl = (fsm_output[7]) & (~ (fsm_output[8])) & (fsm_output[0]) & (VEC_LOOP_j_sva_11_0[0])
      & (COMP_LOOP_acc_14_psp_sva[2:0]==3'b011) & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm
      & (fsm_output[3]) & (fsm_output[9]) & (fsm_output[1]) & (~ (fsm_output[10]));
  assign or_1406_nl = (z_out_7[4:1]!=4'b0111) | (~ (fsm_output[3])) | (fsm_output[9])
      | (fsm_output[1]) | (~ (fsm_output[10]));
  assign or_1404_nl = (fsm_output[3]) | (z_out_7[4:1]!=4'b0111) | (~ (fsm_output[9]))
      | (fsm_output[1]) | (~ (fsm_output[10]));
  assign mux_1622_nl = MUX_s_1_2_2(or_1406_nl, or_1404_nl, fsm_output[0]);
  assign nor_980_nl = ~((fsm_output[8]) | mux_1622_nl);
  assign nor_981_nl = ~((COMP_LOOP_acc_13_psp_sva[1:0]!=2'b01) | (~ (fsm_output[8]))
      | (~ (fsm_output[0])) | (~ (VEC_LOOP_j_sva_11_0[0])) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (~ (VEC_LOOP_j_sva_11_0[1])) | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[1])
      | (fsm_output[10]));
  assign mux_1623_nl = MUX_s_1_2_2(nor_980_nl, nor_981_nl, fsm_output[7]);
  assign mux_1624_nl = MUX_s_1_2_2(and_631_nl, mux_1623_nl, fsm_output[6]);
  assign nor_982_nl = ~((fsm_output[8:7]!=2'b10) | (z_out_7[4:1]!=4'b0111) | (fsm_output[0])
      | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[1]) | (fsm_output[10]));
  assign and_828_nl = (COMP_LOOP_acc_19_psp_sva[1:0]==2'b01) & (fsm_output[0]) &
      (VEC_LOOP_j_sva_11_0[0]) & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm & (VEC_LOOP_j_sva_11_0[1])
      & (fsm_output[3]) & (~ (fsm_output[9])) & (~ (fsm_output[1])) & (fsm_output[10]);
  assign nor_984_nl = ~((z_out_7[4:1]!=4'b0111) | (~ (fsm_output[3])) | (fsm_output[9])
      | (~ (fsm_output[1])) | (fsm_output[10]));
  assign mux_1619_nl = MUX_s_1_2_2(nor_984_nl, nor_975_cse, fsm_output[0]);
  assign mux_1620_nl = MUX_s_1_2_2(and_828_nl, mux_1619_nl, fsm_output[8]);
  assign and_632_nl = (fsm_output[7]) & mux_1620_nl;
  assign mux_1621_nl = MUX_s_1_2_2(nor_982_nl, and_632_nl, fsm_output[6]);
  assign mux_1625_nl = MUX_s_1_2_2(mux_1624_nl, mux_1621_nl, fsm_output[5]);
  assign mux_1632_nl = MUX_s_1_2_2(mux_1631_nl, mux_1625_nl, fsm_output[2]);
  assign or_1395_nl = (z_out_7[4:1]!=4'b0111) | (~ (fsm_output[3])) | (fsm_output[9])
      | (~ (fsm_output[1])) | (fsm_output[10]);
  assign or_1394_nl = (z_out_7[4:1]!=4'b0111) | (fsm_output[3]) | (~ (fsm_output[9]))
      | (~ (fsm_output[1])) | (fsm_output[10]);
  assign mux_1615_nl = MUX_s_1_2_2(or_1395_nl, or_1394_nl, fsm_output[0]);
  assign or_1393_nl = (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b0111) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (fsm_output[3]) | (fsm_output[9]) | not_tmp_260;
  assign or_1391_nl = (COMP_LOOP_acc_16_psp_sva[0]) | (~ (VEC_LOOP_j_sva_11_0[2]))
      | (~ (VEC_LOOP_j_sva_11_0[0])) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) |
      (~ (VEC_LOOP_j_sva_11_0[1])) | (~ (fsm_output[3])) | (~ (fsm_output[9])) |
      (fsm_output[1]) | (fsm_output[10]);
  assign mux_1614_nl = MUX_s_1_2_2(or_1393_nl, or_1391_nl, fsm_output[0]);
  assign mux_1616_nl = MUX_s_1_2_2(mux_1615_nl, mux_1614_nl, fsm_output[8]);
  assign nor_986_nl = ~((fsm_output[7:6]!=2'b01) | mux_1616_nl);
  assign nor_987_nl = ~((fsm_output[8]) | (VEC_LOOP_j_sva_11_0[3]) | (~ (fsm_output[0]))
      | (VEC_LOOP_j_sva_11_0[2:0]!=3'b111) | (fsm_output[3]) | (fsm_output[9]) |
      (fsm_output[1]) | (fsm_output[10]));
  assign or_1386_nl = (z_out_7[4:1]!=4'b0111) | (fsm_output[3]) | (fsm_output[9])
      | (fsm_output[1]) | (~ (fsm_output[10]));
  assign mux_1611_nl = MUX_s_1_2_2(or_1387_cse, or_1386_nl, fsm_output[0]);
  assign nor_988_nl = ~((fsm_output[8]) | mux_1611_nl);
  assign mux_1612_nl = MUX_s_1_2_2(nor_987_nl, nor_988_nl, fsm_output[7]);
  assign nor_989_nl = ~((~((fsm_output[8]) & (fsm_output[0]) & (fsm_output[3]) &
      (z_out_7[4:1]==4'b0111) & (~ (fsm_output[9])))) | not_tmp_260);
  assign nor_990_nl = ~((fsm_output[8]) | (~ (fsm_output[0])) | (~ (VEC_LOOP_j_sva_11_0[0]))
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b011)
      | (~ (fsm_output[3])) | (fsm_output[9]) | (~ (fsm_output[1])) | (fsm_output[10]));
  assign mux_1610_nl = MUX_s_1_2_2(nor_989_nl, nor_990_nl, fsm_output[7]);
  assign mux_1613_nl = MUX_s_1_2_2(mux_1612_nl, mux_1610_nl, fsm_output[6]);
  assign mux_1617_nl = MUX_s_1_2_2(nor_986_nl, mux_1613_nl, fsm_output[5]);
  assign nand_417_nl = ~((COMP_LOOP_acc_1_cse_sva[3:0]==4'b0111) & COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm
      & (~ (fsm_output[0])) & (fsm_output[3]) & (fsm_output[9]) & (~ (fsm_output[1]))
      & (fsm_output[10]));
  assign or_1378_nl = (z_out_7[4:1]!=4'b0111) | (fsm_output[3]) | (fsm_output[9])
      | not_tmp_260;
  assign mux_1606_nl = MUX_s_1_2_2(or_1378_nl, or_1387_cse, fsm_output[0]);
  assign mux_1607_nl = MUX_s_1_2_2(nand_417_nl, mux_1606_nl, fsm_output[8]);
  assign or_1375_nl = (fsm_output[8]) | (fsm_output[0]) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (fsm_output[3]) | (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0111) | (fsm_output[9])
      | (~ (fsm_output[1])) | (fsm_output[10]);
  assign mux_1608_nl = MUX_s_1_2_2(mux_1607_nl, or_1375_nl, fsm_output[7]);
  assign nor_991_nl = ~((fsm_output[6]) | mux_1608_nl);
  assign nor_992_nl = ~((~ (fsm_output[0])) | (z_out_7[4:1]!=4'b0111) | (~ (fsm_output[3]))
      | (fsm_output[9]) | (~ (fsm_output[1])) | (fsm_output[10]));
  assign and_634_nl = (COMP_LOOP_acc_1_cse_10_sva[3:0]==4'b0111) & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm
      & (fsm_output[3]) & (fsm_output[9]) & (fsm_output[1]) & (~ (fsm_output[10]));
  assign nor_993_nl = ~((COMP_LOOP_acc_20_psp_sva[2:0]!=3'b011) | (~ (VEC_LOOP_j_sva_11_0[0]))
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[3]) | (fsm_output[9])
      | not_tmp_260);
  assign mux_1603_nl = MUX_s_1_2_2(and_634_nl, nor_993_nl, fsm_output[0]);
  assign mux_1604_nl = MUX_s_1_2_2(nor_992_nl, mux_1603_nl, fsm_output[8]);
  assign and_633_nl = (fsm_output[7]) & mux_1604_nl;
  assign nor_994_nl = ~((fsm_output[8:7]!=2'b01) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[0]) | (fsm_output[3]) | (COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b0111)
      | (~ (fsm_output[9])) | (fsm_output[1]) | (fsm_output[10]));
  assign mux_1605_nl = MUX_s_1_2_2(and_633_nl, nor_994_nl, fsm_output[6]);
  assign mux_1609_nl = MUX_s_1_2_2(nor_991_nl, mux_1605_nl, fsm_output[5]);
  assign mux_1618_nl = MUX_s_1_2_2(mux_1617_nl, mux_1609_nl, fsm_output[2]);
  assign vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_1632_nl,
      mux_1618_nl, fsm_output[4]);
  assign or_1476_nl = (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b100) | (fsm_output[0]) |
      (VEC_LOOP_j_sva_11_0[0]) | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[9]))
      | (fsm_output[8]) | (~ (fsm_output[10]));
  assign mux_1669_nl = MUX_s_1_2_2(or_1476_nl, or_622_cse, fsm_output[5]);
  assign mux_1670_nl = MUX_s_1_2_2(mux_1669_nl, or_621_cse, fsm_output[4]);
  assign or_1467_nl = (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b100) | (fsm_output[0]) |
      (VEC_LOOP_j_sva_11_0[0]) | (fsm_output[3]) | (~ (fsm_output[6])) | (~ (fsm_output[9]))
      | (fsm_output[8]) | (fsm_output[10]);
  assign mux_1666_nl = MUX_s_1_2_2(or_617_cse, or_1467_nl, fsm_output[5]);
  assign mux_1667_nl = MUX_s_1_2_2(mux_1666_nl, mux_tmp_1644, fsm_output[4]);
  assign mux_1671_nl = MUX_s_1_2_2(mux_1670_nl, mux_1667_nl, fsm_output[7]);
  assign mux_1665_nl = MUX_s_1_2_2(mux_tmp_1643, mux_1088_cse, fsm_output[7]);
  assign mux_1672_nl = MUX_s_1_2_2(mux_1671_nl, mux_1665_nl, fsm_output[2]);
  assign or_1457_nl = (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b1000) | (~ (fsm_output[0]))
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (~ (fsm_output[9])) | (fsm_output[8])
      | (fsm_output[10]);
  assign mux_1658_nl = MUX_s_1_2_2(or_607_cse, or_1457_nl, fsm_output[5]);
  assign mux_1659_nl = MUX_s_1_2_2(or_609_cse, mux_1658_nl, fsm_output[4]);
  assign mux_1657_nl = MUX_s_1_2_2(mux_tmp_1638, nand_25_cse, fsm_output[4]);
  assign mux_1660_nl = MUX_s_1_2_2(mux_1659_nl, mux_1657_nl, fsm_output[7]);
  assign or_1454_nl = (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b10) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b00)
      | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[9])) | (fsm_output[8])
      | (fsm_output[10]);
  assign mux_1652_nl = MUX_s_1_2_2(or_1454_nl, or_601_cse, fsm_output[0]);
  assign mux_1653_nl = MUX_s_1_2_2(mux_1652_nl, or_tmp_1367, fsm_output[5]);
  assign mux_1654_nl = MUX_s_1_2_2(or_tmp_1370, mux_1653_nl, fsm_output[4]);
  assign or_1449_nl = (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1000) | (~ (fsm_output[0]))
      | (fsm_output[3]) | (~ (fsm_output[6])) | (fsm_output[9]) | (fsm_output[8])
      | (fsm_output[10]);
  assign mux_1650_nl = MUX_s_1_2_2(mux_1073_cse, or_1449_nl, fsm_output[5]);
  assign mux_1651_nl = MUX_s_1_2_2(mux_1650_nl, or_596_cse, fsm_output[4]);
  assign mux_1655_nl = MUX_s_1_2_2(mux_1654_nl, mux_1651_nl, fsm_output[7]);
  assign mux_1661_nl = MUX_s_1_2_2(mux_1660_nl, mux_1655_nl, fsm_output[2]);
  assign mux_1673_nl = MUX_s_1_2_2(mux_1672_nl, mux_1661_nl, fsm_output[1]);
  assign or_1446_nl = (fsm_output[5:4]!=2'b00) | (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b100)
      | (fsm_output[0]) | (VEC_LOOP_j_sva_11_0[0]) | (~ (fsm_output[3])) | (fsm_output[6])
      | (~ (fsm_output[9])) | (fsm_output[8]) | (~ (fsm_output[10]));
  assign or_1444_nl = (~ (fsm_output[5])) | (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b100)
      | (fsm_output[0]) | (VEC_LOOP_j_sva_11_0[0]) | (fsm_output[3]) | (~ (fsm_output[6]))
      | (~ (fsm_output[9])) | (fsm_output[8]) | (fsm_output[10]);
  assign mux_1645_nl = MUX_s_1_2_2(or_1444_nl, mux_tmp_1644, fsm_output[4]);
  assign mux_1646_nl = MUX_s_1_2_2(or_1446_nl, mux_1645_nl, fsm_output[7]);
  assign or_1440_nl = (fsm_output[7]) | mux_tmp_1643;
  assign mux_1647_nl = MUX_s_1_2_2(mux_1646_nl, or_1440_nl, fsm_output[2]);
  assign or_1433_nl = (fsm_output[5:4]!=2'b11) | (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b1000)
      | (~ (fsm_output[0])) | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (~ (fsm_output[9]))
      | (fsm_output[8]) | (fsm_output[10]);
  assign or_1432_nl = (fsm_output[4]) | mux_tmp_1638;
  assign mux_1639_nl = MUX_s_1_2_2(or_1433_nl, or_1432_nl, fsm_output[7]);
  assign or_1425_nl = (fsm_output[0]) | (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b10) |
      (VEC_LOOP_j_sva_11_0[1:0]!=2'b00) | (fsm_output[3]) | (fsm_output[6]) | (~
      (fsm_output[9])) | (fsm_output[8]) | (fsm_output[10]);
  assign mux_1634_nl = MUX_s_1_2_2(or_1425_nl, or_tmp_1367, fsm_output[5]);
  assign mux_1635_nl = MUX_s_1_2_2(or_tmp_1370, mux_1634_nl, fsm_output[4]);
  assign or_1422_nl = (fsm_output[5:4]!=2'b10) | (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1000)
      | (~ (fsm_output[0])) | (fsm_output[3]) | (~ (fsm_output[6])) | (fsm_output[9])
      | (fsm_output[8]) | (fsm_output[10]);
  assign mux_1636_nl = MUX_s_1_2_2(mux_1635_nl, or_1422_nl, fsm_output[7]);
  assign mux_1640_nl = MUX_s_1_2_2(mux_1639_nl, mux_1636_nl, fsm_output[2]);
  assign mux_1648_nl = MUX_s_1_2_2(mux_1647_nl, mux_1640_nl, fsm_output[1]);
  assign or_1421_nl = (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b1000);
  assign mux_1674_nl = MUX_s_1_2_2(mux_1673_nl, mux_1648_nl, or_1421_nl);
  assign vec_rsc_0_8_i_wea_d_pff = ~ mux_1674_nl;
  assign nor_950_cse = ~((z_out_7[4:1]!=4'b1000) | (fsm_output[3]) | (~ (fsm_output[9]))
      | (~ (fsm_output[1])) | (fsm_output[10]));
  assign or_1494_cse = (z_out_7[4:1]!=4'b1000) | (~ (fsm_output[3])) | (~ (fsm_output[9]))
      | (fsm_output[1]) | (fsm_output[10]);
  assign nor_949_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b1000) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[0]) | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[1])
      | (~ (fsm_output[10])));
  assign nor_951_nl = ~((~ (fsm_output[3])) | (z_out_7[4:1]!=4'b1000) | (fsm_output[9])
      | (fsm_output[1]) | (fsm_output[10]));
  assign mux_1701_nl = MUX_s_1_2_2(nor_950_cse, nor_951_nl, fsm_output[0]);
  assign mux_1702_nl = MUX_s_1_2_2(nor_949_nl, mux_1701_nl, fsm_output[8]);
  assign and_627_nl = nor_223_cse & mux_1702_nl;
  assign or_1522_nl = (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b1000) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (~ (fsm_output[1])) | (fsm_output[10]);
  assign or_1521_nl = (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b100) | (VEC_LOOP_j_sva_11_0[0])
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[3]) | (fsm_output[9])
      | not_tmp_260;
  assign mux_1699_nl = MUX_s_1_2_2(or_1522_nl, or_1521_nl, fsm_output[0]);
  assign nor_952_nl = ~((fsm_output[8:7]!=2'b00) | mux_1699_nl);
  assign nor_953_nl = ~((~ (fsm_output[8])) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b1000) | (fsm_output[0]) | (fsm_output[3])
      | (fsm_output[9]) | (fsm_output[1]) | (fsm_output[10]));
  assign nor_954_nl = ~((~ (fsm_output[8])) | (fsm_output[0]) | (z_out_7[4:1]!=4'b1000)
      | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[1]) | (~ (fsm_output[10])));
  assign mux_1698_nl = MUX_s_1_2_2(nor_953_nl, nor_954_nl, fsm_output[7]);
  assign mux_1700_nl = MUX_s_1_2_2(nor_952_nl, mux_1698_nl, fsm_output[6]);
  assign mux_1703_nl = MUX_s_1_2_2(and_627_nl, mux_1700_nl, fsm_output[5]);
  assign nor_955_nl = ~((~ (fsm_output[7])) | (fsm_output[8]) | (~ (fsm_output[0]))
      | (VEC_LOOP_j_sva_11_0[0]) | (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b100) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (~ (fsm_output[1])) | (fsm_output[10]));
  assign or_1513_nl = (z_out_7[4:1]!=4'b1000) | (~ (fsm_output[3])) | (fsm_output[9])
      | (fsm_output[1]) | (~ (fsm_output[10]));
  assign or_1511_nl = (fsm_output[3]) | (z_out_7[4:1]!=4'b1000) | (~ (fsm_output[9]))
      | (fsm_output[1]) | (~ (fsm_output[10]));
  assign mux_1694_nl = MUX_s_1_2_2(or_1513_nl, or_1511_nl, fsm_output[0]);
  assign nor_956_nl = ~((fsm_output[8]) | mux_1694_nl);
  assign nor_957_nl = ~((COMP_LOOP_acc_13_psp_sva[1:0]!=2'b10) | (~ (fsm_output[8]))
      | (~ (fsm_output[0])) | (VEC_LOOP_j_sva_11_0[0]) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (VEC_LOOP_j_sva_11_0[1]) | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[1])
      | (fsm_output[10]));
  assign mux_1695_nl = MUX_s_1_2_2(nor_956_nl, nor_957_nl, fsm_output[7]);
  assign mux_1696_nl = MUX_s_1_2_2(nor_955_nl, mux_1695_nl, fsm_output[6]);
  assign nor_958_nl = ~((fsm_output[8:7]!=2'b10) | (z_out_7[4:1]!=4'b1000) | (fsm_output[0])
      | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[1]) | (fsm_output[10]));
  assign nor_959_nl = ~((COMP_LOOP_acc_19_psp_sva[1:0]!=2'b10) | (~ (fsm_output[0]))
      | (VEC_LOOP_j_sva_11_0[0]) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (VEC_LOOP_j_sva_11_0[1])
      | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[1]) | (~ (fsm_output[10])));
  assign nor_960_nl = ~((z_out_7[4:1]!=4'b1000) | (~ (fsm_output[3])) | (fsm_output[9])
      | (~ (fsm_output[1])) | (fsm_output[10]));
  assign mux_1691_nl = MUX_s_1_2_2(nor_960_nl, nor_950_cse, fsm_output[0]);
  assign mux_1692_nl = MUX_s_1_2_2(nor_959_nl, mux_1691_nl, fsm_output[8]);
  assign and_628_nl = (fsm_output[7]) & mux_1692_nl;
  assign mux_1693_nl = MUX_s_1_2_2(nor_958_nl, and_628_nl, fsm_output[6]);
  assign mux_1697_nl = MUX_s_1_2_2(mux_1696_nl, mux_1693_nl, fsm_output[5]);
  assign mux_1704_nl = MUX_s_1_2_2(mux_1703_nl, mux_1697_nl, fsm_output[2]);
  assign or_1502_nl = (z_out_7[4:1]!=4'b1000) | (~ (fsm_output[3])) | (fsm_output[9])
      | (~ (fsm_output[1])) | (fsm_output[10]);
  assign or_1501_nl = (z_out_7[4:1]!=4'b1000) | (fsm_output[3]) | (~ (fsm_output[9]))
      | (~ (fsm_output[1])) | (fsm_output[10]);
  assign mux_1687_nl = MUX_s_1_2_2(or_1502_nl, or_1501_nl, fsm_output[0]);
  assign or_1500_nl = (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b1000) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (fsm_output[3]) | (fsm_output[9]) | not_tmp_260;
  assign or_1498_nl = (~ (COMP_LOOP_acc_16_psp_sva[0])) | (VEC_LOOP_j_sva_11_0[2])
      | (VEC_LOOP_j_sva_11_0[0]) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (VEC_LOOP_j_sva_11_0[1])
      | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[1]) | (fsm_output[10]);
  assign mux_1686_nl = MUX_s_1_2_2(or_1500_nl, or_1498_nl, fsm_output[0]);
  assign mux_1688_nl = MUX_s_1_2_2(mux_1687_nl, mux_1686_nl, fsm_output[8]);
  assign nor_962_nl = ~((fsm_output[7:6]!=2'b01) | mux_1688_nl);
  assign nor_963_nl = ~((fsm_output[8]) | (~ (VEC_LOOP_j_sva_11_0[3])) | (~ (fsm_output[0]))
      | (VEC_LOOP_j_sva_11_0[2:0]!=3'b000) | (fsm_output[3]) | (fsm_output[9]) |
      (fsm_output[1]) | (fsm_output[10]));
  assign or_1493_nl = (z_out_7[4:1]!=4'b1000) | (fsm_output[3]) | (fsm_output[9])
      | (fsm_output[1]) | (~ (fsm_output[10]));
  assign mux_1683_nl = MUX_s_1_2_2(or_1494_cse, or_1493_nl, fsm_output[0]);
  assign nor_964_nl = ~((fsm_output[8]) | mux_1683_nl);
  assign mux_1684_nl = MUX_s_1_2_2(nor_963_nl, nor_964_nl, fsm_output[7]);
  assign nor_965_nl = ~((~ (fsm_output[8])) | (~ (fsm_output[0])) | (~ (fsm_output[3]))
      | (z_out_7[4:1]!=4'b1000) | (fsm_output[9]) | not_tmp_260);
  assign nor_966_nl = ~((fsm_output[8]) | (~ (fsm_output[0])) | (VEC_LOOP_j_sva_11_0[0])
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b100)
      | (~ (fsm_output[3])) | (fsm_output[9]) | (~ (fsm_output[1])) | (fsm_output[10]));
  assign mux_1682_nl = MUX_s_1_2_2(nor_965_nl, nor_966_nl, fsm_output[7]);
  assign mux_1685_nl = MUX_s_1_2_2(mux_1684_nl, mux_1682_nl, fsm_output[6]);
  assign mux_1689_nl = MUX_s_1_2_2(nor_962_nl, mux_1685_nl, fsm_output[5]);
  assign or_1487_nl = (COMP_LOOP_acc_1_cse_sva[3:0]!=4'b1000) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[0]) | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[1])
      | (~ (fsm_output[10]));
  assign or_1485_nl = (z_out_7[4:1]!=4'b1000) | (fsm_output[3]) | (fsm_output[9])
      | not_tmp_260;
  assign mux_1678_nl = MUX_s_1_2_2(or_1485_nl, or_1494_cse, fsm_output[0]);
  assign mux_1679_nl = MUX_s_1_2_2(or_1487_nl, mux_1678_nl, fsm_output[8]);
  assign or_1482_nl = (fsm_output[8]) | (fsm_output[0]) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (fsm_output[3]) | (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1000) | (fsm_output[9])
      | (~ (fsm_output[1])) | (fsm_output[10]);
  assign mux_1680_nl = MUX_s_1_2_2(mux_1679_nl, or_1482_nl, fsm_output[7]);
  assign nor_967_nl = ~((fsm_output[6]) | mux_1680_nl);
  assign nor_968_nl = ~((~ (fsm_output[0])) | (z_out_7[4:1]!=4'b1000) | (~ (fsm_output[3]))
      | (fsm_output[9]) | (~ (fsm_output[1])) | (fsm_output[10]));
  assign nor_969_nl = ~((COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b1000) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (~ (fsm_output[1])) | (fsm_output[10]));
  assign nor_970_nl = ~((COMP_LOOP_acc_20_psp_sva[2:0]!=3'b100) | (VEC_LOOP_j_sva_11_0[0])
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[3]) | (fsm_output[9])
      | not_tmp_260);
  assign mux_1675_nl = MUX_s_1_2_2(nor_969_nl, nor_970_nl, fsm_output[0]);
  assign mux_1676_nl = MUX_s_1_2_2(nor_968_nl, mux_1675_nl, fsm_output[8]);
  assign and_629_nl = (fsm_output[7]) & mux_1676_nl;
  assign nor_971_nl = ~((fsm_output[8:7]!=2'b01) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[0]) | (fsm_output[3]) | (COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b1000)
      | (~ (fsm_output[9])) | (fsm_output[1]) | (fsm_output[10]));
  assign mux_1677_nl = MUX_s_1_2_2(and_629_nl, nor_971_nl, fsm_output[6]);
  assign mux_1681_nl = MUX_s_1_2_2(nor_967_nl, mux_1677_nl, fsm_output[5]);
  assign mux_1690_nl = MUX_s_1_2_2(mux_1689_nl, mux_1681_nl, fsm_output[2]);
  assign vec_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_1704_nl,
      mux_1690_nl, fsm_output[4]);
  assign or_1582_nl = (fsm_output[5:4]!=2'b00) | (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b100)
      | (fsm_output[0]) | (~ (VEC_LOOP_j_sva_11_0[0])) | (~ (fsm_output[3])) | (fsm_output[6])
      | (~ (fsm_output[9])) | (fsm_output[8]) | (~ (fsm_output[10]));
  assign or_1580_nl = (~ (fsm_output[5])) | (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b100)
      | (fsm_output[0]) | (~ (VEC_LOOP_j_sva_11_0[0])) | (fsm_output[3]) | (~ (fsm_output[6]))
      | (~ (fsm_output[9])) | (fsm_output[8]) | (fsm_output[10]);
  assign mux_1742_nl = MUX_s_1_2_2(or_1580_nl, mux_tmp_1728, fsm_output[4]);
  assign mux_1743_nl = MUX_s_1_2_2(or_1582_nl, mux_1742_nl, fsm_output[7]);
  assign or_1579_nl = (fsm_output[7]) | mux_tmp_1726;
  assign mux_1744_nl = MUX_s_1_2_2(mux_1743_nl, or_1579_nl, fsm_output[2]);
  assign or_1578_nl = (fsm_output[5:4]!=2'b11) | (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b1001)
      | (~ (fsm_output[0])) | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (~ (fsm_output[9]))
      | (fsm_output[8]) | (fsm_output[10]);
  assign or_1577_nl = (fsm_output[4]) | mux_tmp_1715;
  assign mux_1740_nl = MUX_s_1_2_2(or_1578_nl, or_1577_nl, fsm_output[7]);
  assign or_1576_nl = (fsm_output[0]) | (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b10) |
      (VEC_LOOP_j_sva_11_0[1:0]!=2'b01) | (fsm_output[3]) | (fsm_output[6]) | (~
      (fsm_output[9])) | (fsm_output[8]) | (fsm_output[10]);
  assign mux_1737_nl = MUX_s_1_2_2(or_1576_nl, or_tmp_1478, fsm_output[5]);
  assign mux_1738_nl = MUX_s_1_2_2(or_tmp_1482, mux_1737_nl, fsm_output[4]);
  assign or_1575_nl = (fsm_output[5:4]!=2'b10) | (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1001)
      | (~ (fsm_output[0])) | (fsm_output[3]) | (~ (fsm_output[6])) | (fsm_output[9])
      | (fsm_output[8]) | (fsm_output[10]);
  assign mux_1739_nl = MUX_s_1_2_2(mux_1738_nl, or_1575_nl, fsm_output[7]);
  assign mux_1741_nl = MUX_s_1_2_2(mux_1740_nl, mux_1739_nl, fsm_output[2]);
  assign mux_1745_nl = MUX_s_1_2_2(mux_1744_nl, mux_1741_nl, fsm_output[1]);
  assign or_1574_nl = (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b100) | (fsm_output[0]) |
      (~ (VEC_LOOP_j_sva_11_0[0])) | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[9]))
      | (fsm_output[8]) | (~ (fsm_output[10]));
  assign mux_1732_nl = MUX_s_1_2_2(or_1574_nl, or_622_cse, fsm_output[5]);
  assign mux_1733_nl = MUX_s_1_2_2(mux_1732_nl, or_621_cse, fsm_output[4]);
  assign or_1565_nl = (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b100) | (fsm_output[0]) |
      (~ (VEC_LOOP_j_sva_11_0[0])) | (fsm_output[3]) | (~ (fsm_output[6])) | (~ (fsm_output[9]))
      | (fsm_output[8]) | (fsm_output[10]);
  assign mux_1729_nl = MUX_s_1_2_2(or_617_cse, or_1565_nl, fsm_output[5]);
  assign mux_1730_nl = MUX_s_1_2_2(mux_1729_nl, mux_tmp_1728, fsm_output[4]);
  assign mux_1734_nl = MUX_s_1_2_2(mux_1733_nl, mux_1730_nl, fsm_output[7]);
  assign mux_1727_nl = MUX_s_1_2_2(mux_tmp_1726, mux_1088_cse, fsm_output[7]);
  assign mux_1735_nl = MUX_s_1_2_2(mux_1734_nl, mux_1727_nl, fsm_output[2]);
  assign or_1546_nl = (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b1001) | (~ (fsm_output[0]))
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (~ (fsm_output[9])) | (fsm_output[8])
      | (fsm_output[10]);
  assign mux_1717_nl = MUX_s_1_2_2(or_607_cse, or_1546_nl, fsm_output[5]);
  assign mux_1718_nl = MUX_s_1_2_2(or_609_cse, mux_1717_nl, fsm_output[4]);
  assign mux_1716_nl = MUX_s_1_2_2(mux_tmp_1715, nand_25_cse, fsm_output[4]);
  assign mux_1719_nl = MUX_s_1_2_2(mux_1718_nl, mux_1716_nl, fsm_output[7]);
  assign or_1537_nl = (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b10) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b01)
      | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[9])) | (fsm_output[8])
      | (fsm_output[10]);
  assign mux_1709_nl = MUX_s_1_2_2(or_1537_nl, or_601_cse, fsm_output[0]);
  assign mux_1710_nl = MUX_s_1_2_2(mux_1709_nl, or_tmp_1478, fsm_output[5]);
  assign mux_1711_nl = MUX_s_1_2_2(or_tmp_1482, mux_1710_nl, fsm_output[4]);
  assign or_1530_nl = (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1001) | (~ (fsm_output[0]))
      | (fsm_output[3]) | (~ (fsm_output[6])) | (fsm_output[9]) | (fsm_output[8])
      | (fsm_output[10]);
  assign mux_1707_nl = MUX_s_1_2_2(mux_1073_cse, or_1530_nl, fsm_output[5]);
  assign mux_1708_nl = MUX_s_1_2_2(mux_1707_nl, or_596_cse, fsm_output[4]);
  assign mux_1712_nl = MUX_s_1_2_2(mux_1711_nl, mux_1708_nl, fsm_output[7]);
  assign mux_1720_nl = MUX_s_1_2_2(mux_1719_nl, mux_1712_nl, fsm_output[2]);
  assign mux_1736_nl = MUX_s_1_2_2(mux_1735_nl, mux_1720_nl, fsm_output[1]);
  assign nor_252_nl = ~((COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b1001));
  assign mux_1746_nl = MUX_s_1_2_2(mux_1745_nl, mux_1736_nl, nor_252_nl);
  assign vec_rsc_0_9_i_wea_d_pff = ~ mux_1746_nl;
  assign nor_925_cse = ~((z_out_7[4:1]!=4'b1001) | (fsm_output[3]) | (~ (fsm_output[9]))
      | (~ (fsm_output[1])) | (fsm_output[10]));
  assign or_1600_cse = (z_out_7[4:1]!=4'b1001) | (~ (fsm_output[3])) | (~ (fsm_output[9]))
      | (fsm_output[1]) | (fsm_output[10]);
  assign nor_924_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b1001) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[0]) | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[1])
      | (~ (fsm_output[10])));
  assign nor_926_nl = ~((~ (fsm_output[3])) | (z_out_7[4:1]!=4'b1001) | (fsm_output[9])
      | (fsm_output[1]) | (fsm_output[10]));
  assign mux_1773_nl = MUX_s_1_2_2(nor_925_cse, nor_926_nl, fsm_output[0]);
  assign mux_1774_nl = MUX_s_1_2_2(nor_924_nl, mux_1773_nl, fsm_output[8]);
  assign and_624_nl = nor_223_cse & mux_1774_nl;
  assign or_1628_nl = (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b1001) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (~ (fsm_output[1])) | (fsm_output[10]);
  assign or_1627_nl = (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b100) | (~ (VEC_LOOP_j_sva_11_0[0]))
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[3]) | (fsm_output[9])
      | not_tmp_260;
  assign mux_1771_nl = MUX_s_1_2_2(or_1628_nl, or_1627_nl, fsm_output[0]);
  assign nor_927_nl = ~((fsm_output[8:7]!=2'b00) | mux_1771_nl);
  assign nor_928_nl = ~((~ (fsm_output[8])) | (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b1001)
      | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) | (fsm_output[0]) | (fsm_output[3])
      | (fsm_output[9]) | (fsm_output[1]) | (fsm_output[10]));
  assign nor_929_nl = ~((~ (fsm_output[8])) | (fsm_output[0]) | (z_out_7[4:1]!=4'b1001)
      | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[1]) | (~ (fsm_output[10])));
  assign mux_1770_nl = MUX_s_1_2_2(nor_928_nl, nor_929_nl, fsm_output[7]);
  assign mux_1772_nl = MUX_s_1_2_2(nor_927_nl, mux_1770_nl, fsm_output[6]);
  assign mux_1775_nl = MUX_s_1_2_2(and_624_nl, mux_1772_nl, fsm_output[5]);
  assign nor_930_nl = ~((~ (fsm_output[7])) | (fsm_output[8]) | (~ (fsm_output[0]))
      | (~ (VEC_LOOP_j_sva_11_0[0])) | (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b100) |
      (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (~ (fsm_output[3])) | (~ (fsm_output[9]))
      | (~ (fsm_output[1])) | (fsm_output[10]));
  assign or_1619_nl = (z_out_7[4:1]!=4'b1001) | (~ (fsm_output[3])) | (fsm_output[9])
      | (fsm_output[1]) | (~ (fsm_output[10]));
  assign or_1617_nl = (fsm_output[3]) | (z_out_7[4:1]!=4'b1001) | (~ (fsm_output[9]))
      | (fsm_output[1]) | (~ (fsm_output[10]));
  assign mux_1766_nl = MUX_s_1_2_2(or_1619_nl, or_1617_nl, fsm_output[0]);
  assign nor_931_nl = ~((fsm_output[8]) | mux_1766_nl);
  assign nor_932_nl = ~((COMP_LOOP_acc_13_psp_sva[1:0]!=2'b10) | (~ (fsm_output[8]))
      | (~ (fsm_output[0])) | (~ (VEC_LOOP_j_sva_11_0[0])) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (VEC_LOOP_j_sva_11_0[1]) | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[1])
      | (fsm_output[10]));
  assign mux_1767_nl = MUX_s_1_2_2(nor_931_nl, nor_932_nl, fsm_output[7]);
  assign mux_1768_nl = MUX_s_1_2_2(nor_930_nl, mux_1767_nl, fsm_output[6]);
  assign nor_933_nl = ~((fsm_output[8:7]!=2'b10) | (z_out_7[4:1]!=4'b1001) | (fsm_output[0])
      | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[1]) | (fsm_output[10]));
  assign nor_934_nl = ~((COMP_LOOP_acc_19_psp_sva[1:0]!=2'b10) | (~ (fsm_output[0]))
      | (~ (VEC_LOOP_j_sva_11_0[0])) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) |
      (VEC_LOOP_j_sva_11_0[1]) | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[1])
      | (~ (fsm_output[10])));
  assign nor_935_nl = ~((z_out_7[4:1]!=4'b1001) | (~ (fsm_output[3])) | (fsm_output[9])
      | (~ (fsm_output[1])) | (fsm_output[10]));
  assign mux_1763_nl = MUX_s_1_2_2(nor_935_nl, nor_925_cse, fsm_output[0]);
  assign mux_1764_nl = MUX_s_1_2_2(nor_934_nl, mux_1763_nl, fsm_output[8]);
  assign and_625_nl = (fsm_output[7]) & mux_1764_nl;
  assign mux_1765_nl = MUX_s_1_2_2(nor_933_nl, and_625_nl, fsm_output[6]);
  assign mux_1769_nl = MUX_s_1_2_2(mux_1768_nl, mux_1765_nl, fsm_output[5]);
  assign mux_1776_nl = MUX_s_1_2_2(mux_1775_nl, mux_1769_nl, fsm_output[2]);
  assign or_1608_nl = (z_out_7[4:1]!=4'b1001) | (~ (fsm_output[3])) | (fsm_output[9])
      | (~ (fsm_output[1])) | (fsm_output[10]);
  assign or_1607_nl = (z_out_7[4:1]!=4'b1001) | (fsm_output[3]) | (~ (fsm_output[9]))
      | (~ (fsm_output[1])) | (fsm_output[10]);
  assign mux_1759_nl = MUX_s_1_2_2(or_1608_nl, or_1607_nl, fsm_output[0]);
  assign or_1606_nl = (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b1001) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (fsm_output[3]) | (fsm_output[9]) | not_tmp_260;
  assign or_1604_nl = (~ (COMP_LOOP_acc_16_psp_sva[0])) | (VEC_LOOP_j_sva_11_0[2])
      | (~ (VEC_LOOP_j_sva_11_0[0])) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) |
      (VEC_LOOP_j_sva_11_0[1]) | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[1])
      | (fsm_output[10]);
  assign mux_1758_nl = MUX_s_1_2_2(or_1606_nl, or_1604_nl, fsm_output[0]);
  assign mux_1760_nl = MUX_s_1_2_2(mux_1759_nl, mux_1758_nl, fsm_output[8]);
  assign nor_937_nl = ~((fsm_output[7:6]!=2'b01) | mux_1760_nl);
  assign nor_938_nl = ~((fsm_output[8]) | (~ (VEC_LOOP_j_sva_11_0[3])) | (~ (fsm_output[0]))
      | (VEC_LOOP_j_sva_11_0[2:0]!=3'b001) | (fsm_output[3]) | (fsm_output[9]) |
      (fsm_output[1]) | (fsm_output[10]));
  assign or_1599_nl = (z_out_7[4:1]!=4'b1001) | (fsm_output[3]) | (fsm_output[9])
      | (fsm_output[1]) | (~ (fsm_output[10]));
  assign mux_1755_nl = MUX_s_1_2_2(or_1600_cse, or_1599_nl, fsm_output[0]);
  assign nor_939_nl = ~((fsm_output[8]) | mux_1755_nl);
  assign mux_1756_nl = MUX_s_1_2_2(nor_938_nl, nor_939_nl, fsm_output[7]);
  assign nor_940_nl = ~((~ (fsm_output[8])) | (~ (fsm_output[0])) | (~ (fsm_output[3]))
      | (z_out_7[4:1]!=4'b1001) | (fsm_output[9]) | not_tmp_260);
  assign nor_941_nl = ~((fsm_output[8]) | (~ (fsm_output[0])) | (~ (VEC_LOOP_j_sva_11_0[0]))
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b100)
      | (~ (fsm_output[3])) | (fsm_output[9]) | (~ (fsm_output[1])) | (fsm_output[10]));
  assign mux_1754_nl = MUX_s_1_2_2(nor_940_nl, nor_941_nl, fsm_output[7]);
  assign mux_1757_nl = MUX_s_1_2_2(mux_1756_nl, mux_1754_nl, fsm_output[6]);
  assign mux_1761_nl = MUX_s_1_2_2(nor_937_nl, mux_1757_nl, fsm_output[5]);
  assign or_1593_nl = (COMP_LOOP_acc_1_cse_sva[3:0]!=4'b1001) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[0]) | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[1])
      | (~ (fsm_output[10]));
  assign or_1591_nl = (z_out_7[4:1]!=4'b1001) | (fsm_output[3]) | (fsm_output[9])
      | not_tmp_260;
  assign mux_1750_nl = MUX_s_1_2_2(or_1591_nl, or_1600_cse, fsm_output[0]);
  assign mux_1751_nl = MUX_s_1_2_2(or_1593_nl, mux_1750_nl, fsm_output[8]);
  assign or_1588_nl = (fsm_output[8]) | (fsm_output[0]) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (fsm_output[3]) | (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1001) | (fsm_output[9])
      | (~ (fsm_output[1])) | (fsm_output[10]);
  assign mux_1752_nl = MUX_s_1_2_2(mux_1751_nl, or_1588_nl, fsm_output[7]);
  assign nor_942_nl = ~((fsm_output[6]) | mux_1752_nl);
  assign nor_943_nl = ~((~ (fsm_output[0])) | (z_out_7[4:1]!=4'b1001) | (~ (fsm_output[3]))
      | (fsm_output[9]) | (~ (fsm_output[1])) | (fsm_output[10]));
  assign nor_944_nl = ~((COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b1001) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (~ (fsm_output[1])) | (fsm_output[10]));
  assign nor_945_nl = ~((COMP_LOOP_acc_20_psp_sva[2:0]!=3'b100) | (~ (VEC_LOOP_j_sva_11_0[0]))
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[3]) | (fsm_output[9])
      | not_tmp_260);
  assign mux_1747_nl = MUX_s_1_2_2(nor_944_nl, nor_945_nl, fsm_output[0]);
  assign mux_1748_nl = MUX_s_1_2_2(nor_943_nl, mux_1747_nl, fsm_output[8]);
  assign and_626_nl = (fsm_output[7]) & mux_1748_nl;
  assign nor_946_nl = ~((fsm_output[8:7]!=2'b01) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[0]) | (fsm_output[3]) | (COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b1001)
      | (~ (fsm_output[9])) | (fsm_output[1]) | (fsm_output[10]));
  assign mux_1749_nl = MUX_s_1_2_2(and_626_nl, nor_946_nl, fsm_output[6]);
  assign mux_1753_nl = MUX_s_1_2_2(nor_942_nl, mux_1749_nl, fsm_output[5]);
  assign mux_1762_nl = MUX_s_1_2_2(mux_1761_nl, mux_1753_nl, fsm_output[2]);
  assign vec_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_1776_nl,
      mux_1762_nl, fsm_output[4]);
  assign or_1689_nl = (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b101) | (fsm_output[0]) |
      (VEC_LOOP_j_sva_11_0[0]) | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[9]))
      | (fsm_output[8]) | (~ (fsm_output[10]));
  assign mux_1813_nl = MUX_s_1_2_2(or_1689_nl, or_622_cse, fsm_output[5]);
  assign mux_1814_nl = MUX_s_1_2_2(mux_1813_nl, or_621_cse, fsm_output[4]);
  assign or_1680_nl = (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b101) | (fsm_output[0]) |
      (VEC_LOOP_j_sva_11_0[0]) | (fsm_output[3]) | (~ (fsm_output[6])) | (~ (fsm_output[9]))
      | (fsm_output[8]) | (fsm_output[10]);
  assign mux_1810_nl = MUX_s_1_2_2(or_617_cse, or_1680_nl, fsm_output[5]);
  assign mux_1811_nl = MUX_s_1_2_2(mux_1810_nl, mux_tmp_1788, fsm_output[4]);
  assign mux_1815_nl = MUX_s_1_2_2(mux_1814_nl, mux_1811_nl, fsm_output[7]);
  assign mux_1809_nl = MUX_s_1_2_2(mux_tmp_1787, mux_1088_cse, fsm_output[7]);
  assign mux_1816_nl = MUX_s_1_2_2(mux_1815_nl, mux_1809_nl, fsm_output[2]);
  assign or_1670_nl = (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b1010) | (~ (fsm_output[0]))
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (~ (fsm_output[9])) | (fsm_output[8])
      | (fsm_output[10]);
  assign mux_1802_nl = MUX_s_1_2_2(or_607_cse, or_1670_nl, fsm_output[5]);
  assign mux_1803_nl = MUX_s_1_2_2(or_609_cse, mux_1802_nl, fsm_output[4]);
  assign mux_1801_nl = MUX_s_1_2_2(mux_tmp_1782, nand_25_cse, fsm_output[4]);
  assign mux_1804_nl = MUX_s_1_2_2(mux_1803_nl, mux_1801_nl, fsm_output[7]);
  assign or_1667_nl = (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b10) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b10)
      | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[9])) | (fsm_output[8])
      | (fsm_output[10]);
  assign mux_1796_nl = MUX_s_1_2_2(or_1667_nl, or_601_cse, fsm_output[0]);
  assign mux_1797_nl = MUX_s_1_2_2(mux_1796_nl, or_tmp_1580, fsm_output[5]);
  assign mux_1798_nl = MUX_s_1_2_2(or_tmp_1583, mux_1797_nl, fsm_output[4]);
  assign or_1662_nl = (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1010) | (~ (fsm_output[0]))
      | (fsm_output[3]) | (~ (fsm_output[6])) | (fsm_output[9]) | (fsm_output[8])
      | (fsm_output[10]);
  assign mux_1794_nl = MUX_s_1_2_2(mux_1073_cse, or_1662_nl, fsm_output[5]);
  assign mux_1795_nl = MUX_s_1_2_2(mux_1794_nl, or_596_cse, fsm_output[4]);
  assign mux_1799_nl = MUX_s_1_2_2(mux_1798_nl, mux_1795_nl, fsm_output[7]);
  assign mux_1805_nl = MUX_s_1_2_2(mux_1804_nl, mux_1799_nl, fsm_output[2]);
  assign mux_1817_nl = MUX_s_1_2_2(mux_1816_nl, mux_1805_nl, fsm_output[1]);
  assign or_1659_nl = (fsm_output[5:4]!=2'b00) | (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b101)
      | (fsm_output[0]) | (VEC_LOOP_j_sva_11_0[0]) | (~ (fsm_output[3])) | (fsm_output[6])
      | (~ (fsm_output[9])) | (fsm_output[8]) | (~ (fsm_output[10]));
  assign or_1657_nl = (~ (fsm_output[5])) | (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b101)
      | (fsm_output[0]) | (VEC_LOOP_j_sva_11_0[0]) | (fsm_output[3]) | (~ (fsm_output[6]))
      | (~ (fsm_output[9])) | (fsm_output[8]) | (fsm_output[10]);
  assign mux_1789_nl = MUX_s_1_2_2(or_1657_nl, mux_tmp_1788, fsm_output[4]);
  assign mux_1790_nl = MUX_s_1_2_2(or_1659_nl, mux_1789_nl, fsm_output[7]);
  assign or_1653_nl = (fsm_output[7]) | mux_tmp_1787;
  assign mux_1791_nl = MUX_s_1_2_2(mux_1790_nl, or_1653_nl, fsm_output[2]);
  assign or_1646_nl = (fsm_output[5:4]!=2'b11) | (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b1010)
      | (~ (fsm_output[0])) | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (~ (fsm_output[9]))
      | (fsm_output[8]) | (fsm_output[10]);
  assign or_1645_nl = (fsm_output[4]) | mux_tmp_1782;
  assign mux_1783_nl = MUX_s_1_2_2(or_1646_nl, or_1645_nl, fsm_output[7]);
  assign or_1638_nl = (fsm_output[0]) | (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b10) |
      (VEC_LOOP_j_sva_11_0[1:0]!=2'b10) | (fsm_output[3]) | (fsm_output[6]) | (~
      (fsm_output[9])) | (fsm_output[8]) | (fsm_output[10]);
  assign mux_1778_nl = MUX_s_1_2_2(or_1638_nl, or_tmp_1580, fsm_output[5]);
  assign mux_1779_nl = MUX_s_1_2_2(or_tmp_1583, mux_1778_nl, fsm_output[4]);
  assign or_1635_nl = (fsm_output[5:4]!=2'b10) | (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1010)
      | (~ (fsm_output[0])) | (fsm_output[3]) | (~ (fsm_output[6])) | (fsm_output[9])
      | (fsm_output[8]) | (fsm_output[10]);
  assign mux_1780_nl = MUX_s_1_2_2(mux_1779_nl, or_1635_nl, fsm_output[7]);
  assign mux_1784_nl = MUX_s_1_2_2(mux_1783_nl, mux_1780_nl, fsm_output[2]);
  assign mux_1792_nl = MUX_s_1_2_2(mux_1791_nl, mux_1784_nl, fsm_output[1]);
  assign or_1634_nl = (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b1010);
  assign mux_1818_nl = MUX_s_1_2_2(mux_1817_nl, mux_1792_nl, or_1634_nl);
  assign vec_rsc_0_10_i_wea_d_pff = ~ mux_1818_nl;
  assign nor_900_cse = ~((z_out_7[4:1]!=4'b1010) | (fsm_output[3]) | (~ (fsm_output[9]))
      | (~ (fsm_output[1])) | (fsm_output[10]));
  assign or_1707_cse = (z_out_7[4:1]!=4'b1010) | (~ (fsm_output[3])) | (~ (fsm_output[9]))
      | (fsm_output[1]) | (fsm_output[10]);
  assign nor_899_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b1010) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[0]) | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[1])
      | (~ (fsm_output[10])));
  assign nor_901_nl = ~((~ (fsm_output[3])) | (z_out_7[4:1]!=4'b1010) | (fsm_output[9])
      | (fsm_output[1]) | (fsm_output[10]));
  assign mux_1845_nl = MUX_s_1_2_2(nor_900_cse, nor_901_nl, fsm_output[0]);
  assign mux_1846_nl = MUX_s_1_2_2(nor_899_nl, mux_1845_nl, fsm_output[8]);
  assign and_621_nl = nor_223_cse & mux_1846_nl;
  assign or_1735_nl = (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b1010) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (~ (fsm_output[1])) | (fsm_output[10]);
  assign or_1734_nl = (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b101) | (VEC_LOOP_j_sva_11_0[0])
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[3]) | (fsm_output[9])
      | not_tmp_260;
  assign mux_1843_nl = MUX_s_1_2_2(or_1735_nl, or_1734_nl, fsm_output[0]);
  assign nor_902_nl = ~((fsm_output[8:7]!=2'b00) | mux_1843_nl);
  assign nor_903_nl = ~((~ (fsm_output[8])) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b1010) | (fsm_output[0]) | (fsm_output[3])
      | (fsm_output[9]) | (fsm_output[1]) | (fsm_output[10]));
  assign nor_904_nl = ~((~ (fsm_output[8])) | (fsm_output[0]) | (z_out_7[4:1]!=4'b1010)
      | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[1]) | (~ (fsm_output[10])));
  assign mux_1842_nl = MUX_s_1_2_2(nor_903_nl, nor_904_nl, fsm_output[7]);
  assign mux_1844_nl = MUX_s_1_2_2(nor_902_nl, mux_1842_nl, fsm_output[6]);
  assign mux_1847_nl = MUX_s_1_2_2(and_621_nl, mux_1844_nl, fsm_output[5]);
  assign nor_905_nl = ~((~ (fsm_output[7])) | (fsm_output[8]) | (~ (fsm_output[0]))
      | (VEC_LOOP_j_sva_11_0[0]) | (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b101) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (~ (fsm_output[1])) | (fsm_output[10]));
  assign or_1726_nl = (z_out_7[4:1]!=4'b1010) | (~ (fsm_output[3])) | (fsm_output[9])
      | (fsm_output[1]) | (~ (fsm_output[10]));
  assign or_1724_nl = (fsm_output[3]) | (z_out_7[4:1]!=4'b1010) | (~ (fsm_output[9]))
      | (fsm_output[1]) | (~ (fsm_output[10]));
  assign mux_1838_nl = MUX_s_1_2_2(or_1726_nl, or_1724_nl, fsm_output[0]);
  assign nor_906_nl = ~((fsm_output[8]) | mux_1838_nl);
  assign nor_907_nl = ~((COMP_LOOP_acc_13_psp_sva[1:0]!=2'b10) | (~ (fsm_output[8]))
      | (~ (fsm_output[0])) | (VEC_LOOP_j_sva_11_0[0]) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (~ (VEC_LOOP_j_sva_11_0[1])) | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[1])
      | (fsm_output[10]));
  assign mux_1839_nl = MUX_s_1_2_2(nor_906_nl, nor_907_nl, fsm_output[7]);
  assign mux_1840_nl = MUX_s_1_2_2(nor_905_nl, mux_1839_nl, fsm_output[6]);
  assign nor_908_nl = ~((fsm_output[8:7]!=2'b10) | (z_out_7[4:1]!=4'b1010) | (fsm_output[0])
      | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[1]) | (fsm_output[10]));
  assign nor_909_nl = ~((COMP_LOOP_acc_19_psp_sva[1:0]!=2'b10) | (~ (fsm_output[0]))
      | (VEC_LOOP_j_sva_11_0[0]) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (~
      (VEC_LOOP_j_sva_11_0[1])) | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[1])
      | (~ (fsm_output[10])));
  assign nor_910_nl = ~((z_out_7[4:1]!=4'b1010) | (~ (fsm_output[3])) | (fsm_output[9])
      | (~ (fsm_output[1])) | (fsm_output[10]));
  assign mux_1835_nl = MUX_s_1_2_2(nor_910_nl, nor_900_cse, fsm_output[0]);
  assign mux_1836_nl = MUX_s_1_2_2(nor_909_nl, mux_1835_nl, fsm_output[8]);
  assign and_622_nl = (fsm_output[7]) & mux_1836_nl;
  assign mux_1837_nl = MUX_s_1_2_2(nor_908_nl, and_622_nl, fsm_output[6]);
  assign mux_1841_nl = MUX_s_1_2_2(mux_1840_nl, mux_1837_nl, fsm_output[5]);
  assign mux_1848_nl = MUX_s_1_2_2(mux_1847_nl, mux_1841_nl, fsm_output[2]);
  assign or_1715_nl = (z_out_7[4:1]!=4'b1010) | (~ (fsm_output[3])) | (fsm_output[9])
      | (~ (fsm_output[1])) | (fsm_output[10]);
  assign or_1714_nl = (z_out_7[4:1]!=4'b1010) | (fsm_output[3]) | (~ (fsm_output[9]))
      | (~ (fsm_output[1])) | (fsm_output[10]);
  assign mux_1831_nl = MUX_s_1_2_2(or_1715_nl, or_1714_nl, fsm_output[0]);
  assign or_1713_nl = (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b1010) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (fsm_output[3]) | (fsm_output[9]) | not_tmp_260;
  assign or_1711_nl = (~ (COMP_LOOP_acc_16_psp_sva[0])) | (VEC_LOOP_j_sva_11_0[2])
      | (VEC_LOOP_j_sva_11_0[0]) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (~
      (VEC_LOOP_j_sva_11_0[1])) | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[1])
      | (fsm_output[10]);
  assign mux_1830_nl = MUX_s_1_2_2(or_1713_nl, or_1711_nl, fsm_output[0]);
  assign mux_1832_nl = MUX_s_1_2_2(mux_1831_nl, mux_1830_nl, fsm_output[8]);
  assign nor_912_nl = ~((fsm_output[7:6]!=2'b01) | mux_1832_nl);
  assign nor_913_nl = ~((fsm_output[8]) | (~ (VEC_LOOP_j_sva_11_0[3])) | (~ (fsm_output[0]))
      | (VEC_LOOP_j_sva_11_0[2:0]!=3'b010) | (fsm_output[3]) | (fsm_output[9]) |
      (fsm_output[1]) | (fsm_output[10]));
  assign or_1706_nl = (z_out_7[4:1]!=4'b1010) | (fsm_output[3]) | (fsm_output[9])
      | (fsm_output[1]) | (~ (fsm_output[10]));
  assign mux_1827_nl = MUX_s_1_2_2(or_1707_cse, or_1706_nl, fsm_output[0]);
  assign nor_914_nl = ~((fsm_output[8]) | mux_1827_nl);
  assign mux_1828_nl = MUX_s_1_2_2(nor_913_nl, nor_914_nl, fsm_output[7]);
  assign nor_915_nl = ~((~ (fsm_output[8])) | (~ (fsm_output[0])) | (~ (fsm_output[3]))
      | (z_out_7[4:1]!=4'b1010) | (fsm_output[9]) | not_tmp_260);
  assign nor_916_nl = ~((fsm_output[8]) | (~ (fsm_output[0])) | (VEC_LOOP_j_sva_11_0[0])
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b101)
      | (~ (fsm_output[3])) | (fsm_output[9]) | (~ (fsm_output[1])) | (fsm_output[10]));
  assign mux_1826_nl = MUX_s_1_2_2(nor_915_nl, nor_916_nl, fsm_output[7]);
  assign mux_1829_nl = MUX_s_1_2_2(mux_1828_nl, mux_1826_nl, fsm_output[6]);
  assign mux_1833_nl = MUX_s_1_2_2(nor_912_nl, mux_1829_nl, fsm_output[5]);
  assign or_1700_nl = (COMP_LOOP_acc_1_cse_sva[3:0]!=4'b1010) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[0]) | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[1])
      | (~ (fsm_output[10]));
  assign or_1698_nl = (z_out_7[4:1]!=4'b1010) | (fsm_output[3]) | (fsm_output[9])
      | not_tmp_260;
  assign mux_1822_nl = MUX_s_1_2_2(or_1698_nl, or_1707_cse, fsm_output[0]);
  assign mux_1823_nl = MUX_s_1_2_2(or_1700_nl, mux_1822_nl, fsm_output[8]);
  assign or_1695_nl = (fsm_output[8]) | (fsm_output[0]) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (fsm_output[3]) | (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1010) | (fsm_output[9])
      | (~ (fsm_output[1])) | (fsm_output[10]);
  assign mux_1824_nl = MUX_s_1_2_2(mux_1823_nl, or_1695_nl, fsm_output[7]);
  assign nor_917_nl = ~((fsm_output[6]) | mux_1824_nl);
  assign nor_918_nl = ~((~ (fsm_output[0])) | (z_out_7[4:1]!=4'b1010) | (~ (fsm_output[3]))
      | (fsm_output[9]) | (~ (fsm_output[1])) | (fsm_output[10]));
  assign nor_919_nl = ~((COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b1010) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (~ (fsm_output[1])) | (fsm_output[10]));
  assign nor_920_nl = ~((COMP_LOOP_acc_20_psp_sva[2:0]!=3'b101) | (VEC_LOOP_j_sva_11_0[0])
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[3]) | (fsm_output[9])
      | not_tmp_260);
  assign mux_1819_nl = MUX_s_1_2_2(nor_919_nl, nor_920_nl, fsm_output[0]);
  assign mux_1820_nl = MUX_s_1_2_2(nor_918_nl, mux_1819_nl, fsm_output[8]);
  assign and_623_nl = (fsm_output[7]) & mux_1820_nl;
  assign nor_921_nl = ~((fsm_output[8:7]!=2'b01) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[0]) | (fsm_output[3]) | (COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b1010)
      | (~ (fsm_output[9])) | (fsm_output[1]) | (fsm_output[10]));
  assign mux_1821_nl = MUX_s_1_2_2(and_623_nl, nor_921_nl, fsm_output[6]);
  assign mux_1825_nl = MUX_s_1_2_2(nor_917_nl, mux_1821_nl, fsm_output[5]);
  assign mux_1834_nl = MUX_s_1_2_2(mux_1833_nl, mux_1825_nl, fsm_output[2]);
  assign vec_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_1848_nl,
      mux_1834_nl, fsm_output[4]);
  assign or_1795_nl = (fsm_output[5:4]!=2'b00) | (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b101)
      | (fsm_output[0]) | (~ (VEC_LOOP_j_sva_11_0[0])) | (~ (fsm_output[3])) | (fsm_output[6])
      | (~ (fsm_output[9])) | (fsm_output[8]) | (~ (fsm_output[10]));
  assign or_1793_nl = (~ (fsm_output[5])) | (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b101)
      | (fsm_output[0]) | (~ (VEC_LOOP_j_sva_11_0[0])) | (fsm_output[3]) | (~ (fsm_output[6]))
      | (~ (fsm_output[9])) | (fsm_output[8]) | (fsm_output[10]);
  assign mux_1886_nl = MUX_s_1_2_2(or_1793_nl, mux_tmp_1872, fsm_output[4]);
  assign mux_1887_nl = MUX_s_1_2_2(or_1795_nl, mux_1886_nl, fsm_output[7]);
  assign or_1792_nl = (fsm_output[7]) | mux_tmp_1870;
  assign mux_1888_nl = MUX_s_1_2_2(mux_1887_nl, or_1792_nl, fsm_output[2]);
  assign nand_319_nl = ~((fsm_output[5:4]==2'b11) & (COMP_LOOP_acc_1_cse_6_sva[3:0]==4'b1011)
      & (fsm_output[0]) & (fsm_output[3]) & (fsm_output[6]) & (fsm_output[9]) & (~
      (fsm_output[8])) & (~ (fsm_output[10])));
  assign or_1790_nl = (fsm_output[4]) | mux_tmp_1859;
  assign mux_1884_nl = MUX_s_1_2_2(nand_319_nl, or_1790_nl, fsm_output[7]);
  assign or_1789_nl = (fsm_output[0]) | (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b10) |
      (VEC_LOOP_j_sva_11_0[1:0]!=2'b11) | (fsm_output[3]) | (fsm_output[6]) | (~
      (fsm_output[9])) | (fsm_output[8]) | (fsm_output[10]);
  assign mux_1881_nl = MUX_s_1_2_2(or_1789_nl, or_tmp_1691, fsm_output[5]);
  assign mux_1882_nl = MUX_s_1_2_2(or_tmp_1695, mux_1881_nl, fsm_output[4]);
  assign or_1788_nl = (fsm_output[5:4]!=2'b10) | (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1011)
      | (~ (fsm_output[0])) | (fsm_output[3]) | (~ (fsm_output[6])) | (fsm_output[9])
      | (fsm_output[8]) | (fsm_output[10]);
  assign mux_1883_nl = MUX_s_1_2_2(mux_1882_nl, or_1788_nl, fsm_output[7]);
  assign mux_1885_nl = MUX_s_1_2_2(mux_1884_nl, mux_1883_nl, fsm_output[2]);
  assign mux_1889_nl = MUX_s_1_2_2(mux_1888_nl, mux_1885_nl, fsm_output[1]);
  assign or_1787_nl = (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b101) | (fsm_output[0]) |
      (~ (VEC_LOOP_j_sva_11_0[0])) | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[9]))
      | (fsm_output[8]) | (~ (fsm_output[10]));
  assign mux_1876_nl = MUX_s_1_2_2(or_1787_nl, or_622_cse, fsm_output[5]);
  assign mux_1877_nl = MUX_s_1_2_2(mux_1876_nl, or_621_cse, fsm_output[4]);
  assign or_1778_nl = (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b101) | (fsm_output[0]) |
      (~ (VEC_LOOP_j_sva_11_0[0])) | (fsm_output[3]) | (~ (fsm_output[6])) | (~ (fsm_output[9]))
      | (fsm_output[8]) | (fsm_output[10]);
  assign mux_1873_nl = MUX_s_1_2_2(or_617_cse, or_1778_nl, fsm_output[5]);
  assign mux_1874_nl = MUX_s_1_2_2(mux_1873_nl, mux_tmp_1872, fsm_output[4]);
  assign mux_1878_nl = MUX_s_1_2_2(mux_1877_nl, mux_1874_nl, fsm_output[7]);
  assign mux_1871_nl = MUX_s_1_2_2(mux_tmp_1870, mux_1088_cse, fsm_output[7]);
  assign mux_1879_nl = MUX_s_1_2_2(mux_1878_nl, mux_1871_nl, fsm_output[2]);
  assign nand_321_nl = ~((COMP_LOOP_acc_1_cse_6_sva[3:0]==4'b1011) & (fsm_output[0])
      & (fsm_output[3]) & (fsm_output[6]) & (fsm_output[9]) & (~ (fsm_output[8]))
      & (~ (fsm_output[10])));
  assign mux_1861_nl = MUX_s_1_2_2(or_607_cse, nand_321_nl, fsm_output[5]);
  assign mux_1862_nl = MUX_s_1_2_2(or_609_cse, mux_1861_nl, fsm_output[4]);
  assign mux_1860_nl = MUX_s_1_2_2(mux_tmp_1859, nand_25_cse, fsm_output[4]);
  assign mux_1863_nl = MUX_s_1_2_2(mux_1862_nl, mux_1860_nl, fsm_output[7]);
  assign or_1750_nl = (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b10) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b11)
      | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[9])) | (fsm_output[8])
      | (fsm_output[10]);
  assign mux_1853_nl = MUX_s_1_2_2(or_1750_nl, or_601_cse, fsm_output[0]);
  assign mux_1854_nl = MUX_s_1_2_2(mux_1853_nl, or_tmp_1691, fsm_output[5]);
  assign mux_1855_nl = MUX_s_1_2_2(or_tmp_1695, mux_1854_nl, fsm_output[4]);
  assign or_1743_nl = (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1011) | (~ (fsm_output[0]))
      | (fsm_output[3]) | (~ (fsm_output[6])) | (fsm_output[9]) | (fsm_output[8])
      | (fsm_output[10]);
  assign mux_1851_nl = MUX_s_1_2_2(mux_1073_cse, or_1743_nl, fsm_output[5]);
  assign mux_1852_nl = MUX_s_1_2_2(mux_1851_nl, or_596_cse, fsm_output[4]);
  assign mux_1856_nl = MUX_s_1_2_2(mux_1855_nl, mux_1852_nl, fsm_output[7]);
  assign mux_1864_nl = MUX_s_1_2_2(mux_1863_nl, mux_1856_nl, fsm_output[2]);
  assign mux_1880_nl = MUX_s_1_2_2(mux_1879_nl, mux_1864_nl, fsm_output[1]);
  assign and_620_nl = (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]==4'b1011);
  assign mux_1890_nl = MUX_s_1_2_2(mux_1889_nl, mux_1880_nl, and_620_nl);
  assign vec_rsc_0_11_i_wea_d_pff = ~ mux_1890_nl;
  assign nor_877_cse = ~((z_out_7[4:1]!=4'b1011) | (fsm_output[3]) | (~ (fsm_output[9]))
      | (~ (fsm_output[1])) | (fsm_output[10]));
  assign or_1813_cse = (z_out_7[4:1]!=4'b1011) | (~ (fsm_output[3])) | (~ (fsm_output[9]))
      | (fsm_output[1]) | (fsm_output[10]);
  assign nor_876_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b1011) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[0]) | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[1])
      | (~ (fsm_output[10])));
  assign nor_878_nl = ~((~ (fsm_output[3])) | (z_out_7[4:1]!=4'b1011) | (fsm_output[9])
      | (fsm_output[1]) | (fsm_output[10]));
  assign mux_1917_nl = MUX_s_1_2_2(nor_877_cse, nor_878_nl, fsm_output[0]);
  assign mux_1918_nl = MUX_s_1_2_2(nor_876_nl, mux_1917_nl, fsm_output[8]);
  assign and_615_nl = nor_223_cse & mux_1918_nl;
  assign nand_316_nl = ~((COMP_LOOP_acc_1_cse_6_sva[3:0]==4'b1011) & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm
      & (fsm_output[3]) & (fsm_output[9]) & (fsm_output[1]) & (~ (fsm_output[10])));
  assign or_1840_nl = (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b101) | (~ (VEC_LOOP_j_sva_11_0[0]))
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[3]) | (fsm_output[9])
      | not_tmp_260;
  assign mux_1915_nl = MUX_s_1_2_2(nand_316_nl, or_1840_nl, fsm_output[0]);
  assign nor_879_nl = ~((fsm_output[8:7]!=2'b00) | mux_1915_nl);
  assign nor_880_nl = ~((~ (fsm_output[8])) | (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b1011)
      | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) | (fsm_output[0]) | (fsm_output[3])
      | (fsm_output[9]) | (fsm_output[1]) | (fsm_output[10]));
  assign nor_881_nl = ~((~ (fsm_output[8])) | (fsm_output[0]) | (z_out_7[4:1]!=4'b1011)
      | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[1]) | (~ (fsm_output[10])));
  assign mux_1914_nl = MUX_s_1_2_2(nor_880_nl, nor_881_nl, fsm_output[7]);
  assign mux_1916_nl = MUX_s_1_2_2(nor_879_nl, mux_1914_nl, fsm_output[6]);
  assign mux_1919_nl = MUX_s_1_2_2(and_615_nl, mux_1916_nl, fsm_output[5]);
  assign and_616_nl = (fsm_output[7]) & (~ (fsm_output[8])) & (fsm_output[0]) & (VEC_LOOP_j_sva_11_0[0])
      & (COMP_LOOP_acc_14_psp_sva[2:0]==3'b101) & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm
      & (fsm_output[3]) & (fsm_output[9]) & (fsm_output[1]) & (~ (fsm_output[10]));
  assign or_1832_nl = (z_out_7[4:1]!=4'b1011) | (~ (fsm_output[3])) | (fsm_output[9])
      | (fsm_output[1]) | (~ (fsm_output[10]));
  assign or_1830_nl = (fsm_output[3]) | (z_out_7[4:1]!=4'b1011) | (~ (fsm_output[9]))
      | (fsm_output[1]) | (~ (fsm_output[10]));
  assign mux_1910_nl = MUX_s_1_2_2(or_1832_nl, or_1830_nl, fsm_output[0]);
  assign nor_882_nl = ~((fsm_output[8]) | mux_1910_nl);
  assign nor_883_nl = ~((COMP_LOOP_acc_13_psp_sva[1:0]!=2'b10) | (~ (fsm_output[8]))
      | (~ (fsm_output[0])) | (~ (VEC_LOOP_j_sva_11_0[0])) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (~ (VEC_LOOP_j_sva_11_0[1])) | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[1])
      | (fsm_output[10]));
  assign mux_1911_nl = MUX_s_1_2_2(nor_882_nl, nor_883_nl, fsm_output[7]);
  assign mux_1912_nl = MUX_s_1_2_2(and_616_nl, mux_1911_nl, fsm_output[6]);
  assign nor_884_nl = ~((fsm_output[8:7]!=2'b10) | (z_out_7[4:1]!=4'b1011) | (fsm_output[0])
      | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[1]) | (fsm_output[10]));
  assign and_827_nl = (COMP_LOOP_acc_19_psp_sva[1:0]==2'b10) & (fsm_output[0]) &
      (VEC_LOOP_j_sva_11_0[0]) & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm & (VEC_LOOP_j_sva_11_0[1])
      & (fsm_output[3]) & (~ (fsm_output[9])) & (~ (fsm_output[1])) & (fsm_output[10]);
  assign nor_886_nl = ~((z_out_7[4:1]!=4'b1011) | (~ (fsm_output[3])) | (fsm_output[9])
      | (~ (fsm_output[1])) | (fsm_output[10]));
  assign mux_1907_nl = MUX_s_1_2_2(nor_886_nl, nor_877_cse, fsm_output[0]);
  assign mux_1908_nl = MUX_s_1_2_2(and_827_nl, mux_1907_nl, fsm_output[8]);
  assign and_617_nl = (fsm_output[7]) & mux_1908_nl;
  assign mux_1909_nl = MUX_s_1_2_2(nor_884_nl, and_617_nl, fsm_output[6]);
  assign mux_1913_nl = MUX_s_1_2_2(mux_1912_nl, mux_1909_nl, fsm_output[5]);
  assign mux_1920_nl = MUX_s_1_2_2(mux_1919_nl, mux_1913_nl, fsm_output[2]);
  assign or_1821_nl = (z_out_7[4:1]!=4'b1011) | (~ (fsm_output[3])) | (fsm_output[9])
      | (~ (fsm_output[1])) | (fsm_output[10]);
  assign or_1820_nl = (z_out_7[4:1]!=4'b1011) | (fsm_output[3]) | (~ (fsm_output[9]))
      | (~ (fsm_output[1])) | (fsm_output[10]);
  assign mux_1903_nl = MUX_s_1_2_2(or_1821_nl, or_1820_nl, fsm_output[0]);
  assign or_1819_nl = (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b1011) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (fsm_output[3]) | (fsm_output[9]) | not_tmp_260;
  assign or_1817_nl = (~ (COMP_LOOP_acc_16_psp_sva[0])) | (VEC_LOOP_j_sva_11_0[2])
      | (~ (VEC_LOOP_j_sva_11_0[0])) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) |
      (~ (VEC_LOOP_j_sva_11_0[1])) | (~ (fsm_output[3])) | (~ (fsm_output[9])) |
      (fsm_output[1]) | (fsm_output[10]);
  assign mux_1902_nl = MUX_s_1_2_2(or_1819_nl, or_1817_nl, fsm_output[0]);
  assign mux_1904_nl = MUX_s_1_2_2(mux_1903_nl, mux_1902_nl, fsm_output[8]);
  assign nor_888_nl = ~((fsm_output[7:6]!=2'b01) | mux_1904_nl);
  assign nor_889_nl = ~((fsm_output[8]) | (~ (VEC_LOOP_j_sva_11_0[3])) | (~ (fsm_output[0]))
      | (VEC_LOOP_j_sva_11_0[2:0]!=3'b011) | (fsm_output[3]) | (fsm_output[9]) |
      (fsm_output[1]) | (fsm_output[10]));
  assign or_1812_nl = (z_out_7[4:1]!=4'b1011) | (fsm_output[3]) | (fsm_output[9])
      | (fsm_output[1]) | (~ (fsm_output[10]));
  assign mux_1899_nl = MUX_s_1_2_2(or_1813_cse, or_1812_nl, fsm_output[0]);
  assign nor_890_nl = ~((fsm_output[8]) | mux_1899_nl);
  assign mux_1900_nl = MUX_s_1_2_2(nor_889_nl, nor_890_nl, fsm_output[7]);
  assign nor_891_nl = ~((~((fsm_output[8]) & (fsm_output[0]) & (fsm_output[3]) &
      (z_out_7[4:1]==4'b1011) & (~ (fsm_output[9])))) | not_tmp_260);
  assign nor_892_nl = ~((fsm_output[8]) | (~ (fsm_output[0])) | (~ (VEC_LOOP_j_sva_11_0[0]))
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b101)
      | (~ (fsm_output[3])) | (fsm_output[9]) | (~ (fsm_output[1])) | (fsm_output[10]));
  assign mux_1898_nl = MUX_s_1_2_2(nor_891_nl, nor_892_nl, fsm_output[7]);
  assign mux_1901_nl = MUX_s_1_2_2(mux_1900_nl, mux_1898_nl, fsm_output[6]);
  assign mux_1905_nl = MUX_s_1_2_2(nor_888_nl, mux_1901_nl, fsm_output[5]);
  assign nand_415_nl = ~((COMP_LOOP_acc_1_cse_sva[3:0]==4'b1011) & COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm
      & (~ (fsm_output[0])) & (fsm_output[3]) & (fsm_output[9]) & (~ (fsm_output[1]))
      & (fsm_output[10]));
  assign or_1804_nl = (z_out_7[4:1]!=4'b1011) | (fsm_output[3]) | (fsm_output[9])
      | not_tmp_260;
  assign mux_1894_nl = MUX_s_1_2_2(or_1804_nl, or_1813_cse, fsm_output[0]);
  assign mux_1895_nl = MUX_s_1_2_2(nand_415_nl, mux_1894_nl, fsm_output[8]);
  assign or_1801_nl = (fsm_output[8]) | (fsm_output[0]) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (fsm_output[3]) | (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1011) | (fsm_output[9])
      | (~ (fsm_output[1])) | (fsm_output[10]);
  assign mux_1896_nl = MUX_s_1_2_2(mux_1895_nl, or_1801_nl, fsm_output[7]);
  assign nor_893_nl = ~((fsm_output[6]) | mux_1896_nl);
  assign nor_894_nl = ~((~ (fsm_output[0])) | (z_out_7[4:1]!=4'b1011) | (~ (fsm_output[3]))
      | (fsm_output[9]) | (~ (fsm_output[1])) | (fsm_output[10]));
  assign and_619_nl = (COMP_LOOP_acc_1_cse_10_sva[3:0]==4'b1011) & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm
      & (fsm_output[3]) & (fsm_output[9]) & (fsm_output[1]) & (~ (fsm_output[10]));
  assign nor_895_nl = ~((COMP_LOOP_acc_20_psp_sva[2:0]!=3'b101) | (~ (VEC_LOOP_j_sva_11_0[0]))
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[3]) | (fsm_output[9])
      | not_tmp_260);
  assign mux_1891_nl = MUX_s_1_2_2(and_619_nl, nor_895_nl, fsm_output[0]);
  assign mux_1892_nl = MUX_s_1_2_2(nor_894_nl, mux_1891_nl, fsm_output[8]);
  assign and_618_nl = (fsm_output[7]) & mux_1892_nl;
  assign nor_896_nl = ~((fsm_output[8:7]!=2'b01) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[0]) | (fsm_output[3]) | (COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b1011)
      | (~ (fsm_output[9])) | (fsm_output[1]) | (fsm_output[10]));
  assign mux_1893_nl = MUX_s_1_2_2(and_618_nl, nor_896_nl, fsm_output[6]);
  assign mux_1897_nl = MUX_s_1_2_2(nor_893_nl, mux_1893_nl, fsm_output[5]);
  assign mux_1906_nl = MUX_s_1_2_2(mux_1905_nl, mux_1897_nl, fsm_output[2]);
  assign vec_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_1920_nl,
      mux_1906_nl, fsm_output[4]);
  assign or_1905_nl = (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b110) | (fsm_output[0]) |
      (VEC_LOOP_j_sva_11_0[0]) | (fsm_output[4]) | (~ (fsm_output[9])) | (~ (fsm_output[3]))
      | (fsm_output[6]) | (~ (fsm_output[10]));
  assign or_1903_nl = (~ (fsm_output[0])) | (fsm_output[4]) | (~ (fsm_output[9]))
      | (~ (fsm_output[3])) | (fsm_output[6]) | (fsm_output[10]);
  assign mux_1958_nl = MUX_s_1_2_2(or_1905_nl, or_1903_nl, fsm_output[5]);
  assign nand_311_nl = ~((fsm_output[4]) & (fsm_output[9]) & (fsm_output[3]) & (fsm_output[6])
      & (~ (fsm_output[10])));
  assign or_1900_nl = (~ (fsm_output[4])) | (fsm_output[9]) | (fsm_output[3]) | not_tmp_378;
  assign mux_1957_nl = MUX_s_1_2_2(nand_311_nl, or_1900_nl, fsm_output[0]);
  assign or_1902_nl = (fsm_output[5]) | mux_1957_nl;
  assign mux_1959_nl = MUX_s_1_2_2(mux_1958_nl, or_1902_nl, fsm_output[8]);
  assign or_1898_nl = (fsm_output[4]) | (~ (fsm_output[9])) | (fsm_output[3]) | (fsm_output[6])
      | (~ (fsm_output[10]));
  assign or_1896_nl = (COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b1100) | (~ (fsm_output[4]))
      | (fsm_output[9]) | not_tmp_381;
  assign mux_1954_nl = MUX_s_1_2_2(or_1898_nl, or_1896_nl, fsm_output[0]);
  assign mux_1955_nl = MUX_s_1_2_2(mux_1954_nl, or_tmp_1812, fsm_output[5]);
  assign mux_1956_nl = MUX_s_1_2_2(mux_1955_nl, or_tmp_1811, fsm_output[8]);
  assign mux_1960_nl = MUX_s_1_2_2(mux_1959_nl, mux_1956_nl, fsm_output[7]);
  assign nand_437_nl = ~((fsm_output[0]) & (fsm_output[4]) & (fsm_output[9]) & (fsm_output[3])
      & (~ (fsm_output[6])) & (fsm_output[10]));
  assign or_1891_nl = (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b1100) | (~ (fsm_output[4]))
      | (~ (fsm_output[9])) | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[10]);
  assign mux_1951_nl = MUX_s_1_2_2(or_tmp_1821, or_1891_nl, fsm_output[0]);
  assign mux_1952_nl = MUX_s_1_2_2(nand_437_nl, mux_1951_nl, fsm_output[5]);
  assign or_1894_nl = (fsm_output[8]) | mux_1952_nl;
  assign or_1890_nl = (~ (VEC_LOOP_j_sva_11_0[3])) | (fsm_output[0]) | (VEC_LOOP_j_sva_11_0[2:0]!=3'b100)
      | (fsm_output[4]) | (fsm_output[9]) | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[10]);
  assign or_1889_nl = (~ (fsm_output[4])) | (fsm_output[9]) | (~ (fsm_output[3]))
      | (~ (fsm_output[6])) | (fsm_output[10]);
  assign or_1888_nl = (~ (fsm_output[4])) | (~ (fsm_output[9])) | (fsm_output[3])
      | (~ (fsm_output[6])) | (fsm_output[10]);
  assign mux_1948_nl = MUX_s_1_2_2(or_1889_nl, or_1888_nl, fsm_output[0]);
  assign mux_1949_nl = MUX_s_1_2_2(or_1890_nl, mux_1948_nl, fsm_output[5]);
  assign mux_1950_nl = MUX_s_1_2_2(mux_1949_nl, nand_tmp_74, fsm_output[8]);
  assign mux_1953_nl = MUX_s_1_2_2(or_1894_nl, mux_1950_nl, fsm_output[7]);
  assign mux_1961_nl = MUX_s_1_2_2(mux_1960_nl, mux_1953_nl, fsm_output[1]);
  assign or_1887_nl = (~ (fsm_output[0])) | (~ (fsm_output[4])) | (fsm_output[9])
      | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[10]);
  assign or_1886_nl = (fsm_output[0]) | (fsm_output[4]) | (fsm_output[9]) | not_tmp_381;
  assign mux_1944_nl = MUX_s_1_2_2(or_1887_nl, or_1886_nl, fsm_output[5]);
  assign or_1884_nl = (fsm_output[0]) | (fsm_output[4]) | (fsm_output[9]) | (fsm_output[3])
      | (~ (fsm_output[6])) | (fsm_output[10]);
  assign or_1883_nl = (~ (fsm_output[0])) | (~ (fsm_output[4])) | (~ (fsm_output[9]))
      | (~ (fsm_output[3])) | (fsm_output[6]) | (fsm_output[10]);
  assign mux_1943_nl = MUX_s_1_2_2(or_1884_nl, or_1883_nl, fsm_output[5]);
  assign mux_1945_nl = MUX_s_1_2_2(mux_1944_nl, mux_1943_nl, fsm_output[8]);
  assign mux_1946_nl = MUX_s_1_2_2(mux_tmp_1927, mux_1945_nl, fsm_output[7]);
  assign or_1882_nl = (~ (fsm_output[0])) | (~ (fsm_output[4])) | (fsm_output[9])
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[10]);
  assign or_1881_nl = (COMP_LOOP_acc_19_psp_sva[1:0]!=2'b11) | (fsm_output[0]) |
      (VEC_LOOP_j_sva_11_0[1:0]!=2'b00) | (~ (fsm_output[4])) | (fsm_output[9]) |
      (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[10]));
  assign mux_1940_nl = MUX_s_1_2_2(or_1882_nl, or_1881_nl, fsm_output[5]);
  assign mux_1941_nl = MUX_s_1_2_2(or_tmp_1797, mux_1940_nl, fsm_output[8]);
  assign or_1879_nl = (fsm_output[4]) | (~ (fsm_output[9])) | (~ (fsm_output[3]))
      | (fsm_output[6]) | (fsm_output[10]);
  assign mux_1937_nl = MUX_s_1_2_2(or_1879_nl, or_tmp_1821, fsm_output[0]);
  assign or_1876_nl = (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1100) | (~ (fsm_output[0]))
      | (fsm_output[4]) | (fsm_output[9]) | (fsm_output[3]) | (~ (fsm_output[6]))
      | (fsm_output[10]);
  assign mux_1938_nl = MUX_s_1_2_2(mux_1937_nl, or_1876_nl, fsm_output[5]);
  assign or_1875_nl = (~ (fsm_output[5])) | (fsm_output[0]) | (~ (fsm_output[4]))
      | (fsm_output[9]) | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[10]));
  assign mux_1939_nl = MUX_s_1_2_2(mux_1938_nl, or_1875_nl, fsm_output[8]);
  assign mux_1942_nl = MUX_s_1_2_2(mux_1941_nl, mux_1939_nl, fsm_output[7]);
  assign mux_1947_nl = MUX_s_1_2_2(mux_1946_nl, mux_1942_nl, fsm_output[1]);
  assign mux_1962_nl = MUX_s_1_2_2(mux_1961_nl, mux_1947_nl, fsm_output[2]);
  assign or_1873_nl = (fsm_output[8]) | (fsm_output[5]) | (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b110)
      | (fsm_output[0]) | (VEC_LOOP_j_sva_11_0[0]) | (fsm_output[4]) | (~ (fsm_output[9]))
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[10]));
  assign or_1871_nl = (~ (fsm_output[0])) | (COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b1100)
      | (~ (fsm_output[4])) | (fsm_output[9]) | not_tmp_381;
  assign mux_1932_nl = MUX_s_1_2_2(or_1871_nl, or_tmp_1812, fsm_output[5]);
  assign mux_1933_nl = MUX_s_1_2_2(mux_1932_nl, or_tmp_1811, fsm_output[8]);
  assign mux_1934_nl = MUX_s_1_2_2(or_1873_nl, mux_1933_nl, fsm_output[7]);
  assign or_1867_nl = (fsm_output[8]) | (~ (fsm_output[5])) | (~ (fsm_output[0]))
      | (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b1100) | (~ (fsm_output[4])) | (~ (fsm_output[9]))
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[10]);
  assign or_1866_nl = (fsm_output[5]) | (~ (VEC_LOOP_j_sva_11_0[3])) | (fsm_output[0])
      | (VEC_LOOP_j_sva_11_0[2:0]!=3'b100) | (fsm_output[4]) | (fsm_output[9]) |
      (fsm_output[3]) | (fsm_output[6]) | (fsm_output[10]);
  assign mux_1930_nl = MUX_s_1_2_2(or_1866_nl, nand_tmp_74, fsm_output[8]);
  assign mux_1931_nl = MUX_s_1_2_2(or_1867_nl, mux_1930_nl, fsm_output[7]);
  assign mux_1935_nl = MUX_s_1_2_2(mux_1934_nl, mux_1931_nl, fsm_output[1]);
  assign or_1862_nl = (fsm_output[7]) | mux_tmp_1927;
  assign or_1850_nl = (~ (fsm_output[5])) | (COMP_LOOP_acc_19_psp_sva[1:0]!=2'b11)
      | (fsm_output[0]) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b00) | (~ (fsm_output[4]))
      | (fsm_output[9]) | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[10]));
  assign mux_1923_nl = MUX_s_1_2_2(or_tmp_1797, or_1850_nl, fsm_output[8]);
  assign or_1848_nl = (fsm_output[8]) | (~ (fsm_output[5])) | (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1100)
      | (~ (fsm_output[0])) | (fsm_output[4]) | (fsm_output[9]) | (fsm_output[3])
      | (~ (fsm_output[6])) | (fsm_output[10]);
  assign mux_1924_nl = MUX_s_1_2_2(mux_1923_nl, or_1848_nl, fsm_output[7]);
  assign mux_1928_nl = MUX_s_1_2_2(or_1862_nl, mux_1924_nl, fsm_output[1]);
  assign mux_1936_nl = MUX_s_1_2_2(mux_1935_nl, mux_1928_nl, fsm_output[2]);
  assign or_1847_nl = (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b1100);
  assign mux_1963_nl = MUX_s_1_2_2(mux_1962_nl, mux_1936_nl, or_1847_nl);
  assign vec_rsc_0_12_i_wea_d_pff = ~ mux_1963_nl;
  assign nor_850_cse = ~((z_out_7[4:1]!=4'b1100) | (fsm_output[3]) | (~ (fsm_output[9]))
      | (~ (fsm_output[1])) | (fsm_output[10]));
  assign or_1923_cse = (z_out_7[4:1]!=4'b1100) | (~ (fsm_output[3])) | (~ (fsm_output[9]))
      | (fsm_output[1]) | (fsm_output[10]);
  assign nor_849_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b1100) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[0]) | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[1])
      | (~ (fsm_output[10])));
  assign nor_851_nl = ~((~ (fsm_output[3])) | (z_out_7[4:1]!=4'b1100) | (fsm_output[9])
      | (fsm_output[1]) | (fsm_output[10]));
  assign mux_1990_nl = MUX_s_1_2_2(nor_850_cse, nor_851_nl, fsm_output[0]);
  assign mux_1991_nl = MUX_s_1_2_2(nor_849_nl, mux_1990_nl, fsm_output[8]);
  assign and_612_nl = nor_223_cse & mux_1991_nl;
  assign or_1951_nl = (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b1100) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (~ (fsm_output[1])) | (fsm_output[10]);
  assign or_1950_nl = (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b110) | (VEC_LOOP_j_sva_11_0[0])
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[3]) | (fsm_output[9])
      | not_tmp_260;
  assign mux_1988_nl = MUX_s_1_2_2(or_1951_nl, or_1950_nl, fsm_output[0]);
  assign nor_852_nl = ~((fsm_output[8:7]!=2'b00) | mux_1988_nl);
  assign nor_853_nl = ~((~ (fsm_output[8])) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b1100) | (fsm_output[0]) | (fsm_output[3])
      | (fsm_output[9]) | (fsm_output[1]) | (fsm_output[10]));
  assign nor_854_nl = ~((~ (fsm_output[8])) | (fsm_output[0]) | (z_out_7[4:1]!=4'b1100)
      | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[1]) | (~ (fsm_output[10])));
  assign mux_1987_nl = MUX_s_1_2_2(nor_853_nl, nor_854_nl, fsm_output[7]);
  assign mux_1989_nl = MUX_s_1_2_2(nor_852_nl, mux_1987_nl, fsm_output[6]);
  assign mux_1992_nl = MUX_s_1_2_2(and_612_nl, mux_1989_nl, fsm_output[5]);
  assign nor_855_nl = ~((~ (fsm_output[7])) | (fsm_output[8]) | (~ (fsm_output[0]))
      | (VEC_LOOP_j_sva_11_0[0]) | (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b110) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (~ (fsm_output[1])) | (fsm_output[10]));
  assign or_1942_nl = (z_out_7[4:1]!=4'b1100) | (~ (fsm_output[3])) | (fsm_output[9])
      | (fsm_output[1]) | (~ (fsm_output[10]));
  assign or_1940_nl = (fsm_output[3]) | (z_out_7[4:1]!=4'b1100) | (~ (fsm_output[9]))
      | (fsm_output[1]) | (~ (fsm_output[10]));
  assign mux_1983_nl = MUX_s_1_2_2(or_1942_nl, or_1940_nl, fsm_output[0]);
  assign nor_856_nl = ~((fsm_output[8]) | mux_1983_nl);
  assign nor_857_nl = ~((COMP_LOOP_acc_13_psp_sva[1:0]!=2'b11) | (~ (fsm_output[8]))
      | (~ (fsm_output[0])) | (VEC_LOOP_j_sva_11_0[0]) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (VEC_LOOP_j_sva_11_0[1]) | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[1])
      | (fsm_output[10]));
  assign mux_1984_nl = MUX_s_1_2_2(nor_856_nl, nor_857_nl, fsm_output[7]);
  assign mux_1985_nl = MUX_s_1_2_2(nor_855_nl, mux_1984_nl, fsm_output[6]);
  assign nor_858_nl = ~((fsm_output[8:7]!=2'b10) | (z_out_7[4:1]!=4'b1100) | (fsm_output[0])
      | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[1]) | (fsm_output[10]));
  assign nor_859_nl = ~((COMP_LOOP_acc_19_psp_sva[1:0]!=2'b11) | (~ (fsm_output[0]))
      | (VEC_LOOP_j_sva_11_0[0]) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (VEC_LOOP_j_sva_11_0[1])
      | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[1]) | (~ (fsm_output[10])));
  assign nor_860_nl = ~((z_out_7[4:1]!=4'b1100) | (~ (fsm_output[3])) | (fsm_output[9])
      | (~ (fsm_output[1])) | (fsm_output[10]));
  assign mux_1980_nl = MUX_s_1_2_2(nor_860_nl, nor_850_cse, fsm_output[0]);
  assign mux_1981_nl = MUX_s_1_2_2(nor_859_nl, mux_1980_nl, fsm_output[8]);
  assign and_613_nl = (fsm_output[7]) & mux_1981_nl;
  assign mux_1982_nl = MUX_s_1_2_2(nor_858_nl, and_613_nl, fsm_output[6]);
  assign mux_1986_nl = MUX_s_1_2_2(mux_1985_nl, mux_1982_nl, fsm_output[5]);
  assign mux_1993_nl = MUX_s_1_2_2(mux_1992_nl, mux_1986_nl, fsm_output[2]);
  assign or_1931_nl = (z_out_7[4:1]!=4'b1100) | (~ (fsm_output[3])) | (fsm_output[9])
      | (~ (fsm_output[1])) | (fsm_output[10]);
  assign or_1930_nl = (z_out_7[4:1]!=4'b1100) | (fsm_output[3]) | (~ (fsm_output[9]))
      | (~ (fsm_output[1])) | (fsm_output[10]);
  assign mux_1976_nl = MUX_s_1_2_2(or_1931_nl, or_1930_nl, fsm_output[0]);
  assign or_1929_nl = (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b1100) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (fsm_output[3]) | (fsm_output[9]) | not_tmp_260;
  assign or_1927_nl = (~ (COMP_LOOP_acc_16_psp_sva[0])) | (~ (VEC_LOOP_j_sva_11_0[2]))
      | (VEC_LOOP_j_sva_11_0[0]) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (VEC_LOOP_j_sva_11_0[1])
      | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[1]) | (fsm_output[10]);
  assign mux_1975_nl = MUX_s_1_2_2(or_1929_nl, or_1927_nl, fsm_output[0]);
  assign mux_1977_nl = MUX_s_1_2_2(mux_1976_nl, mux_1975_nl, fsm_output[8]);
  assign nor_862_nl = ~((fsm_output[7:6]!=2'b01) | mux_1977_nl);
  assign nor_863_nl = ~((fsm_output[8]) | (~ (VEC_LOOP_j_sva_11_0[3])) | (~ (fsm_output[0]))
      | (VEC_LOOP_j_sva_11_0[2:0]!=3'b100) | (fsm_output[3]) | (fsm_output[9]) |
      (fsm_output[1]) | (fsm_output[10]));
  assign or_1922_nl = (z_out_7[4:1]!=4'b1100) | (fsm_output[3]) | (fsm_output[9])
      | (fsm_output[1]) | (~ (fsm_output[10]));
  assign mux_1972_nl = MUX_s_1_2_2(or_1923_cse, or_1922_nl, fsm_output[0]);
  assign nor_864_nl = ~((fsm_output[8]) | mux_1972_nl);
  assign mux_1973_nl = MUX_s_1_2_2(nor_863_nl, nor_864_nl, fsm_output[7]);
  assign nor_865_nl = ~((z_out_7[4:1]!=4'b1100) | (~ (fsm_output[8])) | (~ (fsm_output[0]))
      | (~ (fsm_output[3])) | (fsm_output[9]) | not_tmp_260);
  assign nor_866_nl = ~((fsm_output[8]) | (~ (fsm_output[0])) | (VEC_LOOP_j_sva_11_0[0])
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b110)
      | (~ (fsm_output[3])) | (fsm_output[9]) | (~ (fsm_output[1])) | (fsm_output[10]));
  assign mux_1971_nl = MUX_s_1_2_2(nor_865_nl, nor_866_nl, fsm_output[7]);
  assign mux_1974_nl = MUX_s_1_2_2(mux_1973_nl, mux_1971_nl, fsm_output[6]);
  assign mux_1978_nl = MUX_s_1_2_2(nor_862_nl, mux_1974_nl, fsm_output[5]);
  assign or_1916_nl = (COMP_LOOP_acc_1_cse_sva[3:0]!=4'b1100) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[0]) | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[1])
      | (~ (fsm_output[10]));
  assign or_1914_nl = (z_out_7[4:1]!=4'b1100) | (fsm_output[3]) | (fsm_output[9])
      | not_tmp_260;
  assign mux_1967_nl = MUX_s_1_2_2(or_1914_nl, or_1923_cse, fsm_output[0]);
  assign mux_1968_nl = MUX_s_1_2_2(or_1916_nl, mux_1967_nl, fsm_output[8]);
  assign or_1911_nl = (fsm_output[8]) | (fsm_output[0]) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (fsm_output[3]) | (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1100) | (fsm_output[9])
      | (~ (fsm_output[1])) | (fsm_output[10]);
  assign mux_1969_nl = MUX_s_1_2_2(mux_1968_nl, or_1911_nl, fsm_output[7]);
  assign nor_867_nl = ~((fsm_output[6]) | mux_1969_nl);
  assign nor_868_nl = ~((~ (fsm_output[0])) | (z_out_7[4:1]!=4'b1100) | (~ (fsm_output[3]))
      | (fsm_output[9]) | (~ (fsm_output[1])) | (fsm_output[10]));
  assign nor_869_nl = ~((COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b1100) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (~ (fsm_output[1])) | (fsm_output[10]));
  assign nor_870_nl = ~((COMP_LOOP_acc_20_psp_sva[2:0]!=3'b110) | (VEC_LOOP_j_sva_11_0[0])
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[3]) | (fsm_output[9])
      | not_tmp_260);
  assign mux_1964_nl = MUX_s_1_2_2(nor_869_nl, nor_870_nl, fsm_output[0]);
  assign mux_1965_nl = MUX_s_1_2_2(nor_868_nl, mux_1964_nl, fsm_output[8]);
  assign and_614_nl = (fsm_output[7]) & mux_1965_nl;
  assign nor_871_nl = ~((fsm_output[8:7]!=2'b01) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[0]) | (fsm_output[3]) | (COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b1100)
      | (~ (fsm_output[9])) | (fsm_output[1]) | (fsm_output[10]));
  assign mux_1966_nl = MUX_s_1_2_2(and_614_nl, nor_871_nl, fsm_output[6]);
  assign mux_1970_nl = MUX_s_1_2_2(nor_867_nl, mux_1966_nl, fsm_output[5]);
  assign mux_1979_nl = MUX_s_1_2_2(mux_1978_nl, mux_1970_nl, fsm_output[2]);
  assign vec_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_1993_nl,
      mux_1979_nl, fsm_output[4]);
  assign or_2011_nl = (fsm_output[5:4]!=2'b00) | (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b110)
      | (fsm_output[0]) | (~ (VEC_LOOP_j_sva_11_0[0])) | (~ (fsm_output[3])) | (fsm_output[6])
      | (~ (fsm_output[9])) | (fsm_output[8]) | (~ (fsm_output[10]));
  assign or_2009_nl = (~ (fsm_output[5])) | (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b110)
      | (fsm_output[0]) | (~ (VEC_LOOP_j_sva_11_0[0])) | (fsm_output[3]) | (~ (fsm_output[6]))
      | (~ (fsm_output[9])) | (fsm_output[8]) | (fsm_output[10]);
  assign mux_2031_nl = MUX_s_1_2_2(or_2009_nl, mux_tmp_2017, fsm_output[4]);
  assign mux_2032_nl = MUX_s_1_2_2(or_2011_nl, mux_2031_nl, fsm_output[7]);
  assign or_2008_nl = (fsm_output[7]) | mux_tmp_2015;
  assign mux_2033_nl = MUX_s_1_2_2(mux_2032_nl, or_2008_nl, fsm_output[2]);
  assign nand_305_nl = ~((fsm_output[5:4]==2'b11) & (COMP_LOOP_acc_1_cse_6_sva[3:0]==4'b1101)
      & (fsm_output[0]) & (fsm_output[3]) & (fsm_output[6]) & (fsm_output[9]) & (~
      (fsm_output[8])) & (~ (fsm_output[10])));
  assign or_2006_nl = (fsm_output[4]) | mux_tmp_2004;
  assign mux_2029_nl = MUX_s_1_2_2(nand_305_nl, or_2006_nl, fsm_output[7]);
  assign or_2005_nl = (fsm_output[0]) | (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b11) |
      (VEC_LOOP_j_sva_11_0[1:0]!=2'b01) | (fsm_output[3]) | (fsm_output[6]) | (~
      (fsm_output[9])) | (fsm_output[8]) | (fsm_output[10]);
  assign mux_2026_nl = MUX_s_1_2_2(or_2005_nl, or_tmp_1907, fsm_output[5]);
  assign mux_2027_nl = MUX_s_1_2_2(or_tmp_1911, mux_2026_nl, fsm_output[4]);
  assign or_2004_nl = (fsm_output[5:4]!=2'b10) | (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1101)
      | (~ (fsm_output[0])) | (fsm_output[3]) | (~ (fsm_output[6])) | (fsm_output[9])
      | (fsm_output[8]) | (fsm_output[10]);
  assign mux_2028_nl = MUX_s_1_2_2(mux_2027_nl, or_2004_nl, fsm_output[7]);
  assign mux_2030_nl = MUX_s_1_2_2(mux_2029_nl, mux_2028_nl, fsm_output[2]);
  assign mux_2034_nl = MUX_s_1_2_2(mux_2033_nl, mux_2030_nl, fsm_output[1]);
  assign or_2003_nl = (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b110) | (fsm_output[0]) |
      (~ (VEC_LOOP_j_sva_11_0[0])) | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[9]))
      | (fsm_output[8]) | (~ (fsm_output[10]));
  assign mux_2021_nl = MUX_s_1_2_2(or_2003_nl, or_622_cse, fsm_output[5]);
  assign mux_2022_nl = MUX_s_1_2_2(mux_2021_nl, or_621_cse, fsm_output[4]);
  assign or_1994_nl = (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b110) | (fsm_output[0]) |
      (~ (VEC_LOOP_j_sva_11_0[0])) | (fsm_output[3]) | (~ (fsm_output[6])) | (~ (fsm_output[9]))
      | (fsm_output[8]) | (fsm_output[10]);
  assign mux_2018_nl = MUX_s_1_2_2(or_617_cse, or_1994_nl, fsm_output[5]);
  assign mux_2019_nl = MUX_s_1_2_2(mux_2018_nl, mux_tmp_2017, fsm_output[4]);
  assign mux_2023_nl = MUX_s_1_2_2(mux_2022_nl, mux_2019_nl, fsm_output[7]);
  assign mux_2016_nl = MUX_s_1_2_2(mux_tmp_2015, mux_1088_cse, fsm_output[7]);
  assign mux_2024_nl = MUX_s_1_2_2(mux_2023_nl, mux_2016_nl, fsm_output[2]);
  assign nand_307_nl = ~((COMP_LOOP_acc_1_cse_6_sva[3:0]==4'b1101) & (fsm_output[0])
      & (fsm_output[3]) & (fsm_output[6]) & (fsm_output[9]) & (~ (fsm_output[8]))
      & (~ (fsm_output[10])));
  assign mux_2006_nl = MUX_s_1_2_2(or_607_cse, nand_307_nl, fsm_output[5]);
  assign mux_2007_nl = MUX_s_1_2_2(or_609_cse, mux_2006_nl, fsm_output[4]);
  assign mux_2005_nl = MUX_s_1_2_2(mux_tmp_2004, nand_25_cse, fsm_output[4]);
  assign mux_2008_nl = MUX_s_1_2_2(mux_2007_nl, mux_2005_nl, fsm_output[7]);
  assign or_1966_nl = (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b11) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b01)
      | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[9])) | (fsm_output[8])
      | (fsm_output[10]);
  assign mux_1998_nl = MUX_s_1_2_2(or_1966_nl, or_601_cse, fsm_output[0]);
  assign mux_1999_nl = MUX_s_1_2_2(mux_1998_nl, or_tmp_1907, fsm_output[5]);
  assign mux_2000_nl = MUX_s_1_2_2(or_tmp_1911, mux_1999_nl, fsm_output[4]);
  assign or_1959_nl = (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1101) | (~ (fsm_output[0]))
      | (fsm_output[3]) | (~ (fsm_output[6])) | (fsm_output[9]) | (fsm_output[8])
      | (fsm_output[10]);
  assign mux_1996_nl = MUX_s_1_2_2(mux_1073_cse, or_1959_nl, fsm_output[5]);
  assign mux_1997_nl = MUX_s_1_2_2(mux_1996_nl, or_596_cse, fsm_output[4]);
  assign mux_2001_nl = MUX_s_1_2_2(mux_2000_nl, mux_1997_nl, fsm_output[7]);
  assign mux_2009_nl = MUX_s_1_2_2(mux_2008_nl, mux_2001_nl, fsm_output[2]);
  assign mux_2025_nl = MUX_s_1_2_2(mux_2024_nl, mux_2009_nl, fsm_output[1]);
  assign and_611_nl = (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]==4'b1101);
  assign mux_2035_nl = MUX_s_1_2_2(mux_2034_nl, mux_2025_nl, and_611_nl);
  assign vec_rsc_0_13_i_wea_d_pff = ~ mux_2035_nl;
  assign nor_827_cse = ~((z_out_7[4:1]!=4'b1101) | (fsm_output[3]) | (~ (fsm_output[9]))
      | (~ (fsm_output[1])) | (fsm_output[10]));
  assign or_2029_cse = (z_out_7[4:1]!=4'b1101) | (~ (fsm_output[3])) | (~ (fsm_output[9]))
      | (fsm_output[1]) | (fsm_output[10]);
  assign nor_826_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b1101) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[0]) | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[1])
      | (~ (fsm_output[10])));
  assign nor_828_nl = ~((~ (fsm_output[3])) | (z_out_7[4:1]!=4'b1101) | (fsm_output[9])
      | (fsm_output[1]) | (fsm_output[10]));
  assign mux_2062_nl = MUX_s_1_2_2(nor_827_cse, nor_828_nl, fsm_output[0]);
  assign mux_2063_nl = MUX_s_1_2_2(nor_826_nl, mux_2062_nl, fsm_output[8]);
  assign and_606_nl = nor_223_cse & mux_2063_nl;
  assign nand_302_nl = ~((COMP_LOOP_acc_1_cse_6_sva[3:0]==4'b1101) & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm
      & (fsm_output[3]) & (fsm_output[9]) & (fsm_output[1]) & (~ (fsm_output[10])));
  assign or_2056_nl = (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b110) | (~ (VEC_LOOP_j_sva_11_0[0]))
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[3]) | (fsm_output[9])
      | not_tmp_260;
  assign mux_2060_nl = MUX_s_1_2_2(nand_302_nl, or_2056_nl, fsm_output[0]);
  assign nor_829_nl = ~((fsm_output[8:7]!=2'b00) | mux_2060_nl);
  assign nor_830_nl = ~((~ (fsm_output[8])) | (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b1101)
      | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) | (fsm_output[0]) | (fsm_output[3])
      | (fsm_output[9]) | (fsm_output[1]) | (fsm_output[10]));
  assign nor_831_nl = ~((~ (fsm_output[8])) | (fsm_output[0]) | (z_out_7[4:1]!=4'b1101)
      | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[1]) | (~ (fsm_output[10])));
  assign mux_2059_nl = MUX_s_1_2_2(nor_830_nl, nor_831_nl, fsm_output[7]);
  assign mux_2061_nl = MUX_s_1_2_2(nor_829_nl, mux_2059_nl, fsm_output[6]);
  assign mux_2064_nl = MUX_s_1_2_2(and_606_nl, mux_2061_nl, fsm_output[5]);
  assign and_607_nl = (fsm_output[7]) & (~ (fsm_output[8])) & (fsm_output[0]) & (VEC_LOOP_j_sva_11_0[0])
      & (COMP_LOOP_acc_14_psp_sva[2:0]==3'b110) & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm
      & (fsm_output[3]) & (fsm_output[9]) & (fsm_output[1]) & (~ (fsm_output[10]));
  assign or_2048_nl = (z_out_7[4:1]!=4'b1101) | (~ (fsm_output[3])) | (fsm_output[9])
      | (fsm_output[1]) | (~ (fsm_output[10]));
  assign or_2046_nl = (fsm_output[3]) | (z_out_7[4:1]!=4'b1101) | (~ (fsm_output[9]))
      | (fsm_output[1]) | (~ (fsm_output[10]));
  assign mux_2055_nl = MUX_s_1_2_2(or_2048_nl, or_2046_nl, fsm_output[0]);
  assign nor_832_nl = ~((fsm_output[8]) | mux_2055_nl);
  assign nor_833_nl = ~((COMP_LOOP_acc_13_psp_sva[1:0]!=2'b11) | (~ (fsm_output[8]))
      | (~ (fsm_output[0])) | (~ (VEC_LOOP_j_sva_11_0[0])) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (VEC_LOOP_j_sva_11_0[1]) | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[1])
      | (fsm_output[10]));
  assign mux_2056_nl = MUX_s_1_2_2(nor_832_nl, nor_833_nl, fsm_output[7]);
  assign mux_2057_nl = MUX_s_1_2_2(and_607_nl, mux_2056_nl, fsm_output[6]);
  assign nor_834_nl = ~((fsm_output[8:7]!=2'b10) | (z_out_7[4:1]!=4'b1101) | (fsm_output[0])
      | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[1]) | (fsm_output[10]));
  assign and_826_nl = (COMP_LOOP_acc_19_psp_sva[1:0]==2'b11) & (fsm_output[0]) &
      (VEC_LOOP_j_sva_11_0[0]) & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm & (~ (VEC_LOOP_j_sva_11_0[1]))
      & (fsm_output[3]) & (~ (fsm_output[9])) & (~ (fsm_output[1])) & (fsm_output[10]);
  assign nor_836_nl = ~((z_out_7[4:1]!=4'b1101) | (~ (fsm_output[3])) | (fsm_output[9])
      | (~ (fsm_output[1])) | (fsm_output[10]));
  assign mux_2052_nl = MUX_s_1_2_2(nor_836_nl, nor_827_cse, fsm_output[0]);
  assign mux_2053_nl = MUX_s_1_2_2(and_826_nl, mux_2052_nl, fsm_output[8]);
  assign and_608_nl = (fsm_output[7]) & mux_2053_nl;
  assign mux_2054_nl = MUX_s_1_2_2(nor_834_nl, and_608_nl, fsm_output[6]);
  assign mux_2058_nl = MUX_s_1_2_2(mux_2057_nl, mux_2054_nl, fsm_output[5]);
  assign mux_2065_nl = MUX_s_1_2_2(mux_2064_nl, mux_2058_nl, fsm_output[2]);
  assign or_2037_nl = (z_out_7[4:1]!=4'b1101) | (~ (fsm_output[3])) | (fsm_output[9])
      | (~ (fsm_output[1])) | (fsm_output[10]);
  assign or_2036_nl = (z_out_7[4:1]!=4'b1101) | (fsm_output[3]) | (~ (fsm_output[9]))
      | (~ (fsm_output[1])) | (fsm_output[10]);
  assign mux_2048_nl = MUX_s_1_2_2(or_2037_nl, or_2036_nl, fsm_output[0]);
  assign or_2035_nl = (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b1101) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (fsm_output[3]) | (fsm_output[9]) | not_tmp_260;
  assign or_2033_nl = (~ (COMP_LOOP_acc_16_psp_sva[0])) | (~ (VEC_LOOP_j_sva_11_0[2]))
      | (~ (VEC_LOOP_j_sva_11_0[0])) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) |
      (VEC_LOOP_j_sva_11_0[1]) | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[1])
      | (fsm_output[10]);
  assign mux_2047_nl = MUX_s_1_2_2(or_2035_nl, or_2033_nl, fsm_output[0]);
  assign mux_2049_nl = MUX_s_1_2_2(mux_2048_nl, mux_2047_nl, fsm_output[8]);
  assign nor_838_nl = ~((fsm_output[7:6]!=2'b01) | mux_2049_nl);
  assign nor_839_nl = ~((fsm_output[8]) | (~ (VEC_LOOP_j_sva_11_0[3])) | (~ (fsm_output[0]))
      | (VEC_LOOP_j_sva_11_0[2:0]!=3'b101) | (fsm_output[3]) | (fsm_output[9]) |
      (fsm_output[1]) | (fsm_output[10]));
  assign or_2028_nl = (z_out_7[4:1]!=4'b1101) | (fsm_output[3]) | (fsm_output[9])
      | (fsm_output[1]) | (~ (fsm_output[10]));
  assign mux_2044_nl = MUX_s_1_2_2(or_2029_cse, or_2028_nl, fsm_output[0]);
  assign nor_840_nl = ~((fsm_output[8]) | mux_2044_nl);
  assign mux_2045_nl = MUX_s_1_2_2(nor_839_nl, nor_840_nl, fsm_output[7]);
  assign nor_841_nl = ~((~((z_out_7[4:1]==4'b1101) & (fsm_output[8]) & (fsm_output[0])
      & (fsm_output[3]) & (~ (fsm_output[9])))) | not_tmp_260);
  assign nor_842_nl = ~((fsm_output[8]) | (~ (fsm_output[0])) | (~ (VEC_LOOP_j_sva_11_0[0]))
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b110)
      | (~ (fsm_output[3])) | (fsm_output[9]) | (~ (fsm_output[1])) | (fsm_output[10]));
  assign mux_2043_nl = MUX_s_1_2_2(nor_841_nl, nor_842_nl, fsm_output[7]);
  assign mux_2046_nl = MUX_s_1_2_2(mux_2045_nl, mux_2043_nl, fsm_output[6]);
  assign mux_2050_nl = MUX_s_1_2_2(nor_838_nl, mux_2046_nl, fsm_output[5]);
  assign nand_413_nl = ~((COMP_LOOP_acc_1_cse_sva[3:0]==4'b1101) & COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm
      & (~ (fsm_output[0])) & (fsm_output[3]) & (fsm_output[9]) & (~ (fsm_output[1]))
      & (fsm_output[10]));
  assign or_2020_nl = (z_out_7[4:1]!=4'b1101) | (fsm_output[3]) | (fsm_output[9])
      | not_tmp_260;
  assign mux_2039_nl = MUX_s_1_2_2(or_2020_nl, or_2029_cse, fsm_output[0]);
  assign mux_2040_nl = MUX_s_1_2_2(nand_413_nl, mux_2039_nl, fsm_output[8]);
  assign or_2017_nl = (fsm_output[8]) | (fsm_output[0]) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (fsm_output[3]) | (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1101) | (fsm_output[9])
      | (~ (fsm_output[1])) | (fsm_output[10]);
  assign mux_2041_nl = MUX_s_1_2_2(mux_2040_nl, or_2017_nl, fsm_output[7]);
  assign nor_843_nl = ~((fsm_output[6]) | mux_2041_nl);
  assign nor_844_nl = ~((~ (fsm_output[0])) | (z_out_7[4:1]!=4'b1101) | (~ (fsm_output[3]))
      | (fsm_output[9]) | (~ (fsm_output[1])) | (fsm_output[10]));
  assign and_610_nl = (COMP_LOOP_acc_1_cse_10_sva[3:0]==4'b1101) & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm
      & (fsm_output[3]) & (fsm_output[9]) & (fsm_output[1]) & (~ (fsm_output[10]));
  assign nor_845_nl = ~((COMP_LOOP_acc_20_psp_sva[2:0]!=3'b110) | (~ (VEC_LOOP_j_sva_11_0[0]))
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[3]) | (fsm_output[9])
      | not_tmp_260);
  assign mux_2036_nl = MUX_s_1_2_2(and_610_nl, nor_845_nl, fsm_output[0]);
  assign mux_2037_nl = MUX_s_1_2_2(nor_844_nl, mux_2036_nl, fsm_output[8]);
  assign and_609_nl = (fsm_output[7]) & mux_2037_nl;
  assign nor_846_nl = ~((fsm_output[8:7]!=2'b01) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[0]) | (fsm_output[3]) | (COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b1101)
      | (~ (fsm_output[9])) | (fsm_output[1]) | (fsm_output[10]));
  assign mux_2038_nl = MUX_s_1_2_2(and_609_nl, nor_846_nl, fsm_output[6]);
  assign mux_2042_nl = MUX_s_1_2_2(nor_843_nl, mux_2038_nl, fsm_output[5]);
  assign mux_2051_nl = MUX_s_1_2_2(mux_2050_nl, mux_2042_nl, fsm_output[2]);
  assign vec_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_2065_nl,
      mux_2051_nl, fsm_output[4]);
  assign or_2118_nl = (fsm_output[0]) | (VEC_LOOP_j_sva_11_0[0]) | (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b111)
      | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[9])) | (fsm_output[8])
      | (~ (fsm_output[10]));
  assign mux_2102_nl = MUX_s_1_2_2(or_2118_nl, or_622_cse, fsm_output[5]);
  assign mux_2103_nl = MUX_s_1_2_2(mux_2102_nl, or_621_cse, fsm_output[4]);
  assign or_2109_nl = (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b111) | (fsm_output[0]) |
      (VEC_LOOP_j_sva_11_0[0]) | (fsm_output[3]) | (~ (fsm_output[6])) | (~ (fsm_output[9]))
      | (fsm_output[8]) | (fsm_output[10]);
  assign mux_2099_nl = MUX_s_1_2_2(or_617_cse, or_2109_nl, fsm_output[5]);
  assign mux_2100_nl = MUX_s_1_2_2(mux_2099_nl, mux_tmp_2077, fsm_output[4]);
  assign mux_2104_nl = MUX_s_1_2_2(mux_2103_nl, mux_2100_nl, fsm_output[7]);
  assign mux_2098_nl = MUX_s_1_2_2(mux_tmp_2076, mux_1088_cse, fsm_output[7]);
  assign mux_2105_nl = MUX_s_1_2_2(mux_2104_nl, mux_2098_nl, fsm_output[2]);
  assign nand_297_nl = ~((COMP_LOOP_acc_1_cse_6_sva[3:0]==4'b1110) & (fsm_output[0])
      & (fsm_output[3]) & (fsm_output[6]) & (fsm_output[9]) & (~ (fsm_output[8]))
      & (~ (fsm_output[10])));
  assign mux_2091_nl = MUX_s_1_2_2(or_607_cse, nand_297_nl, fsm_output[5]);
  assign mux_2092_nl = MUX_s_1_2_2(or_609_cse, mux_2091_nl, fsm_output[4]);
  assign mux_2090_nl = MUX_s_1_2_2(mux_tmp_2071, nand_25_cse, fsm_output[4]);
  assign mux_2093_nl = MUX_s_1_2_2(mux_2092_nl, mux_2090_nl, fsm_output[7]);
  assign or_2096_nl = (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b11) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b10)
      | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[9])) | (fsm_output[8])
      | (fsm_output[10]);
  assign mux_2085_nl = MUX_s_1_2_2(or_2096_nl, or_601_cse, fsm_output[0]);
  assign mux_2086_nl = MUX_s_1_2_2(mux_2085_nl, or_tmp_2009, fsm_output[5]);
  assign mux_2087_nl = MUX_s_1_2_2(or_tmp_2012, mux_2086_nl, fsm_output[4]);
  assign or_2091_nl = (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1110) | (~ (fsm_output[0]))
      | (fsm_output[3]) | (~ (fsm_output[6])) | (fsm_output[9]) | (fsm_output[8])
      | (fsm_output[10]);
  assign mux_2083_nl = MUX_s_1_2_2(mux_1073_cse, or_2091_nl, fsm_output[5]);
  assign mux_2084_nl = MUX_s_1_2_2(mux_2083_nl, or_596_cse, fsm_output[4]);
  assign mux_2088_nl = MUX_s_1_2_2(mux_2087_nl, mux_2084_nl, fsm_output[7]);
  assign mux_2094_nl = MUX_s_1_2_2(mux_2093_nl, mux_2088_nl, fsm_output[2]);
  assign mux_2106_nl = MUX_s_1_2_2(mux_2105_nl, mux_2094_nl, fsm_output[1]);
  assign or_2088_nl = (fsm_output[4]) | (fsm_output[5]) | (fsm_output[0]) | (VEC_LOOP_j_sva_11_0[0])
      | (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b111) | (~ (fsm_output[3])) | (fsm_output[6])
      | (~ (fsm_output[9])) | (fsm_output[8]) | (~ (fsm_output[10]));
  assign or_2086_nl = (~ (fsm_output[5])) | (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b111)
      | (fsm_output[0]) | (VEC_LOOP_j_sva_11_0[0]) | (fsm_output[3]) | (~ (fsm_output[6]))
      | (~ (fsm_output[9])) | (fsm_output[8]) | (fsm_output[10]);
  assign mux_2078_nl = MUX_s_1_2_2(or_2086_nl, mux_tmp_2077, fsm_output[4]);
  assign mux_2079_nl = MUX_s_1_2_2(or_2088_nl, mux_2078_nl, fsm_output[7]);
  assign or_2082_nl = (fsm_output[7]) | mux_tmp_2076;
  assign mux_2080_nl = MUX_s_1_2_2(mux_2079_nl, or_2082_nl, fsm_output[2]);
  assign nand_298_nl = ~((fsm_output[5:4]==2'b11) & (COMP_LOOP_acc_1_cse_6_sva[3:0]==4'b1110)
      & (fsm_output[0]) & (fsm_output[3]) & (fsm_output[6]) & (fsm_output[9]) & (~
      (fsm_output[8])) & (~ (fsm_output[10])));
  assign or_2074_nl = (fsm_output[4]) | mux_tmp_2071;
  assign mux_2072_nl = MUX_s_1_2_2(nand_298_nl, or_2074_nl, fsm_output[7]);
  assign or_2067_nl = (fsm_output[0]) | (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b11) |
      (VEC_LOOP_j_sva_11_0[1:0]!=2'b10) | (fsm_output[3]) | (fsm_output[6]) | (~
      (fsm_output[9])) | (fsm_output[8]) | (fsm_output[10]);
  assign mux_2067_nl = MUX_s_1_2_2(or_2067_nl, or_tmp_2009, fsm_output[5]);
  assign mux_2068_nl = MUX_s_1_2_2(or_tmp_2012, mux_2067_nl, fsm_output[4]);
  assign or_2064_nl = (fsm_output[5:4]!=2'b10) | (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1110)
      | (~ (fsm_output[0])) | (fsm_output[3]) | (~ (fsm_output[6])) | (fsm_output[9])
      | (fsm_output[8]) | (fsm_output[10]);
  assign mux_2069_nl = MUX_s_1_2_2(mux_2068_nl, or_2064_nl, fsm_output[7]);
  assign mux_2073_nl = MUX_s_1_2_2(mux_2072_nl, mux_2069_nl, fsm_output[2]);
  assign mux_2081_nl = MUX_s_1_2_2(mux_2080_nl, mux_2073_nl, fsm_output[1]);
  assign nand_299_nl = ~((COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]==4'b1110));
  assign mux_2107_nl = MUX_s_1_2_2(mux_2106_nl, mux_2081_nl, nand_299_nl);
  assign vec_rsc_0_14_i_wea_d_pff = ~ mux_2107_nl;
  assign nor_804_cse = ~((z_out_7[4:1]!=4'b1110) | (fsm_output[3]) | (~ (fsm_output[9]))
      | (~ (fsm_output[1])) | (fsm_output[10]));
  assign or_2136_cse = (z_out_7[4:1]!=4'b1110) | (~ (fsm_output[3])) | (~ (fsm_output[9]))
      | (fsm_output[1]) | (fsm_output[10]);
  assign nor_803_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b1110) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[0]) | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[1])
      | (~ (fsm_output[10])));
  assign nor_805_nl = ~((z_out_7[4:1]!=4'b1110) | (~ (fsm_output[3])) | (fsm_output[9])
      | (fsm_output[1]) | (fsm_output[10]));
  assign mux_2134_nl = MUX_s_1_2_2(nor_804_cse, nor_805_nl, fsm_output[0]);
  assign mux_2135_nl = MUX_s_1_2_2(nor_803_nl, mux_2134_nl, fsm_output[8]);
  assign and_601_nl = nor_223_cse & mux_2135_nl;
  assign nand_293_nl = ~((COMP_LOOP_acc_1_cse_6_sva[3:0]==4'b1110) & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm
      & (fsm_output[3]) & (fsm_output[9]) & (fsm_output[1]) & (~ (fsm_output[10])));
  assign or_2163_nl = (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b111) | (VEC_LOOP_j_sva_11_0[0])
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[3]) | (fsm_output[9])
      | not_tmp_260;
  assign mux_2132_nl = MUX_s_1_2_2(nand_293_nl, or_2163_nl, fsm_output[0]);
  assign nor_806_nl = ~((fsm_output[8:7]!=2'b00) | mux_2132_nl);
  assign nor_807_nl = ~((~ (fsm_output[8])) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b1110) | (fsm_output[0]) | (fsm_output[3])
      | (fsm_output[9]) | (fsm_output[1]) | (fsm_output[10]));
  assign nor_808_nl = ~((~ (fsm_output[8])) | (fsm_output[0]) | (z_out_7[4:1]!=4'b1110)
      | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[1]) | (~ (fsm_output[10])));
  assign mux_2131_nl = MUX_s_1_2_2(nor_807_nl, nor_808_nl, fsm_output[7]);
  assign mux_2133_nl = MUX_s_1_2_2(nor_806_nl, mux_2131_nl, fsm_output[6]);
  assign mux_2136_nl = MUX_s_1_2_2(and_601_nl, mux_2133_nl, fsm_output[5]);
  assign and_602_nl = (fsm_output[7]) & (~ (fsm_output[8])) & (fsm_output[0]) & (~
      (VEC_LOOP_j_sva_11_0[0])) & (COMP_LOOP_acc_14_psp_sva[2:0]==3'b111) & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm
      & (fsm_output[3]) & (fsm_output[9]) & (fsm_output[1]) & (~ (fsm_output[10]));
  assign or_2155_nl = (z_out_7[4:1]!=4'b1110) | (~ (fsm_output[3])) | (fsm_output[9])
      | (fsm_output[1]) | (~ (fsm_output[10]));
  assign or_2153_nl = (fsm_output[3]) | (z_out_7[4:1]!=4'b1110) | (~ (fsm_output[9]))
      | (fsm_output[1]) | (~ (fsm_output[10]));
  assign mux_2127_nl = MUX_s_1_2_2(or_2155_nl, or_2153_nl, fsm_output[0]);
  assign nor_809_nl = ~((fsm_output[8]) | mux_2127_nl);
  assign nor_810_nl = ~((COMP_LOOP_acc_13_psp_sva[1:0]!=2'b11) | (~ (fsm_output[8]))
      | (~ (fsm_output[0])) | (VEC_LOOP_j_sva_11_0[0]) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (~ (VEC_LOOP_j_sva_11_0[1])) | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[1])
      | (fsm_output[10]));
  assign mux_2128_nl = MUX_s_1_2_2(nor_809_nl, nor_810_nl, fsm_output[7]);
  assign mux_2129_nl = MUX_s_1_2_2(and_602_nl, mux_2128_nl, fsm_output[6]);
  assign nor_811_nl = ~((fsm_output[8:7]!=2'b10) | (z_out_7[4:1]!=4'b1110) | (fsm_output[0])
      | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[1]) | (fsm_output[10]));
  assign and_825_nl = (COMP_LOOP_acc_19_psp_sva[1:0]==2'b11) & (fsm_output[0]) &
      (~ (VEC_LOOP_j_sva_11_0[0])) & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm & (VEC_LOOP_j_sva_11_0[1])
      & (fsm_output[3]) & (~ (fsm_output[9])) & (~ (fsm_output[1])) & (fsm_output[10]);
  assign nor_813_nl = ~((z_out_7[4:1]!=4'b1110) | (~ (fsm_output[3])) | (fsm_output[9])
      | (~ (fsm_output[1])) | (fsm_output[10]));
  assign mux_2124_nl = MUX_s_1_2_2(nor_813_nl, nor_804_cse, fsm_output[0]);
  assign mux_2125_nl = MUX_s_1_2_2(and_825_nl, mux_2124_nl, fsm_output[8]);
  assign and_603_nl = (fsm_output[7]) & mux_2125_nl;
  assign mux_2126_nl = MUX_s_1_2_2(nor_811_nl, and_603_nl, fsm_output[6]);
  assign mux_2130_nl = MUX_s_1_2_2(mux_2129_nl, mux_2126_nl, fsm_output[5]);
  assign mux_2137_nl = MUX_s_1_2_2(mux_2136_nl, mux_2130_nl, fsm_output[2]);
  assign or_2144_nl = (z_out_7[4:1]!=4'b1110) | (~ (fsm_output[3])) | (fsm_output[9])
      | (~ (fsm_output[1])) | (fsm_output[10]);
  assign or_2143_nl = (z_out_7[4:1]!=4'b1110) | (fsm_output[3]) | (~ (fsm_output[9]))
      | (~ (fsm_output[1])) | (fsm_output[10]);
  assign mux_2120_nl = MUX_s_1_2_2(or_2144_nl, or_2143_nl, fsm_output[0]);
  assign or_2142_nl = (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b1110) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (fsm_output[3]) | (fsm_output[9]) | not_tmp_260;
  assign or_2140_nl = (~ (COMP_LOOP_acc_16_psp_sva[0])) | (~ (VEC_LOOP_j_sva_11_0[2]))
      | (VEC_LOOP_j_sva_11_0[0]) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (~
      (VEC_LOOP_j_sva_11_0[1])) | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[1])
      | (fsm_output[10]);
  assign mux_2119_nl = MUX_s_1_2_2(or_2142_nl, or_2140_nl, fsm_output[0]);
  assign mux_2121_nl = MUX_s_1_2_2(mux_2120_nl, mux_2119_nl, fsm_output[8]);
  assign nor_815_nl = ~((fsm_output[7:6]!=2'b01) | mux_2121_nl);
  assign nor_816_nl = ~((fsm_output[8]) | (~ (VEC_LOOP_j_sva_11_0[3])) | (~ (fsm_output[0]))
      | (VEC_LOOP_j_sva_11_0[2:0]!=3'b110) | (fsm_output[3]) | (fsm_output[9]) |
      (fsm_output[1]) | (fsm_output[10]));
  assign or_2135_nl = (z_out_7[4:1]!=4'b1110) | (fsm_output[3]) | (fsm_output[9])
      | (fsm_output[1]) | (~ (fsm_output[10]));
  assign mux_2116_nl = MUX_s_1_2_2(or_2136_cse, or_2135_nl, fsm_output[0]);
  assign nor_817_nl = ~((fsm_output[8]) | mux_2116_nl);
  assign mux_2117_nl = MUX_s_1_2_2(nor_816_nl, nor_817_nl, fsm_output[7]);
  assign nor_818_nl = ~((~((z_out_7[4:1]==4'b1110) & (fsm_output[8]) & (fsm_output[0])
      & (fsm_output[3]) & (~ (fsm_output[9])))) | not_tmp_260);
  assign nor_819_nl = ~((fsm_output[8]) | (~ (fsm_output[0])) | (VEC_LOOP_j_sva_11_0[0])
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b111)
      | (~ (fsm_output[3])) | (fsm_output[9]) | (~ (fsm_output[1])) | (fsm_output[10]));
  assign mux_2115_nl = MUX_s_1_2_2(nor_818_nl, nor_819_nl, fsm_output[7]);
  assign mux_2118_nl = MUX_s_1_2_2(mux_2117_nl, mux_2115_nl, fsm_output[6]);
  assign mux_2122_nl = MUX_s_1_2_2(nor_815_nl, mux_2118_nl, fsm_output[5]);
  assign nand_411_nl = ~((COMP_LOOP_acc_1_cse_sva[3:0]==4'b1110) & COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm
      & (~ (fsm_output[0])) & (fsm_output[3]) & (fsm_output[9]) & (~ (fsm_output[1]))
      & (fsm_output[10]));
  assign or_2127_nl = (z_out_7[4:1]!=4'b1110) | (fsm_output[3]) | (fsm_output[9])
      | not_tmp_260;
  assign mux_2111_nl = MUX_s_1_2_2(or_2127_nl, or_2136_cse, fsm_output[0]);
  assign mux_2112_nl = MUX_s_1_2_2(nand_411_nl, mux_2111_nl, fsm_output[8]);
  assign or_2124_nl = (fsm_output[8]) | (fsm_output[0]) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (fsm_output[3]) | (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1110) | (fsm_output[9])
      | (~ (fsm_output[1])) | (fsm_output[10]);
  assign mux_2113_nl = MUX_s_1_2_2(mux_2112_nl, or_2124_nl, fsm_output[7]);
  assign nor_820_nl = ~((fsm_output[6]) | mux_2113_nl);
  assign nor_821_nl = ~((~ (fsm_output[0])) | (z_out_7[4:1]!=4'b1110) | (~ (fsm_output[3]))
      | (fsm_output[9]) | (~ (fsm_output[1])) | (fsm_output[10]));
  assign and_605_nl = (COMP_LOOP_acc_1_cse_10_sva[3:0]==4'b1110) & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm
      & (fsm_output[3]) & (fsm_output[9]) & (fsm_output[1]) & (~ (fsm_output[10]));
  assign nor_822_nl = ~((COMP_LOOP_acc_20_psp_sva[2:0]!=3'b111) | (VEC_LOOP_j_sva_11_0[0])
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[3]) | (fsm_output[9])
      | not_tmp_260);
  assign mux_2108_nl = MUX_s_1_2_2(and_605_nl, nor_822_nl, fsm_output[0]);
  assign mux_2109_nl = MUX_s_1_2_2(nor_821_nl, mux_2108_nl, fsm_output[8]);
  assign and_604_nl = (fsm_output[7]) & mux_2109_nl;
  assign nor_823_nl = ~((fsm_output[8:7]!=2'b01) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[0]) | (fsm_output[3]) | (COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b1110)
      | (~ (fsm_output[9])) | (fsm_output[1]) | (fsm_output[10]));
  assign mux_2110_nl = MUX_s_1_2_2(and_604_nl, nor_823_nl, fsm_output[6]);
  assign mux_2114_nl = MUX_s_1_2_2(nor_820_nl, mux_2110_nl, fsm_output[5]);
  assign mux_2123_nl = MUX_s_1_2_2(mux_2122_nl, mux_2114_nl, fsm_output[2]);
  assign vec_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_2137_nl,
      mux_2123_nl, fsm_output[4]);
  assign or_2224_nl = (fsm_output[4]) | (fsm_output[5]) | (fsm_output[0]) | (~ (VEC_LOOP_j_sva_11_0[0]))
      | (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b111) | (~ (fsm_output[3])) | (fsm_output[6])
      | (~ (fsm_output[9])) | (fsm_output[8]) | (~ (fsm_output[10]));
  assign or_2222_nl = (~ (fsm_output[5])) | (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b111)
      | (fsm_output[0]) | (~ (VEC_LOOP_j_sva_11_0[0])) | (fsm_output[3]) | (~ (fsm_output[6]))
      | (~ (fsm_output[9])) | (fsm_output[8]) | (fsm_output[10]);
  assign mux_2175_nl = MUX_s_1_2_2(or_2222_nl, mux_tmp_2161, fsm_output[4]);
  assign mux_2176_nl = MUX_s_1_2_2(or_2224_nl, mux_2175_nl, fsm_output[7]);
  assign or_2221_nl = (fsm_output[7]) | mux_tmp_2159;
  assign mux_2177_nl = MUX_s_1_2_2(mux_2176_nl, or_2221_nl, fsm_output[2]);
  assign nand_284_nl = ~((fsm_output[5:4]==2'b11) & (COMP_LOOP_acc_1_cse_6_sva[3:0]==4'b1111)
      & (fsm_output[0]) & (fsm_output[3]) & (fsm_output[6]) & (fsm_output[9]) & (~
      (fsm_output[8])) & (~ (fsm_output[10])));
  assign or_2219_nl = (fsm_output[4]) | mux_tmp_2148;
  assign mux_2173_nl = MUX_s_1_2_2(nand_284_nl, or_2219_nl, fsm_output[7]);
  assign or_2218_nl = (fsm_output[0]) | (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b11) |
      (VEC_LOOP_j_sva_11_0[1:0]!=2'b11) | (fsm_output[3]) | (fsm_output[6]) | (~
      (fsm_output[9])) | (fsm_output[8]) | (fsm_output[10]);
  assign mux_2170_nl = MUX_s_1_2_2(or_2218_nl, or_tmp_2120, fsm_output[5]);
  assign mux_2171_nl = MUX_s_1_2_2(or_tmp_2124, mux_2170_nl, fsm_output[4]);
  assign or_2217_nl = (fsm_output[5:4]!=2'b10) | (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1111)
      | (~ (fsm_output[0])) | (fsm_output[3]) | (~ (fsm_output[6])) | (fsm_output[9])
      | (fsm_output[8]) | (fsm_output[10]);
  assign mux_2172_nl = MUX_s_1_2_2(mux_2171_nl, or_2217_nl, fsm_output[7]);
  assign mux_2174_nl = MUX_s_1_2_2(mux_2173_nl, mux_2172_nl, fsm_output[2]);
  assign mux_2178_nl = MUX_s_1_2_2(mux_2177_nl, mux_2174_nl, fsm_output[1]);
  assign nand_438_nl = ~((~ (fsm_output[0])) & (VEC_LOOP_j_sva_11_0[0]) & (COMP_LOOP_acc_20_psp_sva[2:0]==3'b111)
      & (fsm_output[3]) & (~ (fsm_output[6])) & (fsm_output[9]) & (~ (fsm_output[8]))
      & (fsm_output[10]));
  assign mux_2165_nl = MUX_s_1_2_2(nand_438_nl, or_622_cse, fsm_output[5]);
  assign mux_2166_nl = MUX_s_1_2_2(mux_2165_nl, or_621_cse, fsm_output[4]);
  assign or_2207_nl = (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b111) | (fsm_output[0]) |
      (~ (VEC_LOOP_j_sva_11_0[0])) | (fsm_output[3]) | (~ (fsm_output[6])) | (~ (fsm_output[9]))
      | (fsm_output[8]) | (fsm_output[10]);
  assign mux_2162_nl = MUX_s_1_2_2(or_617_cse, or_2207_nl, fsm_output[5]);
  assign mux_2163_nl = MUX_s_1_2_2(mux_2162_nl, mux_tmp_2161, fsm_output[4]);
  assign mux_2167_nl = MUX_s_1_2_2(mux_2166_nl, mux_2163_nl, fsm_output[7]);
  assign mux_2160_nl = MUX_s_1_2_2(mux_tmp_2159, mux_1088_cse, fsm_output[7]);
  assign mux_2168_nl = MUX_s_1_2_2(mux_2167_nl, mux_2160_nl, fsm_output[2]);
  assign nand_286_nl = ~((COMP_LOOP_acc_1_cse_6_sva[3:0]==4'b1111) & (fsm_output[0])
      & (fsm_output[3]) & (fsm_output[6]) & (fsm_output[9]) & (~ (fsm_output[8]))
      & (~ (fsm_output[10])));
  assign mux_2150_nl = MUX_s_1_2_2(or_607_cse, nand_286_nl, fsm_output[5]);
  assign mux_2151_nl = MUX_s_1_2_2(or_609_cse, mux_2150_nl, fsm_output[4]);
  assign mux_2149_nl = MUX_s_1_2_2(mux_tmp_2148, nand_25_cse, fsm_output[4]);
  assign mux_2152_nl = MUX_s_1_2_2(mux_2151_nl, mux_2149_nl, fsm_output[7]);
  assign or_2179_nl = (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b11) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b11)
      | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[9])) | (fsm_output[8])
      | (fsm_output[10]);
  assign mux_2142_nl = MUX_s_1_2_2(or_2179_nl, or_601_cse, fsm_output[0]);
  assign mux_2143_nl = MUX_s_1_2_2(mux_2142_nl, or_tmp_2120, fsm_output[5]);
  assign mux_2144_nl = MUX_s_1_2_2(or_tmp_2124, mux_2143_nl, fsm_output[4]);
  assign or_2172_nl = (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1111) | (~ (fsm_output[0]))
      | (fsm_output[3]) | (~ (fsm_output[6])) | (fsm_output[9]) | (fsm_output[8])
      | (fsm_output[10]);
  assign mux_2140_nl = MUX_s_1_2_2(mux_1073_cse, or_2172_nl, fsm_output[5]);
  assign mux_2141_nl = MUX_s_1_2_2(mux_2140_nl, or_596_cse, fsm_output[4]);
  assign mux_2145_nl = MUX_s_1_2_2(mux_2144_nl, mux_2141_nl, fsm_output[7]);
  assign mux_2153_nl = MUX_s_1_2_2(mux_2152_nl, mux_2145_nl, fsm_output[2]);
  assign mux_2169_nl = MUX_s_1_2_2(mux_2168_nl, mux_2153_nl, fsm_output[1]);
  assign and_600_nl = (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]==4'b1111);
  assign mux_2179_nl = MUX_s_1_2_2(mux_2178_nl, mux_2169_nl, and_600_nl);
  assign vec_rsc_0_15_i_wea_d_pff = ~ mux_2179_nl;
  assign and_591_cse = (z_out_7[4:1]==4'b1111) & (~ (fsm_output[3])) & (fsm_output[9])
      & (fsm_output[1]) & (~ (fsm_output[10]));
  assign nand_278_cse = ~((z_out_7[4:1]==4'b1111) & (fsm_output[3]) & (fsm_output[9])
      & (~ (fsm_output[1])) & (~ (fsm_output[10])));
  assign and_823_nl = (COMP_LOOP_acc_1_cse_12_sva[3:0]==4'b1111) & COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm
      & (~ (fsm_output[0])) & (fsm_output[3]) & (~ (fsm_output[9])) & (~ (fsm_output[1]))
      & (fsm_output[10]);
  assign nor_786_nl = ~((~ (fsm_output[3])) | (z_out_7[4:1]!=4'b1111) | (fsm_output[9])
      | (fsm_output[1]) | (fsm_output[10]));
  assign mux_2206_nl = MUX_s_1_2_2(and_591_cse, nor_786_nl, fsm_output[0]);
  assign mux_2207_nl = MUX_s_1_2_2(and_823_nl, mux_2206_nl, fsm_output[8]);
  assign and_590_nl = nor_223_cse & mux_2207_nl;
  assign nand_269_nl = ~((COMP_LOOP_acc_1_cse_6_sva[3:0]==4'b1111) & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm
      & (fsm_output[3]) & (fsm_output[9]) & (fsm_output[1]) & (~ (fsm_output[10])));
  assign or_2269_nl = (~((COMP_LOOP_acc_17_psp_sva[2:0]==3'b111) & (VEC_LOOP_j_sva_11_0[0])
      & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm & (~ (fsm_output[3])) & (~ (fsm_output[9]))))
      | not_tmp_260;
  assign mux_2204_nl = MUX_s_1_2_2(nand_269_nl, or_2269_nl, fsm_output[0]);
  assign nor_787_nl = ~((fsm_output[8:7]!=2'b00) | mux_2204_nl);
  assign nor_788_nl = ~((~ (fsm_output[8])) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b1111) | (fsm_output[0]) | (fsm_output[3])
      | (fsm_output[9]) | (fsm_output[1]) | (fsm_output[10]));
  assign nor_789_nl = ~((~ (fsm_output[8])) | (fsm_output[0]) | (z_out_7[4:1]!=4'b1111)
      | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[1]) | (~ (fsm_output[10])));
  assign mux_2203_nl = MUX_s_1_2_2(nor_788_nl, nor_789_nl, fsm_output[7]);
  assign mux_2205_nl = MUX_s_1_2_2(nor_787_nl, mux_2203_nl, fsm_output[6]);
  assign mux_2208_nl = MUX_s_1_2_2(and_590_nl, mux_2205_nl, fsm_output[5]);
  assign and_592_nl = (fsm_output[7]) & (~ (fsm_output[8])) & (fsm_output[0]) & (VEC_LOOP_j_sva_11_0[0])
      & (COMP_LOOP_acc_14_psp_sva[2:0]==3'b111) & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm
      & (fsm_output[3]) & (fsm_output[9]) & (fsm_output[1]) & (~ (fsm_output[10]));
  assign nand_436_nl = ~((z_out_7[4:1]==4'b1111) & (fsm_output[3]) & (~ (fsm_output[9]))
      & (~ (fsm_output[1])) & (fsm_output[10]));
  assign nand_434_nl = ~((~ (fsm_output[3])) & (z_out_7[4:1]==4'b1111) & (fsm_output[9])
      & (~ (fsm_output[1])) & (fsm_output[10]));
  assign mux_2199_nl = MUX_s_1_2_2(nand_436_nl, nand_434_nl, fsm_output[0]);
  assign nor_790_nl = ~((fsm_output[8]) | mux_2199_nl);
  assign nor_791_nl = ~((COMP_LOOP_acc_13_psp_sva[1:0]!=2'b11) | (~ (fsm_output[8]))
      | (~ (fsm_output[0])) | (~ (VEC_LOOP_j_sva_11_0[0])) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (~ (VEC_LOOP_j_sva_11_0[1])) | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[1])
      | (fsm_output[10]));
  assign mux_2200_nl = MUX_s_1_2_2(nor_790_nl, nor_791_nl, fsm_output[7]);
  assign mux_2201_nl = MUX_s_1_2_2(and_592_nl, mux_2200_nl, fsm_output[6]);
  assign nor_792_nl = ~((fsm_output[8:7]!=2'b10) | (z_out_7[4:1]!=4'b1111) | (fsm_output[0])
      | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[1]) | (fsm_output[10]));
  assign and_824_nl = (COMP_LOOP_acc_19_psp_sva[1:0]==2'b11) & (fsm_output[0]) &
      (VEC_LOOP_j_sva_11_0[0]) & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm & (VEC_LOOP_j_sva_11_0[1])
      & (fsm_output[3]) & (~ (fsm_output[9])) & (~ (fsm_output[1])) & (fsm_output[10]);
  assign and_594_nl = (z_out_7[4:1]==4'b1111) & (fsm_output[3]) & (~ (fsm_output[9]))
      & (fsm_output[1]) & (~ (fsm_output[10]));
  assign mux_2196_nl = MUX_s_1_2_2(and_594_nl, and_591_cse, fsm_output[0]);
  assign mux_2197_nl = MUX_s_1_2_2(and_824_nl, mux_2196_nl, fsm_output[8]);
  assign and_593_nl = (fsm_output[7]) & mux_2197_nl;
  assign mux_2198_nl = MUX_s_1_2_2(nor_792_nl, and_593_nl, fsm_output[6]);
  assign mux_2202_nl = MUX_s_1_2_2(mux_2201_nl, mux_2198_nl, fsm_output[5]);
  assign mux_2209_nl = MUX_s_1_2_2(mux_2208_nl, mux_2202_nl, fsm_output[2]);
  assign nand_274_nl = ~((z_out_7[4:1]==4'b1111) & (fsm_output[3]) & (~ (fsm_output[9]))
      & (fsm_output[1]) & (~ (fsm_output[10])));
  assign nand_275_nl = ~((z_out_7[4:1]==4'b1111) & (~ (fsm_output[3])) & (fsm_output[9])
      & (fsm_output[1]) & (~ (fsm_output[10])));
  assign mux_2192_nl = MUX_s_1_2_2(nand_274_nl, nand_275_nl, fsm_output[0]);
  assign or_2248_nl = (~((COMP_LOOP_acc_1_cse_14_sva[3:0]==4'b1111) & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm
      & (~ (fsm_output[3])) & (~ (fsm_output[9])))) | not_tmp_260;
  assign nand_277_nl = ~((COMP_LOOP_acc_16_psp_sva[0]) & (VEC_LOOP_j_sva_11_0[2])
      & (VEC_LOOP_j_sva_11_0[0]) & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm & (VEC_LOOP_j_sva_11_0[1])
      & (fsm_output[3]) & (fsm_output[9]) & (~ (fsm_output[1])) & (~ (fsm_output[10])));
  assign mux_2191_nl = MUX_s_1_2_2(or_2248_nl, nand_277_nl, fsm_output[0]);
  assign mux_2193_nl = MUX_s_1_2_2(mux_2192_nl, mux_2191_nl, fsm_output[8]);
  assign nor_794_nl = ~((fsm_output[7:6]!=2'b01) | mux_2193_nl);
  assign nor_795_nl = ~((fsm_output[8]) | (~ (VEC_LOOP_j_sva_11_0[3])) | (~ (fsm_output[0]))
      | (VEC_LOOP_j_sva_11_0[2:0]!=3'b111) | (fsm_output[3]) | (fsm_output[9]) |
      (fsm_output[1]) | (fsm_output[10]));
  assign or_2241_nl = (z_out_7[4:1]!=4'b1111) | (fsm_output[3]) | (fsm_output[9])
      | (fsm_output[1]) | (~ (fsm_output[10]));
  assign mux_2188_nl = MUX_s_1_2_2(nand_278_cse, or_2241_nl, fsm_output[0]);
  assign nor_796_nl = ~((fsm_output[8]) | mux_2188_nl);
  assign mux_2189_nl = MUX_s_1_2_2(nor_795_nl, nor_796_nl, fsm_output[7]);
  assign nor_797_nl = ~((~((z_out_7[4:1]==4'b1111) & (fsm_output[8]) & (fsm_output[0])
      & (fsm_output[3]) & (~ (fsm_output[9])))) | not_tmp_260);
  assign and_596_nl = (~ (fsm_output[8])) & (fsm_output[0]) & (VEC_LOOP_j_sva_11_0[0])
      & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm & (COMP_LOOP_acc_11_psp_sva[2:0]==3'b111)
      & (fsm_output[3]) & (~ (fsm_output[9])) & (fsm_output[1]) & (~ (fsm_output[10]));
  assign mux_2187_nl = MUX_s_1_2_2(nor_797_nl, and_596_nl, fsm_output[7]);
  assign mux_2190_nl = MUX_s_1_2_2(mux_2189_nl, mux_2187_nl, fsm_output[6]);
  assign mux_2194_nl = MUX_s_1_2_2(nor_794_nl, mux_2190_nl, fsm_output[5]);
  assign nand_409_nl = ~((COMP_LOOP_acc_1_cse_sva[3:0]==4'b1111) & COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm
      & (~ (fsm_output[0])) & (fsm_output[3]) & (fsm_output[9]) & (~ (fsm_output[1]))
      & (fsm_output[10]));
  assign or_2233_nl = (z_out_7[4:1]!=4'b1111) | (fsm_output[3]) | (fsm_output[9])
      | not_tmp_260;
  assign mux_2183_nl = MUX_s_1_2_2(or_2233_nl, nand_278_cse, fsm_output[0]);
  assign mux_2184_nl = MUX_s_1_2_2(nand_409_nl, mux_2183_nl, fsm_output[8]);
  assign or_2230_nl = (fsm_output[8]) | (fsm_output[0]) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (fsm_output[3]) | (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1111) | (fsm_output[9])
      | (~ (fsm_output[1])) | (fsm_output[10]);
  assign mux_2185_nl = MUX_s_1_2_2(mux_2184_nl, or_2230_nl, fsm_output[7]);
  assign nor_798_nl = ~((fsm_output[6]) | mux_2185_nl);
  assign and_598_nl = (fsm_output[0]) & (z_out_7[4:1]==4'b1111) & (fsm_output[3])
      & (~ (fsm_output[9])) & (fsm_output[1]) & (~ (fsm_output[10]));
  assign and_599_nl = (COMP_LOOP_acc_1_cse_10_sva[3:0]==4'b1111) & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm
      & (fsm_output[3]) & (fsm_output[9]) & (fsm_output[1]) & (~ (fsm_output[10]));
  assign nor_799_nl = ~((~((COMP_LOOP_acc_20_psp_sva[2:0]==3'b111) & (VEC_LOOP_j_sva_11_0[0])
      & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm & (~ (fsm_output[3])) & (~ (fsm_output[9]))))
      | not_tmp_260);
  assign mux_2180_nl = MUX_s_1_2_2(and_599_nl, nor_799_nl, fsm_output[0]);
  assign mux_2181_nl = MUX_s_1_2_2(and_598_nl, mux_2180_nl, fsm_output[8]);
  assign and_597_nl = (fsm_output[7]) & mux_2181_nl;
  assign nor_800_nl = ~((fsm_output[8:7]!=2'b01) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[0]) | (fsm_output[3]) | (COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b1111)
      | (~ (fsm_output[9])) | (fsm_output[1]) | (fsm_output[10]));
  assign mux_2182_nl = MUX_s_1_2_2(and_597_nl, nor_800_nl, fsm_output[6]);
  assign mux_2186_nl = MUX_s_1_2_2(nor_798_nl, mux_2182_nl, fsm_output[5]);
  assign mux_2195_nl = MUX_s_1_2_2(mux_2194_nl, mux_2186_nl, fsm_output[2]);
  assign vec_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_2209_nl,
      mux_2195_nl, fsm_output[4]);
  assign and_dcpl_348 = ~((fsm_output[3:2]!=2'b00));
  assign and_dcpl_350 = and_dcpl_348 & (~ (fsm_output[1])) & and_dcpl_107;
  assign and_dcpl_351 = ~((fsm_output[8:7]!=2'b00));
  assign and_dcpl_353 = (fsm_output[4]) & (~ (fsm_output[10]));
  assign and_dcpl_354 = and_dcpl_353 & (~ (fsm_output[9]));
  assign and_dcpl_356 = and_dcpl_354 & and_dcpl_351 & (fsm_output[5]) & and_dcpl_350;
  assign and_dcpl_358 = (fsm_output[3:2]==2'b10);
  assign and_dcpl_359 = and_dcpl_358 & (fsm_output[1]);
  assign and_dcpl_361 = and_dcpl_351 & (~ (fsm_output[5]));
  assign and_850_cse = and_dcpl_354 & and_dcpl_361 & and_dcpl_359 & and_dcpl_121;
  assign and_dcpl_365 = and_459_cse & (fsm_output[1]);
  assign and_dcpl_368 = (~ (fsm_output[8])) & (fsm_output[7]) & (fsm_output[5]);
  assign and_857_cse = and_dcpl_354 & and_dcpl_368 & and_dcpl_365 & and_dcpl_107;
  assign and_dcpl_373 = (fsm_output[8:7]==2'b11);
  assign and_dcpl_374 = and_dcpl_373 & (~ (fsm_output[5]));
  assign and_dcpl_375 = ~((fsm_output[4]) | (fsm_output[10]));
  assign and_dcpl_376 = and_dcpl_375 & (~ (fsm_output[9]));
  assign and_dcpl_378 = and_dcpl_376 & and_dcpl_374 & and_dcpl_358 & (~ (fsm_output[1]))
      & and_dcpl_107;
  assign and_dcpl_380 = and_dcpl_373 & (fsm_output[5]);
  assign and_869_cse = and_dcpl_376 & and_dcpl_380 & and_dcpl_365 & and_dcpl_121;
  assign and_dcpl_384 = and_dcpl_348 & (fsm_output[1]);
  assign and_dcpl_386 = and_dcpl_353 & (fsm_output[9]);
  assign and_875_cse = and_dcpl_386 & and_dcpl_361 & and_dcpl_384 & nor_tmp_217;
  assign and_dcpl_391 = (fsm_output[8:7]==2'b10);
  assign and_dcpl_392 = and_dcpl_391 & (~ (fsm_output[5]));
  assign and_dcpl_394 = and_dcpl_386 & and_dcpl_392 & and_459_cse & (~ (fsm_output[1]))
      & and_dcpl_107;
  assign and_dcpl_397 = and_dcpl_375 & (fsm_output[9]);
  assign and_886_cse = and_dcpl_397 & and_dcpl_374 & and_dcpl_384 & and_dcpl_99;
  assign and_dcpl_401 = (fsm_output[3:1]==3'b011);
  assign and_dcpl_404 = and_dcpl_397 & and_dcpl_380 & and_dcpl_401 & nor_tmp_217;
  assign and_dcpl_406 = (fsm_output[4]) & (fsm_output[10]) & (~ (fsm_output[9]));
  assign and_dcpl_408 = and_dcpl_406 & and_dcpl_368 & and_dcpl_350;
  assign and_dcpl_411 = and_dcpl_406 & and_dcpl_392 & and_dcpl_401 & and_dcpl_99;
  assign and_dcpl_415 = and_dcpl_406 & and_dcpl_391 & (fsm_output[5]) & and_dcpl_359
      & nor_tmp_217;
  assign and_dcpl_430 = (fsm_output[8]) & (~ (fsm_output[7])) & (~ (fsm_output[5]));
  assign and_dcpl_433 = and_dcpl_353 & (fsm_output[9]) & and_dcpl_430 & (fsm_output[3:1]==3'b110)
      & and_dcpl_107;
  assign and_dcpl_441 = (fsm_output[10]) & (fsm_output[4]) & (~ (fsm_output[9]))
      & and_dcpl_430 & (~ (fsm_output[3])) & (fsm_output[2]) & (fsm_output[1]) &
      (~ (fsm_output[6])) & (~ (fsm_output[0]));
  assign and_dcpl_480 = (fsm_output[3:1]==3'b010);
  assign and_dcpl_502 = ~((fsm_output[8]) | (fsm_output[7]) | (fsm_output[5]));
  assign and_dcpl_503 = (fsm_output[10]) & (~ (fsm_output[4]));
  assign and_dcpl_511 = and_dcpl_503 & (fsm_output[9]) & and_dcpl_502 & and_dcpl_480
      & (fsm_output[6]) & (fsm_output[0]);
  assign and_dcpl_517 = (fsm_output[8]) & (fsm_output[7]) & (fsm_output[5]);
  assign and_dcpl_555 = (~ (fsm_output[10])) & (fsm_output[4]) & (~ (fsm_output[9]))
      & and_dcpl_351 & (fsm_output[5]) & (~ (fsm_output[3])) & (~ (fsm_output[2]))
      & (~ (fsm_output[1])) & (~ (fsm_output[6])) & (fsm_output[0]);
  assign not_tmp_930 = ~((fsm_output[6]) & (fsm_output[2]) & (fsm_output[7]));
  assign nand_450_nl = ~((fsm_output[9]) & (fsm_output[3]) & (fsm_output[6]) & (fsm_output[2])
      & (fsm_output[7]));
  assign or_3357_nl = (~ (fsm_output[9])) | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[2])
      | (fsm_output[7]);
  assign mux_tmp = MUX_s_1_2_2(nand_450_nl, or_3357_nl, fsm_output[1]);
  assign not_tmp_933 = ~((fsm_output[2]) & (fsm_output[7]));
  assign nand_439_nl = ~((fsm_output[0]) & (~ mux_tmp));
  assign or_3373_nl = (fsm_output[0]) | (~ (fsm_output[1])) | (fsm_output[9]) | (fsm_output[3])
      | not_tmp_930;
  assign mux_3721_nl = MUX_s_1_2_2(nand_439_nl, or_3373_nl, fsm_output[10]);
  assign or_3371_nl = (fsm_output[0]) | (fsm_output[1]) | (fsm_output[9]) | (fsm_output[3])
      | not_tmp_930;
  assign or_3369_nl = (fsm_output[0]) | (~ (fsm_output[1])) | (~ (fsm_output[9]))
      | (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[2]) | (fsm_output[7]);
  assign mux_3720_nl = MUX_s_1_2_2(or_3371_nl, or_3369_nl, fsm_output[10]);
  assign mux_3722_nl = MUX_s_1_2_2(mux_3721_nl, mux_3720_nl, fsm_output[4]);
  assign or_3367_nl = (fsm_output[1]) | (~ (fsm_output[9])) | (~ (fsm_output[3]))
      | (~ (fsm_output[6])) | (fsm_output[2]) | (fsm_output[7]);
  assign or_3366_nl = (~ (fsm_output[1])) | (fsm_output[9]) | (~ (fsm_output[3]))
      | (~ (fsm_output[6])) | (~ (fsm_output[2])) | (fsm_output[7]);
  assign mux_3718_nl = MUX_s_1_2_2(or_3367_nl, or_3366_nl, fsm_output[0]);
  assign or_3365_nl = (~ (fsm_output[0])) | (fsm_output[1]) | (fsm_output[9]) | (fsm_output[3])
      | (~ (fsm_output[6])) | (fsm_output[2]) | (fsm_output[7]);
  assign mux_3719_nl = MUX_s_1_2_2(mux_3718_nl, or_3365_nl, fsm_output[10]);
  assign or_3368_nl = (fsm_output[4]) | mux_3719_nl;
  assign mux_3723_nl = MUX_s_1_2_2(mux_3722_nl, or_3368_nl, fsm_output[5]);
  assign nor_1381_nl = ~((~ (fsm_output[1])) | (fsm_output[9]) | (~ (fsm_output[3]))
      | (fsm_output[6]) | not_tmp_933);
  assign nor_1382_nl = ~((~ (fsm_output[1])) | (~ (fsm_output[9])) | (fsm_output[3])
      | (fsm_output[6]) | not_tmp_933);
  assign mux_3715_nl = MUX_s_1_2_2(nor_1381_nl, nor_1382_nl, fsm_output[0]);
  assign nor_1383_nl = ~((fsm_output[0]) | (fsm_output[1]) | (fsm_output[9]) | (fsm_output[3])
      | (fsm_output[6]) | (fsm_output[2]) | (~ (fsm_output[7])));
  assign mux_3716_nl = MUX_s_1_2_2(mux_3715_nl, nor_1383_nl, fsm_output[10]);
  assign nand_445_nl = ~((fsm_output[4]) & mux_3716_nl);
  assign or_3358_nl = (~ (fsm_output[10])) | (~ (fsm_output[0])) | (~ (fsm_output[1]))
      | (fsm_output[9]) | (~ (fsm_output[3])) | (fsm_output[6]) | (fsm_output[2])
      | (fsm_output[7]);
  assign or_3356_nl = (fsm_output[1]) | (fsm_output[9]) | (~ (fsm_output[3])) | (fsm_output[6])
      | (fsm_output[2]) | (fsm_output[7]);
  assign mux_3712_nl = MUX_s_1_2_2(mux_tmp, or_3356_nl, fsm_output[0]);
  assign or_3355_nl = (~ (fsm_output[0])) | (fsm_output[1]) | (fsm_output[9]) | (fsm_output[3])
      | not_tmp_930;
  assign mux_3713_nl = MUX_s_1_2_2(mux_3712_nl, or_3355_nl, fsm_output[10]);
  assign mux_3714_nl = MUX_s_1_2_2(or_3358_nl, mux_3713_nl, fsm_output[4]);
  assign mux_3717_nl = MUX_s_1_2_2(nand_445_nl, mux_3714_nl, fsm_output[5]);
  assign mux_3724_itm = MUX_s_1_2_2(mux_3723_nl, mux_3717_nl, fsm_output[8]);
  assign and_dcpl_564 = ~((fsm_output[10]) | (fsm_output[4]) | (fsm_output[9]) |
      (~ and_dcpl_351) | (fsm_output[5]) | (~ (fsm_output[3])) | (fsm_output[2])
      | (~ (fsm_output[1])) | (fsm_output[6]) | (fsm_output[0]));
  assign and_dcpl_568 = and_dcpl_348 & (~ (fsm_output[1])) & (~ (fsm_output[6]))
      & (fsm_output[0]);
  assign and_dcpl_574 = (fsm_output[4]) & (~ (fsm_output[10])) & (~ (fsm_output[9]))
      & and_dcpl_351 & (fsm_output[5]) & and_dcpl_568;
  assign or_tmp_3188 = (fsm_output[10:6]!=5'b01000);
  assign or_tmp_3189 = (fsm_output[10:6]!=5'b01001);
  assign mux_tmp_3724 = MUX_s_1_2_2(or_tmp_3189, or_tmp_3188, fsm_output[2]);
  assign or_tmp_3191 = (fsm_output[6]) | (fsm_output[9]) | (fsm_output[8]) | (fsm_output[10]);
  assign or_tmp_3193 = (fsm_output[6]) | (fsm_output[9]) | not_tmp_51;
  assign mux_tmp_3725 = MUX_s_1_2_2(or_tmp_3193, or_tmp_3191, fsm_output[7]);
  assign or_tmp_3195 = (~ (fsm_output[6])) | (fsm_output[9]) | not_tmp_51;
  assign or_tmp_3196 = (~ (fsm_output[6])) | (fsm_output[9]) | (~ (fsm_output[8]))
      | (fsm_output[10]);
  assign mux_tmp_3728 = MUX_s_1_2_2(or_tmp_3196, or_tmp_3195, fsm_output[7]);
  assign or_tmp_3200 = (fsm_output[10:6]!=5'b10000);
  assign or_tmp_3202 = (fsm_output[10:6]!=5'b10001);
  assign or_tmp_3203 = (~ (fsm_output[6])) | (fsm_output[9]) | (fsm_output[8]) |
      (fsm_output[10]);
  assign mux_tmp_3733 = MUX_s_1_2_2(or_tmp_3195, or_tmp_3203, fsm_output[7]);
  assign or_tmp_3204 = (fsm_output[10:6]!=5'b01101);
  assign or_tmp_3205 = (fsm_output[10:6]!=5'b01110);
  assign mux_tmp_3735 = MUX_s_1_2_2(or_tmp_3205, or_tmp_3204, fsm_output[2]);
  assign nand_455_nl = ~((fsm_output[6]) & (fsm_output[9]) & (~ (fsm_output[8]))
      & (fsm_output[10]));
  assign mux_tmp_3737 = MUX_s_1_2_2(nand_455_nl, or_tmp_3196, fsm_output[7]);
  assign or_tmp_3211 = (fsm_output[10:6]!=5'b01011);
  assign or_3396_nl = (fsm_output[10:6]!=5'b01010);
  assign mux_tmp_3742 = MUX_s_1_2_2(or_tmp_3211, or_3396_nl, fsm_output[2]);
  assign or_tmp_3212 = (fsm_output[6]) | (fsm_output[9]) | (~ (fsm_output[8])) |
      (fsm_output[10]);
  assign mux_tmp_3743 = MUX_s_1_2_2(or_tmp_3212, or_tmp_3193, fsm_output[7]);
  assign or_tmp_3213 = ~((fsm_output[10:6]==5'b01111));
  assign or_tmp_3218 = (fsm_output[10:6]!=5'b01100);
  assign mux_tmp_3751 = MUX_s_1_2_2(or_tmp_3200, or_tmp_3213, fsm_output[2]);
  assign or_3406_nl = (~ (fsm_output[6])) | (fsm_output[9]) | (fsm_output[8]) | (~
      (fsm_output[10]));
  assign mux_tmp_3753 = MUX_s_1_2_2(or_tmp_3203, or_3406_nl, fsm_output[7]);
  assign or_3409_nl = (fsm_output[6]) | (fsm_output[9]) | (fsm_output[8]) | (~ (fsm_output[10]));
  assign mux_tmp_3762 = MUX_s_1_2_2(or_tmp_3191, or_3409_nl, fsm_output[7]);
  assign or_3413_nl = (fsm_output[6]) | (~ (fsm_output[9])) | (fsm_output[8]) | (~
      (fsm_output[10]));
  assign mux_3771_nl = MUX_s_1_2_2(or_3413_nl, or_tmp_3212, fsm_output[7]);
  assign mux_tmp_3771 = MUX_s_1_2_2(mux_3771_nl, mux_tmp_3728, fsm_output[2]);
  assign or_3420_nl = (fsm_output[10:6]!=5'b11010);
  assign mux_3783_nl = MUX_s_1_2_2(or_3420_nl, mux_tmp_3737, fsm_output[2]);
  assign or_3418_nl = (fsm_output[10:6]!=5'b00011);
  assign mux_3782_nl = MUX_s_1_2_2(mux_tmp_3743, or_3418_nl, fsm_output[2]);
  assign mux_3784_nl = MUX_s_1_2_2(mux_3783_nl, mux_3782_nl, fsm_output[4]);
  assign mux_3780_nl = MUX_s_1_2_2(mux_tmp_3762, or_tmp_3202, fsm_output[2]);
  assign mux_3781_nl = MUX_s_1_2_2(mux_tmp_3742, mux_3780_nl, fsm_output[4]);
  assign mux_3785_nl = MUX_s_1_2_2(mux_3784_nl, mux_3781_nl, fsm_output[5]);
  assign or_3417_nl = (fsm_output[7]) | (~ (fsm_output[6])) | (fsm_output[9]) | not_tmp_51;
  assign mux_3777_nl = MUX_s_1_2_2(or_3417_nl, mux_tmp_3725, fsm_output[2]);
  assign mux_3778_nl = MUX_s_1_2_2(mux_tmp_3735, mux_3777_nl, fsm_output[4]);
  assign or_3415_nl = (fsm_output[2]) | (fsm_output[7]) | (~ (fsm_output[6])) | (fsm_output[9])
      | (fsm_output[8]) | (~ (fsm_output[10]));
  assign mux_3776_nl = MUX_s_1_2_2(or_3415_nl, mux_tmp_3771, fsm_output[4]);
  assign mux_3779_nl = MUX_s_1_2_2(mux_3778_nl, mux_3776_nl, fsm_output[5]);
  assign mux_3786_nl = MUX_s_1_2_2(mux_3785_nl, mux_3779_nl, fsm_output[0]);
  assign mux_3770_nl = MUX_s_1_2_2(or_tmp_3204, or_tmp_3218, fsm_output[2]);
  assign mux_3773_nl = MUX_s_1_2_2(mux_tmp_3771, mux_3770_nl, fsm_output[4]);
  assign or_3411_nl = (fsm_output[10:6]!=5'b10011);
  assign mux_3768_nl = MUX_s_1_2_2(or_tmp_3189, or_3411_nl, fsm_output[2]);
  assign mux_3769_nl = MUX_s_1_2_2(mux_3768_nl, mux_tmp_3751, fsm_output[4]);
  assign mux_3774_nl = MUX_s_1_2_2(mux_3773_nl, mux_3769_nl, fsm_output[5]);
  assign mux_3765_nl = MUX_s_1_2_2(or_tmp_3218, or_tmp_3211, fsm_output[2]);
  assign mux_3764_nl = MUX_s_1_2_2(mux_tmp_3753, mux_tmp_3762, fsm_output[2]);
  assign mux_3766_nl = MUX_s_1_2_2(mux_3765_nl, mux_3764_nl, fsm_output[4]);
  assign mux_3761_nl = MUX_s_1_2_2(or_tmp_3188, mux_tmp_3737, fsm_output[2]);
  assign or_3407_nl = (fsm_output[10:6]!=5'b00100);
  assign mux_3760_nl = MUX_s_1_2_2(or_3407_nl, or_tmp_3205, fsm_output[2]);
  assign mux_3762_nl = MUX_s_1_2_2(mux_3761_nl, mux_3760_nl, fsm_output[4]);
  assign mux_3767_nl = MUX_s_1_2_2(mux_3766_nl, mux_3762_nl, fsm_output[5]);
  assign mux_3775_nl = MUX_s_1_2_2(mux_3774_nl, mux_3767_nl, fsm_output[0]);
  assign mux_3787_nl = MUX_s_1_2_2(mux_3786_nl, mux_3775_nl, fsm_output[3]);
  assign mux_3755_nl = MUX_s_1_2_2(mux_tmp_3725, mux_tmp_3753, fsm_output[2]);
  assign mux_3756_nl = MUX_s_1_2_2(mux_3755_nl, mux_tmp_3724, fsm_output[4]);
  assign or_3403_nl = (~ (fsm_output[7])) | (fsm_output[6]) | (fsm_output[9]) | not_tmp_51;
  assign mux_3751_nl = MUX_s_1_2_2(or_tmp_3218, or_3403_nl, fsm_output[2]);
  assign mux_3753_nl = MUX_s_1_2_2(mux_tmp_3751, mux_3751_nl, fsm_output[4]);
  assign mux_3757_nl = MUX_s_1_2_2(mux_3756_nl, mux_3753_nl, fsm_output[5]);
  assign or_3401_nl = (fsm_output[10:6]!=5'b10010);
  assign mux_3748_nl = MUX_s_1_2_2(or_tmp_3188, or_3401_nl, fsm_output[2]);
  assign mux_3747_nl = MUX_s_1_2_2(or_tmp_3213, or_tmp_3205, fsm_output[2]);
  assign mux_3749_nl = MUX_s_1_2_2(mux_3748_nl, mux_3747_nl, fsm_output[4]);
  assign mux_3745_nl = MUX_s_1_2_2(mux_tmp_3743, mux_tmp_3733, fsm_output[2]);
  assign mux_3746_nl = MUX_s_1_2_2(mux_3745_nl, mux_tmp_3742, fsm_output[4]);
  assign mux_3750_nl = MUX_s_1_2_2(mux_3749_nl, mux_3746_nl, fsm_output[5]);
  assign mux_3758_nl = MUX_s_1_2_2(mux_3757_nl, mux_3750_nl, fsm_output[0]);
  assign or_3395_nl = (~ (fsm_output[2])) | (~ (fsm_output[7])) | (fsm_output[6])
      | (~ (fsm_output[9])) | (fsm_output[8]) | (fsm_output[10]);
  assign or_3392_nl = (fsm_output[10:6]!=5'b00110);
  assign mux_3739_nl = MUX_s_1_2_2(mux_tmp_3737, or_3392_nl, fsm_output[2]);
  assign mux_3740_nl = MUX_s_1_2_2(or_3395_nl, mux_3739_nl, fsm_output[4]);
  assign mux_3735_nl = MUX_s_1_2_2(mux_tmp_3733, mux_tmp_3725, fsm_output[2]);
  assign mux_3737_nl = MUX_s_1_2_2(mux_tmp_3735, mux_3735_nl, fsm_output[4]);
  assign mux_3741_nl = MUX_s_1_2_2(mux_3740_nl, mux_3737_nl, fsm_output[5]);
  assign mux_3731_nl = MUX_s_1_2_2(or_tmp_3202, or_tmp_3200, fsm_output[2]);
  assign or_3384_nl = (fsm_output[10:6]!=5'b11000);
  assign mux_3730_nl = MUX_s_1_2_2(or_3384_nl, mux_tmp_3728, fsm_output[2]);
  assign mux_3732_nl = MUX_s_1_2_2(mux_3731_nl, mux_3730_nl, fsm_output[4]);
  assign or_3376_nl = (fsm_output[10:6]!=5'b00001);
  assign mux_3727_nl = MUX_s_1_2_2(mux_tmp_3725, or_3376_nl, fsm_output[2]);
  assign mux_3728_nl = MUX_s_1_2_2(mux_3727_nl, mux_tmp_3724, fsm_output[4]);
  assign mux_3733_nl = MUX_s_1_2_2(mux_3732_nl, mux_3728_nl, fsm_output[5]);
  assign mux_3742_nl = MUX_s_1_2_2(mux_3741_nl, mux_3733_nl, fsm_output[0]);
  assign mux_3759_nl = MUX_s_1_2_2(mux_3758_nl, mux_3742_nl, fsm_output[3]);
  assign mux_3788_itm = MUX_s_1_2_2(mux_3787_nl, mux_3759_nl, fsm_output[1]);
  assign and_dcpl_579 = (~ (fsm_output[4])) & (~ (fsm_output[10])) & (~ (fsm_output[9]))
      & and_dcpl_351 & (~ (fsm_output[5])) & and_dcpl_568;
  assign and_dcpl_588 = (~ (fsm_output[4])) & (fsm_output[10]) & (fsm_output[9])
      & (~ (fsm_output[8])) & (fsm_output[7]) & (~ (fsm_output[5])) & and_dcpl_348
      & (fsm_output[1]) & (~ (fsm_output[6])) & (~ (fsm_output[0]));
  assign and_dcpl_591 = and_dcpl_348 & (~ (fsm_output[1]));
  assign and_dcpl_592 = and_dcpl_591 & and_dcpl_107;
  assign and_dcpl_598 = and_dcpl_354 & and_dcpl_351 & (fsm_output[5]) & and_dcpl_592;
  assign and_dcpl_614 = (fsm_output[3:2]==2'b01);
  assign and_dcpl_615 = and_dcpl_614 & (~ (fsm_output[1]));
  assign and_dcpl_618 = and_dcpl_391 & (fsm_output[5]);
  assign and_dcpl_622 = and_dcpl_376 & and_dcpl_618 & and_dcpl_615 & and_dcpl_99;
  assign and_dcpl_623 = and_dcpl_358 & (~ (fsm_output[1]));
  assign and_dcpl_624 = and_dcpl_623 & and_dcpl_107;
  assign and_dcpl_628 = and_dcpl_376 & and_dcpl_374 & and_dcpl_624;
  assign and_dcpl_641 = and_dcpl_386 & and_dcpl_368 & and_dcpl_623 & and_dcpl_99;
  assign and_dcpl_642 = and_459_cse & (~ (fsm_output[1]));
  assign and_dcpl_646 = and_dcpl_386 & and_dcpl_392 & and_dcpl_642 & and_dcpl_107;
  assign and_dcpl_651 = and_dcpl_614 & (fsm_output[1]);
  assign and_dcpl_654 = and_dcpl_397 & and_dcpl_380 & and_dcpl_651 & nor_tmp_217;
  assign and_dcpl_657 = and_dcpl_503 & (~ (fsm_output[9]));
  assign and_dcpl_659 = and_dcpl_657 & and_dcpl_361 & and_dcpl_642 & and_dcpl_121;
  assign and_dcpl_663 = and_dcpl_406 & and_dcpl_368 & and_dcpl_592;
  assign and_dcpl_666 = and_dcpl_406 & and_dcpl_392 & and_dcpl_651 & and_dcpl_99;
  assign and_dcpl_669 = and_dcpl_406 & and_dcpl_618 & and_dcpl_359 & nor_tmp_217;
  assign and_dcpl_672 = and_dcpl_657 & and_dcpl_380 & and_dcpl_591 & and_dcpl_121;
  assign and_dcpl_676 = and_dcpl_503 & (fsm_output[9]) & and_dcpl_361 & and_dcpl_615
      & nor_tmp_217;
  assign and_dcpl_678 = and_dcpl_376 & and_dcpl_361 & and_dcpl_624;
  assign and_dcpl_688 = ~((fsm_output!=11'b00100100100));
  assign and_dcpl_698 = (~ (fsm_output[4])) & (fsm_output[10]) & (~ (fsm_output[9]))
      & and_dcpl_351 & (~ (fsm_output[5])) & (fsm_output[3]) & (fsm_output[2]) &
      (~ (fsm_output[1])) & (fsm_output[6]) & (~ (fsm_output[0]));
  assign nor_1369_nl = ~((fsm_output[10]) | (~((fsm_output[9]) & (fsm_output[1])
      & (fsm_output[0]) & (fsm_output[3]) & (fsm_output[8]) & (fsm_output[6]))));
  assign nor_1370_nl = ~((fsm_output[1]) | (fsm_output[0]) | (fsm_output[3]) | nand_257_cse);
  assign nor_1371_nl = ~((~ (fsm_output[1])) | (fsm_output[0]) | (~ (fsm_output[3]))
      | (fsm_output[8]) | (fsm_output[6]));
  assign mux_3799_nl = MUX_s_1_2_2(nor_1370_nl, nor_1371_nl, fsm_output[9]);
  assign and_1249_nl = (fsm_output[10]) & mux_3799_nl;
  assign mux_3800_nl = MUX_s_1_2_2(nor_1369_nl, and_1249_nl, fsm_output[2]);
  assign and_1248_nl = (fsm_output[4]) & mux_3800_nl;
  assign or_3441_nl = (fsm_output[10]) | (fsm_output[9]) | (~ (fsm_output[1])) |
      (fsm_output[0]) | (fsm_output[3]) | nand_257_cse;
  assign or_3439_nl = (~ (fsm_output[9])) | (fsm_output[1]) | (fsm_output[0]) | (~
      (fsm_output[3])) | (fsm_output[8]) | (fsm_output[6]);
  assign or_3438_nl = (fsm_output[9]) | (fsm_output[1]) | (~ (fsm_output[0])) | (fsm_output[3])
      | (fsm_output[8]) | (fsm_output[6]);
  assign mux_3797_nl = MUX_s_1_2_2(or_3439_nl, or_3438_nl, fsm_output[10]);
  assign mux_3798_nl = MUX_s_1_2_2(or_3441_nl, mux_3797_nl, fsm_output[2]);
  assign nor_1372_nl = ~((fsm_output[4]) | mux_3798_nl);
  assign mux_3801_nl = MUX_s_1_2_2(and_1248_nl, nor_1372_nl, fsm_output[5]);
  assign nor_1373_nl = ~((~ (fsm_output[9])) | (fsm_output[1]) | (fsm_output[0])
      | (fsm_output[3]) | nand_257_cse);
  assign nor_1374_nl = ~((fsm_output[9]) | (~ (fsm_output[1])) | (fsm_output[0])
      | (~ (fsm_output[3])) | (fsm_output[8]) | (fsm_output[6]));
  assign mux_3793_nl = MUX_s_1_2_2(nor_1373_nl, nor_1374_nl, fsm_output[10]);
  assign nor_1375_nl = ~((fsm_output[10]) | (fsm_output[9]) | (~ (fsm_output[1]))
      | (~ (fsm_output[0])) | (fsm_output[3]) | nand_257_cse);
  assign mux_3794_nl = MUX_s_1_2_2(mux_3793_nl, nor_1375_nl, fsm_output[2]);
  assign or_3431_nl = (fsm_output[1]) | (fsm_output[0]) | (~ (fsm_output[3])) | (fsm_output[8])
      | (fsm_output[6]);
  assign or_3430_nl = (fsm_output[1]) | (~ (fsm_output[0])) | (fsm_output[3]) | (fsm_output[8])
      | (fsm_output[6]);
  assign mux_3792_nl = MUX_s_1_2_2(or_3431_nl, or_3430_nl, fsm_output[9]);
  assign nor_1376_nl = ~((fsm_output[2]) | (fsm_output[10]) | mux_3792_nl);
  assign mux_3795_nl = MUX_s_1_2_2(mux_3794_nl, nor_1376_nl, fsm_output[4]);
  assign and_1250_nl = (fsm_output[2]) & (fsm_output[10]) & (~ (fsm_output[9])) &
      (fsm_output[1]) & (fsm_output[0]) & (fsm_output[3]) & (~ (fsm_output[8])) &
      (fsm_output[6]);
  assign nor_1378_nl = ~((~ (fsm_output[10])) | (fsm_output[9]) | (fsm_output[1])
      | (~ (fsm_output[0])) | (~ (fsm_output[3])) | (~ (fsm_output[8])) | (fsm_output[6]));
  assign or_3424_nl = (fsm_output[1]) | (~ (fsm_output[0])) | (~ (fsm_output[3]))
      | (fsm_output[8]) | (~ (fsm_output[6]));
  assign or_3422_nl = (~ (fsm_output[1])) | (fsm_output[0]) | (fsm_output[3]) | (fsm_output[8])
      | (~ (fsm_output[6]));
  assign mux_3789_nl = MUX_s_1_2_2(or_3424_nl, or_3422_nl, fsm_output[9]);
  assign nor_1379_nl = ~((fsm_output[10]) | mux_3789_nl);
  assign mux_3790_nl = MUX_s_1_2_2(nor_1378_nl, nor_1379_nl, fsm_output[2]);
  assign mux_3791_nl = MUX_s_1_2_2(and_1250_nl, mux_3790_nl, fsm_output[4]);
  assign mux_3796_nl = MUX_s_1_2_2(mux_3795_nl, mux_3791_nl, fsm_output[5]);
  assign not_tmp_980 = MUX_s_1_2_2(mux_3801_nl, mux_3796_nl, fsm_output[7]);
  assign and_dcpl_707 = (fsm_output[4]) & (~ (fsm_output[10])) & (~ (fsm_output[9]))
      & and_dcpl_351 & (fsm_output[5]) & (~ (fsm_output[3])) & (~ (fsm_output[2]))
      & (fsm_output[1]) & (~ (fsm_output[6])) & (fsm_output[0]);
  assign and_dcpl_717 = and_dcpl_353 & (fsm_output[9]) & (~ (fsm_output[8])) & (fsm_output[7])
      & (fsm_output[5]) & and_dcpl_358 & (~ (fsm_output[1])) & and_dcpl_99;
  assign and_dcpl_727 = (fsm_output[10]) & (~ (fsm_output[4])) & (~ (fsm_output[9]))
      & and_dcpl_373 & (fsm_output[5]) & and_dcpl_348 & (~ (fsm_output[1])) & and_dcpl_121;
  assign and_dcpl_734 = and_dcpl_353 & (~ (fsm_output[9])) & (~ (fsm_output[8]))
      & (~ (fsm_output[7])) & (~ (fsm_output[5])) & and_dcpl_358 & (fsm_output[1])
      & and_dcpl_121;
  assign and_dcpl_741 = (~ (fsm_output[10])) & (~ (fsm_output[4])) & (fsm_output[9])
      & and_dcpl_373 & (~ (fsm_output[5])) & and_dcpl_348 & (fsm_output[1]) & and_dcpl_99;
  assign COMP_LOOP_or_55_ssc = and_857_cse | and_dcpl_628 | and_875_cse | and_dcpl_672;
  assign COMP_LOOP_or_56_ssc = and_dcpl_622 | and_dcpl_641 | and_dcpl_659 | and_dcpl_676;
  assign COMP_LOOP_or_57_ssc = and_869_cse | and_dcpl_654 | and_dcpl_663 | and_dcpl_669;
  assign COMP_LOOP_or_58_ssc = and_dcpl_646 | and_dcpl_666;
  assign or_tmp = (fsm_output[9]) | (~ (fsm_output[4]));
  assign nor_tmp = (fsm_output[2]) & (fsm_output[4]);
  assign mux_tmp_3818 = MUX_s_1_2_2((~ (fsm_output[4])), (fsm_output[4]), fsm_output[2]);
  assign not_tmp_1007 = ~((fsm_output[2]) | (fsm_output[4]));
  assign mux_tmp_3819 = MUX_s_1_2_2(not_tmp_1007, mux_tmp_3818, fsm_output[0]);
  assign mux_tmp_3822 = MUX_s_1_2_2(mux_tmp_3818, nor_tmp, or_2348_cse);
  assign or_tmp_3291 = and_563_cse | (fsm_output[4]);
  assign or_tmp_3293 = (fsm_output[9]) | (~ or_tmp_3291);
  assign nor_tmp_535 = ((fsm_output[9]) | (fsm_output[2])) & (fsm_output[4]);
  assign nor_tmp_536 = or_2348_cse & (fsm_output[2]) & (fsm_output[4]);
  assign mux_tmp_3828 = MUX_s_1_2_2((~ or_tmp_3291), nor_tmp_536, fsm_output[9]);
  assign mux_tmp_3834 = MUX_s_1_2_2(mux_tmp_3822, (fsm_output[4]), fsm_output[9]);
  assign nor_tmp_539 = or_3280_cse & (fsm_output[4]);
  assign nor_tmp_540 = or_2385_cse & (fsm_output[4]);
  assign or_tmp_3303 = and_573_cse | (fsm_output[2]) | (fsm_output[4]);
  assign or_tmp_3304 = ((fsm_output[9]) & (fsm_output[2])) | (fsm_output[4]);
  assign mux_tmp_3846 = MUX_s_1_2_2(mux_tmp_3818, nor_tmp, fsm_output[0]);
  assign mux_tmp_3853 = MUX_s_1_2_2((~ or_tmp_3291), nor_tmp_540, fsm_output[9]);
  assign not_tmp_1021 = ~(((fsm_output[9]) & (fsm_output[1]) & (fsm_output[0]) &
      (fsm_output[2])) | (fsm_output[4]));
  assign nor_1460_nl = ~((fsm_output[0]) | (fsm_output[2]) | (fsm_output[4]));
  assign and_1267_nl = (fsm_output[0]) & (fsm_output[2]) & (fsm_output[4]);
  assign mux_tmp_3861 = MUX_s_1_2_2(nor_1460_nl, and_1267_nl, fsm_output[1]);
  assign mux_tmp_3878 = MUX_s_1_2_2(mux_tmp_3819, mux_tmp_3846, fsm_output[1]);
  assign or_tmp_3320 = (fsm_output[1]) | (~ COMP_LOOP_nor_11_itm) | (~ (fsm_output[8]))
      | (fsm_output[10]) | (fsm_output[9]) | (fsm_output[4]);
  assign not_tmp_1034 = ~((fsm_output[9]) & (fsm_output[4]));
  assign or_tmp_3327 = (fsm_output[10]) | not_tmp_1034;
  assign mux_3898_nl = MUX_s_1_2_2(or_tmp_3327, or_tmp_2652, fsm_output[8]);
  assign or_3516_nl = (~ COMP_LOOP_nor_11_itm) | (fsm_output[8]) | (fsm_output[10])
      | not_tmp_1034;
  assign mux_tmp_3898 = MUX_s_1_2_2(mux_3898_nl, or_3516_nl, fsm_output[1]);
  assign or_tmp_3332 = (fsm_output[8]) | (fsm_output[10]) | (~ (fsm_output[9])) |
      (fsm_output[4]);
  assign nand_470_nl = ~(COMP_LOOP_nor_11_itm & (fsm_output[8]) & (fsm_output[10])
      & (~ (fsm_output[9])) & (fsm_output[4]));
  assign mux_3902_nl = MUX_s_1_2_2(or_tmp_3332, nand_470_nl, fsm_output[1]);
  assign nand_tmp = ~((fsm_output[6]) & (~ mux_3902_nl));
  assign mux_tmp_3902 = MUX_s_1_2_2(or_tmp_195, or_tmp_3327, fsm_output[8]);
  assign or_3531_nl = (fsm_output[8]) | (~ (fsm_output[10])) | (fsm_output[9]) |
      (fsm_output[4]);
  assign mux_3906_nl = MUX_s_1_2_2(or_tmp, or_2747_cse, fsm_output[10]);
  assign or_3530_nl = (fsm_output[8]) | mux_3906_nl;
  assign mux_tmp_3906 = MUX_s_1_2_2(or_3531_nl, or_3530_nl, COMP_LOOP_nor_11_itm);
  assign or_tmp_3343 = (~ (fsm_output[1])) | (fsm_output[8]) | (fsm_output[10]) |
      (fsm_output[9]) | (fsm_output[4]);
  assign mux_tmp_3915 = MUX_s_1_2_2(or_2415_cse, or_tmp_182, fsm_output[8]);
  assign or_tmp_3369 = (fsm_output[8]) | (fsm_output[10]) | (fsm_output[9]) | (~
      (fsm_output[4]));
  assign COMP_LOOP_or_60_itm = and_850_cse | and_857_cse | and_dcpl_378 | and_869_cse
      | and_875_cse | and_dcpl_394 | and_886_cse | and_dcpl_404 | and_dcpl_408 |
      and_dcpl_411 | and_dcpl_415;
  assign COMP_LOOP_or_24_itm = and_dcpl_433 | and_dcpl_441;
  assign COMP_LOOP_COMP_LOOP_or_6_cse = (~ and_dcpl_441) | (and_dcpl_353 & (~ (fsm_output[9]))
      & and_dcpl_351 & (fsm_output[5]) & nor_738_cse & and_dcpl_107) | and_dcpl_433;
  assign COMP_LOOP_or_67_itm = and_dcpl_688 | and_dcpl_698;
  assign COMP_LOOP_COMP_LOOP_or_9_cse = (~(and_dcpl_688 | and_dcpl_698)) | not_tmp_980
      | and_dcpl_707;
  assign COMP_LOOP_nor_680_itm = ~(not_tmp_980 | and_dcpl_707);
  always @(posedge clk) begin
    if ( ~ not_tmp_219 ) begin
      p_sva <= p_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( (and_dcpl_103 & and_dcpl_98) | STAGE_LOOP_i_3_0_sva_mx0c1 ) begin
      STAGE_LOOP_i_3_0_sva <= MUX_v_4_2_2(4'b0001, STAGE_LOOP_i_3_0_sva_2, STAGE_LOOP_i_3_0_sva_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ not_tmp_219 ) begin
      r_sva <= r_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_vec_rsc_triosy_0_15_obj_ld_cse <= 1'b0;
      COMP_LOOP_nor_11_itm <= 1'b0;
      modExp_exp_1_7_1_sva <= 1'b0;
      COMP_LOOP_nor_12_itm <= 1'b0;
      COMP_LOOP_nor_134_itm <= 1'b0;
      COMP_LOOP_nor_137_itm <= 1'b0;
      COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_nor_1_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_139_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_140_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_141_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_143_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_144_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_145_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_146_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_147_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_148_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_149_itm <= 1'b0;
    end
    else begin
      reg_vec_rsc_triosy_0_15_obj_ld_cse <= and_dcpl_111 & and_dcpl_97 & and_dcpl_50
          & (~ STAGE_LOOP_acc_itm_2_1);
      COMP_LOOP_nor_11_itm <= (COMP_LOOP_mux1h_428_nl & (mux_2888_nl | (fsm_output[0])))
          | (mux_2983_nl & (fsm_output[0]));
      modExp_exp_1_7_1_sva <= COMP_LOOP_mux1h_464_nl & (~ mux_3396_nl);
      COMP_LOOP_nor_12_itm <= (COMP_LOOP_mux1h_474_nl & (~(mux_3417_nl & (fsm_output[1]))))
          | (~(mux_3513_nl | (fsm_output[1])));
      COMP_LOOP_nor_134_itm <= (COMP_LOOP_mux1h_477_nl & mux_3584_nl) | mux_3591_nl;
      COMP_LOOP_nor_137_itm <= (COMP_LOOP_mux1h_479_nl & (mux_3598_nl | (fsm_output[10])))
          | mux_3605_nl;
      COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm <= COMP_LOOP_mux1h_480_nl & (~ and_dcpl_283);
      COMP_LOOP_COMP_LOOP_nor_1_itm <= ~((z_out_7[4:1]!=4'b0000));
      COMP_LOOP_COMP_LOOP_and_139_itm <= (z_out_7[4:1]==4'b0101);
      COMP_LOOP_COMP_LOOP_and_140_itm <= (z_out_7[4:1]==4'b0110);
      COMP_LOOP_COMP_LOOP_and_141_itm <= (z_out_7[4:1]==4'b0111);
      COMP_LOOP_COMP_LOOP_and_143_itm <= (z_out_7[4:1]==4'b1001);
      COMP_LOOP_COMP_LOOP_and_144_itm <= (z_out_7[4:1]==4'b1010);
      COMP_LOOP_COMP_LOOP_and_145_itm <= (z_out_7[4:1]==4'b1011);
      COMP_LOOP_COMP_LOOP_and_146_itm <= (z_out_7[4:1]==4'b1100);
      COMP_LOOP_COMP_LOOP_and_147_itm <= (z_out_7[4:1]==4'b1101);
      COMP_LOOP_COMP_LOOP_and_148_itm <= (z_out_7[4:1]==4'b1110);
      COMP_LOOP_COMP_LOOP_and_149_itm <= (z_out_7[4:1]==4'b1111);
    end
  end
  always @(posedge clk) begin
    modulo_result_rem_cmp_a <= MUX1HOT_v_64_6_2(z_out_10, operator_64_false_acc_mut_63_0,
        COMP_LOOP_10_acc_8_itm, COMP_LOOP_1_modExp_1_while_if_mul_mut_1, COMP_LOOP_10_mul_mut,
        z_out_5, {modulo_result_or_nl , (~ mux_2303_nl) , (~ mux_2378_nl) , mux_2394_nl
        , (~ mux_2461_nl) , (~ mux_2475_itm)});
    modulo_result_rem_cmp_b <= p_sva;
    operator_66_true_div_cmp_a <= MUX_v_65_2_2(z_out_6, ({operator_64_false_acc_mut_64
        , operator_64_false_acc_mut_63_0}), and_dcpl_266);
    operator_66_true_div_cmp_b_9_0 <= MUX_v_10_2_2(STAGE_LOOP_lshift_psp_sva_mx0w0,
        STAGE_LOOP_lshift_psp_sva, and_dcpl_266);
  end
  always @(posedge clk) begin
    if ( ~ mux_2495_nl ) begin
      STAGE_LOOP_lshift_psp_sva <= STAGE_LOOP_lshift_psp_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ mux_3896_nl ) begin
      operator_64_false_acc_mut_64 <= operator_64_false_mux1h_2_rgt[64];
    end
  end
  always @(posedge clk) begin
    if ( ~ mux_3949_nl ) begin
      operator_64_false_acc_mut_63_0 <= operator_64_false_mux1h_2_rgt[63:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      VEC_LOOP_j_sva_11_0 <= 12'b000000000000;
    end
    else if ( and_dcpl_273 | VEC_LOOP_j_sva_11_0_mx0c1 ) begin
      VEC_LOOP_j_sva_11_0 <= MUX_v_12_2_2(12'b000000000000, (z_out_6[11:0]), VEC_LOOP_j_sva_11_0_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_k_9_4_sva_4_0 <= 5'b00000;
    end
    else if ( ~(mux_3952_nl | (fsm_output[8])) ) begin
      COMP_LOOP_k_9_4_sva_4_0 <= MUX_v_5_2_2(5'b00000, (COMP_LOOP_k_9_4_sva_2[4:0]),
          or_3477_nl);
    end
  end
  always @(posedge clk) begin
    if ( (modExp_while_and_3 | modExp_while_and_5 | modExp_result_sva_mx0c0 | (~
        mux_2675_nl)) & (modExp_result_sva_mx0c0 | modExp_result_and_rgt | modExp_result_and_1_rgt)
        ) begin
      modExp_result_sva <= MUX1HOT_v_64_3_2(64'b0000000000000000000000000000000000000000000000000000000000000001,
          modulo_result_rem_cmp_z, (z_out_6[63:0]), {modExp_result_sva_mx0c0 , modExp_result_and_rgt
          , modExp_result_and_1_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      tmp_10_lpi_4_dfm <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( MUX_s_1_2_2((~ mux_2740_nl), mux_2705_nl, fsm_output[9]) ) begin
      tmp_10_lpi_4_dfm <= MUX1HOT_v_64_17_2(({1'b0 , operator_64_false_slc_modExp_exp_63_1_3}),
          vec_rsc_0_0_i_qa_d, vec_rsc_0_1_i_qa_d, vec_rsc_0_2_i_qa_d, vec_rsc_0_3_i_qa_d,
          vec_rsc_0_4_i_qa_d, vec_rsc_0_5_i_qa_d, vec_rsc_0_6_i_qa_d, vec_rsc_0_7_i_qa_d,
          vec_rsc_0_8_i_qa_d, vec_rsc_0_9_i_qa_d, vec_rsc_0_10_i_qa_d, vec_rsc_0_11_i_qa_d,
          vec_rsc_0_12_i_qa_d, vec_rsc_0_13_i_qa_d, vec_rsc_0_14_i_qa_d, vec_rsc_0_15_i_qa_d,
          {and_dcpl_273 , COMP_LOOP_or_8_nl , COMP_LOOP_or_9_nl , COMP_LOOP_or_10_nl
          , COMP_LOOP_or_11_nl , COMP_LOOP_or_12_nl , COMP_LOOP_or_13_nl , COMP_LOOP_or_14_nl
          , COMP_LOOP_or_15_nl , COMP_LOOP_or_16_nl , COMP_LOOP_or_17_nl , COMP_LOOP_or_18_nl
          , COMP_LOOP_or_19_nl , COMP_LOOP_or_20_nl , COMP_LOOP_or_21_nl , COMP_LOOP_or_22_nl
          , COMP_LOOP_or_23_nl});
    end
  end
  always @(posedge clk) begin
    if ( MUX_s_1_2_2(mux_2867_nl, mux_2822_nl, fsm_output[9]) ) begin
      COMP_LOOP_10_mul_mut <= MUX1HOT_v_64_21_2(r_sva, modulo_result_rem_cmp_z, (z_out_6[63:0]),
          modExp_result_sva, vec_rsc_0_0_i_qa_d, vec_rsc_0_1_i_qa_d, vec_rsc_0_2_i_qa_d,
          vec_rsc_0_3_i_qa_d, vec_rsc_0_4_i_qa_d, vec_rsc_0_5_i_qa_d, vec_rsc_0_6_i_qa_d,
          vec_rsc_0_7_i_qa_d, vec_rsc_0_8_i_qa_d, vec_rsc_0_9_i_qa_d, vec_rsc_0_10_i_qa_d,
          vec_rsc_0_11_i_qa_d, vec_rsc_0_12_i_qa_d, vec_rsc_0_13_i_qa_d, vec_rsc_0_14_i_qa_d,
          vec_rsc_0_15_i_qa_d, COMP_LOOP_1_modExp_1_while_if_mul_mut_1, {and_340_nl
          , COMP_LOOP_or_30_nl , COMP_LOOP_or_31_nl , not_tmp_596 , COMP_LOOP_and_277_nl
          , COMP_LOOP_COMP_LOOP_and_932_nl , COMP_LOOP_COMP_LOOP_and_934_nl , COMP_LOOP_and_1_nl
          , COMP_LOOP_COMP_LOOP_and_936_nl , COMP_LOOP_and_2_nl , COMP_LOOP_and_3_nl
          , COMP_LOOP_and_4_nl , COMP_LOOP_COMP_LOOP_and_930_nl , COMP_LOOP_and_5_nl
          , COMP_LOOP_and_6_nl , COMP_LOOP_and_7_nl , COMP_LOOP_and_8_nl , COMP_LOOP_and_9_nl
          , COMP_LOOP_and_10_nl , COMP_LOOP_and_11_nl , mux_114_nl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_137_itm <= 1'b0;
    end
    else if ( and_dcpl_260 | and_dcpl_332 | and_dcpl_126 | and_dcpl_141 | and_dcpl_147
        | and_dcpl_158 | and_dcpl_164 | and_dcpl_175 | and_dcpl_182 | and_dcpl_192
        | and_dcpl_198 | and_dcpl_206 | and_dcpl_217 | and_dcpl_225 | and_dcpl_232
        | and_dcpl_242 | and_dcpl_247 | and_dcpl_255 ) begin
      COMP_LOOP_COMP_LOOP_and_137_itm <= MUX1HOT_s_1_3_2((~ (z_out_5[63])), (~ (z_out_8_8_7[1])),
          COMP_LOOP_COMP_LOOP_and_17_nl, {and_dcpl_260 , and_dcpl_332 , COMP_LOOP_or_32_cse});
    end
  end
  always @(posedge clk) begin
    if ( mux_3181_nl | (~ mux_2475_itm) ) begin
      COMP_LOOP_10_acc_8_itm <= MUX_v_64_2_2(COMP_LOOP_1_acc_8_nl, z_out_10, mux_2475_itm);
    end
  end
  always @(posedge clk) begin
    if ( ~(or_tmp_9 | (~ (fsm_output[0])) | (fsm_output[6]) | (fsm_output[7]) | (~
        (fsm_output[5])) | (fsm_output[2]) | (fsm_output[8]) | (~ (fsm_output[4]))
        | (fsm_output[9])) ) begin
      COMP_LOOP_acc_psp_sva <= COMP_LOOP_acc_psp_sva_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_nor_itm <= 1'b0;
    end
    else if ( ~ not_tmp_708 ) begin
      COMP_LOOP_COMP_LOOP_nor_itm <= ~((VEC_LOOP_j_sva_11_0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_305_itm <= 1'b0;
    end
    else if ( ~ not_tmp_708 ) begin
      COMP_LOOP_COMP_LOOP_and_305_itm <= (COMP_LOOP_acc_1_cse_6_sva_1[3:0]==4'b0110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_62_itm <= 1'b0;
    end
    else if ( ~ not_tmp_708 ) begin
      COMP_LOOP_COMP_LOOP_and_62_itm <= (COMP_LOOP_acc_1_cse_2_sva_1[3:0]==4'b0011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_2_itm <= 1'b0;
    end
    else if ( ~ not_tmp_708 ) begin
      COMP_LOOP_COMP_LOOP_and_2_itm <= (VEC_LOOP_j_sva_11_0[3:0]==4'b0011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_64_itm <= 1'b0;
    end
    else if ( ~ not_tmp_708 ) begin
      COMP_LOOP_COMP_LOOP_and_64_itm <= (COMP_LOOP_acc_1_cse_2_sva_1[3:0]==4'b0101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_4_itm <= 1'b0;
    end
    else if ( ~ not_tmp_708 ) begin
      COMP_LOOP_COMP_LOOP_and_4_itm <= (VEC_LOOP_j_sva_11_0[3:0]==4'b0101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_5_itm <= 1'b0;
    end
    else if ( ~ not_tmp_708 ) begin
      COMP_LOOP_COMP_LOOP_and_5_itm <= (VEC_LOOP_j_sva_11_0[3:0]==4'b0110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_6_itm <= 1'b0;
    end
    else if ( ~ not_tmp_708 ) begin
      COMP_LOOP_COMP_LOOP_and_6_itm <= (VEC_LOOP_j_sva_11_0[3:0]==4'b0111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_68_itm <= 1'b0;
    end
    else if ( ~ not_tmp_708 ) begin
      COMP_LOOP_COMP_LOOP_and_68_itm <= (COMP_LOOP_acc_1_cse_2_sva_1[3:0]==4'b1001);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_8_itm <= 1'b0;
    end
    else if ( ~ not_tmp_708 ) begin
      COMP_LOOP_COMP_LOOP_and_8_itm <= (VEC_LOOP_j_sva_11_0[3:0]==4'b1001);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_9_itm <= 1'b0;
    end
    else if ( ~ not_tmp_708 ) begin
      COMP_LOOP_COMP_LOOP_and_9_itm <= (VEC_LOOP_j_sva_11_0[3:0]==4'b1010);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_10_itm <= 1'b0;
    end
    else if ( MUX_s_1_2_2(nor_nl, and_1253_nl, fsm_output[9]) ) begin
      COMP_LOOP_COMP_LOOP_and_10_itm <= MUX_s_1_2_2(COMP_LOOP_COMP_LOOP_and_10_nl,
          (~ (readslicef_10_1_9(COMP_LOOP_1_acc_nl))), and_dcpl_255);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_11_itm <= 1'b0;
    end
    else if ( ~ not_tmp_708 ) begin
      COMP_LOOP_COMP_LOOP_and_11_itm <= (VEC_LOOP_j_sva_11_0[3:0]==4'b1100);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_12_itm <= 1'b0;
    end
    else if ( ~ not_tmp_708 ) begin
      COMP_LOOP_COMP_LOOP_and_12_itm <= (VEC_LOOP_j_sva_11_0[3:0]==4'b1101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_13_itm <= 1'b0;
    end
    else if ( ~ not_tmp_708 ) begin
      COMP_LOOP_COMP_LOOP_and_13_itm <= (VEC_LOOP_j_sva_11_0[3:0]==4'b1110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_14_itm <= 1'b0;
    end
    else if ( ~ not_tmp_708 ) begin
      COMP_LOOP_COMP_LOOP_and_14_itm <= (VEC_LOOP_j_sva_11_0[3:0]==4'b1111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_1_cse_6_sva <= 12'b000000000000;
    end
    else if ( mux_3224_nl | (fsm_output[10]) ) begin
      COMP_LOOP_acc_1_cse_6_sva <= COMP_LOOP_acc_1_cse_6_sva_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_1_cse_2_sva <= 12'b000000000000;
    end
    else if ( mux_3234_nl | (fsm_output[10:8]!=3'b000) ) begin
      COMP_LOOP_acc_1_cse_2_sva <= COMP_LOOP_acc_1_cse_2_sva_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_11_psp_sva <= 11'b00000000000;
    end
    else if ( ~((~ mux_3242_nl) & nor_601_cse) ) begin
      COMP_LOOP_acc_11_psp_sva <= nl_COMP_LOOP_acc_11_psp_sva[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_1_cse_4_sva <= 12'b000000000000;
    end
    else if ( ~(mux_3243_nl & nor_601_cse) ) begin
      COMP_LOOP_acc_1_cse_4_sva <= z_out_5[11:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_13_psp_sva <= 10'b0000000000;
    end
    else if ( mux_3249_nl | (fsm_output[10]) ) begin
      COMP_LOOP_acc_13_psp_sva <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_14_psp_sva <= 11'b00000000000;
    end
    else if ( mux_3251_nl | (fsm_output[10]) ) begin
      COMP_LOOP_acc_14_psp_sva <= nl_COMP_LOOP_acc_14_psp_sva[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_1_cse_8_sva <= 12'b000000000000;
    end
    else if ( mux_3255_nl | (fsm_output[10]) ) begin
      COMP_LOOP_acc_1_cse_8_sva <= nl_COMP_LOOP_acc_1_cse_8_sva[11:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_16_psp_sva <= 9'b000000000;
    end
    else if ( mux_3263_nl | (fsm_output[10]) ) begin
      COMP_LOOP_acc_16_psp_sva <= z_out_7[8:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_1_cse_10_sva <= 12'b000000000000;
    end
    else if ( MUX_s_1_2_2(mux_3267_nl, mux_3264_nl, fsm_output[4]) ) begin
      COMP_LOOP_acc_1_cse_10_sva <= nl_COMP_LOOP_acc_1_cse_10_sva[11:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_17_psp_sva <= 11'b00000000000;
    end
    else if ( MUX_s_1_2_2(mux_3276_nl, (fsm_output[10]), fsm_output[9]) ) begin
      COMP_LOOP_acc_17_psp_sva <= nl_COMP_LOOP_acc_17_psp_sva[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_1_cse_12_sva <= 12'b000000000000;
    end
    else if ( MUX_s_1_2_2(mux_3288_nl, mux_3287_nl, fsm_output[4]) ) begin
      COMP_LOOP_acc_1_cse_12_sva <= nl_COMP_LOOP_acc_1_cse_12_sva[11:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_19_psp_sva <= 10'b0000000000;
    end
    else if ( MUX_s_1_2_2(mux_3292_nl, (fsm_output[10]), fsm_output[9]) ) begin
      COMP_LOOP_acc_19_psp_sva <= z_out_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_1_cse_14_sva <= 12'b000000000000;
    end
    else if ( MUX_s_1_2_2(mux_3297_nl, (fsm_output[10]), fsm_output[9]) ) begin
      COMP_LOOP_acc_1_cse_14_sva <= nl_COMP_LOOP_acc_1_cse_14_sva[11:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_20_psp_sva <= 11'b00000000000;
    end
    else if ( MUX_s_1_2_2(nor_1420_nl, and_1254_nl, fsm_output[9]) ) begin
      COMP_LOOP_acc_20_psp_sva <= nl_COMP_LOOP_acc_20_psp_sva[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_1_cse_sva <= 12'b000000000000;
    end
    else if ( MUX_s_1_2_2(mux_3304_nl, and_816_cse, or_2935_cse) ) begin
      COMP_LOOP_acc_1_cse_sva <= nl_COMP_LOOP_acc_1_cse_sva[11:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      modExp_exp_1_6_1_sva <= 1'b0;
      modExp_exp_1_5_1_sva <= 1'b0;
      modExp_exp_1_4_1_sva <= 1'b0;
    end
    else if ( mux_3369_itm ) begin
      modExp_exp_1_6_1_sva <= MUX1HOT_s_1_3_2((COMP_LOOP_k_9_4_sva_4_0[2]), modExp_exp_1_7_1_sva,
          (COMP_LOOP_k_9_4_sva_4_0[3]), {and_dcpl_283 , not_tmp_776 , not_tmp_762});
      modExp_exp_1_5_1_sva <= MUX1HOT_s_1_3_2((COMP_LOOP_k_9_4_sva_4_0[1]), modExp_exp_1_6_1_sva,
          (COMP_LOOP_k_9_4_sva_4_0[2]), {and_dcpl_283 , not_tmp_776 , not_tmp_762});
      modExp_exp_1_4_1_sva <= MUX1HOT_s_1_3_2((COMP_LOOP_k_9_4_sva_4_0[0]), modExp_exp_1_5_1_sva,
          (COMP_LOOP_k_9_4_sva_4_0[1]), {and_dcpl_283 , not_tmp_776 , not_tmp_762});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_10_cse_12_1_1_sva <= 12'b000000000000;
    end
    else if ( COMP_LOOP_or_32_cse ) begin
      COMP_LOOP_acc_10_cse_12_1_1_sva <= z_out_7[12:1];
    end
  end
  always @(posedge clk) begin
    if ( and_dcpl_126 | not_tmp_519 | and_dcpl_141 | and_dcpl_158 | and_dcpl_164
        | and_dcpl_175 | and_dcpl_192 | and_dcpl_198 | and_dcpl_206 | and_dcpl_225
        | and_dcpl_232 | and_dcpl_242 ) begin
      COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm <= MUX_s_1_2_2((z_out[9]), (z_out_8_8_7[1]),
          not_tmp_519);
    end
  end
  assign modulo_result_or_nl = and_dcpl_260 | not_tmp_519;
  assign mux_2296_nl = MUX_s_1_2_2(and_dcpl_123, (fsm_output[3]), and_573_cse);
  assign mux_2297_nl = MUX_s_1_2_2(or_tmp_2233, (~ mux_2296_nl), fsm_output[6]);
  assign mux_2298_nl = MUX_s_1_2_2(mux_2297_nl, mux_tmp_2220, fsm_output[7]);
  assign mux_2295_nl = MUX_s_1_2_2((~ and_tmp_10), mux_tmp_2218, fsm_output[7]);
  assign mux_2299_nl = MUX_s_1_2_2((~ mux_2298_nl), mux_2295_nl, fsm_output[5]);
  assign mux_2291_nl = MUX_s_1_2_2((fsm_output[3]), or_tmp_2260, fsm_output[1]);
  assign mux_2292_nl = MUX_s_1_2_2(mux_tmp_2254, mux_2291_nl, fsm_output[6]);
  assign nand_264_nl = ~((fsm_output[6]) & nor_tmp_295);
  assign mux_2293_nl = MUX_s_1_2_2(mux_2292_nl, nand_264_nl, fsm_output[7]);
  assign mux_2294_nl = MUX_s_1_2_2(mux_2293_nl, mux_tmp_2290, fsm_output[5]);
  assign mux_2300_nl = MUX_s_1_2_2(mux_2299_nl, mux_2294_nl, fsm_output[2]);
  assign mux_2286_nl = MUX_s_1_2_2(mux_tmp_2285, or_tmp_2223, fsm_output[7]);
  assign mux_2283_nl = MUX_s_1_2_2(or_tmp_2230, (~ nor_tmp_6), fsm_output[6]);
  assign mux_2282_nl = MUX_s_1_2_2(nor_tmp_295, (fsm_output[10]), fsm_output[6]);
  assign mux_2284_nl = MUX_s_1_2_2(mux_2283_nl, mux_2282_nl, fsm_output[7]);
  assign mux_2287_nl = MUX_s_1_2_2(mux_2286_nl, mux_2284_nl, fsm_output[5]);
  assign mux_2278_nl = MUX_s_1_2_2(and_dcpl_101, nor_tmp_6, fsm_output[6]);
  assign mux_2280_nl = MUX_s_1_2_2(mux_28_cse, (~ mux_2278_nl), fsm_output[7]);
  assign nand_265_nl = ~((and_574_cse | (fsm_output[3])) & (fsm_output[10]));
  assign mux_2276_nl = MUX_s_1_2_2((fsm_output[10]), or_tmp_2248, fsm_output[6]);
  assign mux_2277_nl = MUX_s_1_2_2(nand_265_nl, mux_2276_nl, fsm_output[7]);
  assign mux_2281_nl = MUX_s_1_2_2(mux_2280_nl, mux_2277_nl, fsm_output[5]);
  assign mux_2288_nl = MUX_s_1_2_2(mux_2287_nl, mux_2281_nl, fsm_output[2]);
  assign mux_2301_nl = MUX_s_1_2_2(mux_2300_nl, mux_2288_nl, fsm_output[8]);
  assign mux_2272_nl = MUX_s_1_2_2(or_tmp_14, nand_tmp_92, fsm_output[7]);
  assign mux_2270_nl = MUX_s_1_2_2((~ (fsm_output[3])), nor_tmp_6, fsm_output[6]);
  assign mux_2271_nl = MUX_s_1_2_2(mux_2270_nl, or_tmp_14, fsm_output[7]);
  assign mux_2273_nl = MUX_s_1_2_2(mux_2272_nl, mux_2271_nl, fsm_output[5]);
  assign mux_2267_nl = MUX_s_1_2_2((~ nor_tmp_291), mux_tmp_2250, fsm_output[6]);
  assign mux_2268_nl = MUX_s_1_2_2(or_tmp_2257, mux_2267_nl, fsm_output[7]);
  assign mux_2266_nl = MUX_s_1_2_2(mux_tmp_2265, or_tmp_2255, fsm_output[7]);
  assign mux_2269_nl = MUX_s_1_2_2(mux_2268_nl, mux_2266_nl, fsm_output[5]);
  assign mux_2274_nl = MUX_s_1_2_2(mux_2273_nl, mux_2269_nl, fsm_output[2]);
  assign nor_778_nl = ~((fsm_output[6]) | nor_tmp_6);
  assign mux_2261_nl = MUX_s_1_2_2(nor_tmp_9, or_tmp_2253, fsm_output[6]);
  assign mux_2262_nl = MUX_s_1_2_2(nor_778_nl, mux_2261_nl, fsm_output[7]);
  assign mux_2259_nl = MUX_s_1_2_2(or_tmp_2253, (~ mux_tmp_2251), fsm_output[6]);
  assign mux_2258_nl = MUX_s_1_2_2((~ or_tmp_2238), nor_tmp_6, fsm_output[6]);
  assign mux_2260_nl = MUX_s_1_2_2(mux_2259_nl, mux_2258_nl, fsm_output[7]);
  assign mux_2263_nl = MUX_s_1_2_2(mux_2262_nl, mux_2260_nl, fsm_output[5]);
  assign nor_779_nl = ~((fsm_output[6]) | nor_tmp_9);
  assign mux_2255_nl = MUX_s_1_2_2(or_tmp_2233, (~ mux_tmp_2254), fsm_output[6]);
  assign mux_2256_nl = MUX_s_1_2_2(nor_779_nl, mux_2255_nl, fsm_output[7]);
  assign mux_2252_nl = MUX_s_1_2_2(mux_tmp_2251, mux_tmp_2250, fsm_output[6]);
  assign mux_2253_nl = MUX_s_1_2_2((~ mux_2252_nl), and_tmp_10, fsm_output[7]);
  assign mux_2257_nl = MUX_s_1_2_2(mux_2256_nl, mux_2253_nl, fsm_output[5]);
  assign mux_2264_nl = MUX_s_1_2_2(mux_2263_nl, mux_2257_nl, fsm_output[2]);
  assign mux_2275_nl = MUX_s_1_2_2(mux_2274_nl, (~ mux_2264_nl), fsm_output[8]);
  assign mux_2302_nl = MUX_s_1_2_2(mux_2301_nl, mux_2275_nl, fsm_output[4]);
  assign mux_2245_nl = MUX_s_1_2_2(mux_tmp_2239, nor_tmp_6, fsm_output[6]);
  assign or_2306_nl = (fsm_output[7]) | mux_2245_nl;
  assign mux_2244_nl = MUX_s_1_2_2(not_tmp_426, or_tmp_2246, fsm_output[7]);
  assign mux_2246_nl = MUX_s_1_2_2(or_2306_nl, mux_2244_nl, fsm_output[5]);
  assign mux_2242_nl = MUX_s_1_2_2(nor_tmp_286, or_tmp_2237, fsm_output[7]);
  assign mux_2241_nl = MUX_s_1_2_2(nand_tmp_92, or_tmp_14, fsm_output[7]);
  assign mux_2243_nl = MUX_s_1_2_2(mux_2242_nl, mux_2241_nl, fsm_output[5]);
  assign mux_2247_nl = MUX_s_1_2_2(mux_2246_nl, mux_2243_nl, fsm_output[2]);
  assign mux_2235_nl = MUX_s_1_2_2(or_tmp_2220, or_tmp_21, fsm_output[6]);
  assign or_2300_nl = (fsm_output[6]) | (fsm_output[0]) | (fsm_output[1]) | (fsm_output[3])
      | (fsm_output[10]);
  assign mux_2236_nl = MUX_s_1_2_2(mux_2235_nl, or_2300_nl, fsm_output[7]);
  assign nand_91_nl = ~((fsm_output[7]) & (~((((fsm_output[6]) | (fsm_output[1]))
      & (fsm_output[3])) | (fsm_output[10]))));
  assign mux_2237_nl = MUX_s_1_2_2(mux_2236_nl, nand_91_nl, fsm_output[5]);
  assign mux_2233_nl = MUX_s_1_2_2(or_tmp_237, or_tmp_2238, fsm_output[6]);
  assign or_2297_nl = (fsm_output[7]) | mux_2233_nl;
  assign or_2293_nl = ((fsm_output[6]) & (fsm_output[1])) | (fsm_output[3]) | (fsm_output[10]);
  assign mux_2232_nl = MUX_s_1_2_2(or_tmp_2237, or_2293_nl, fsm_output[7]);
  assign mux_2234_nl = MUX_s_1_2_2(or_2297_nl, mux_2232_nl, fsm_output[5]);
  assign mux_2238_nl = MUX_s_1_2_2(mux_2237_nl, mux_2234_nl, fsm_output[2]);
  assign mux_2248_nl = MUX_s_1_2_2(mux_2247_nl, mux_2238_nl, fsm_output[8]);
  assign mux_2225_nl = MUX_s_1_2_2(and_dcpl_101, nor_tmp_6, fsm_output[1]);
  assign mux_2226_nl = MUX_s_1_2_2(and_dcpl_102, mux_2225_nl, fsm_output[0]);
  assign mux_2227_nl = MUX_s_1_2_2(and_dcpl_101, mux_2226_nl, fsm_output[6]);
  assign mux_2228_nl = MUX_s_1_2_2((~ mux_2227_nl), or_tmp_4, fsm_output[7]);
  assign mux_2224_nl = MUX_s_1_2_2(mux_tmp_2223, or_tmp_2223, fsm_output[7]);
  assign mux_2229_nl = MUX_s_1_2_2(mux_2228_nl, mux_2224_nl, fsm_output[5]);
  assign mux_2221_nl = MUX_s_1_2_2((~ mux_tmp_2220), or_tmp_4, fsm_output[7]);
  assign or_2288_nl = (fsm_output[6]) | or_tmp_2230;
  assign mux_2219_nl = MUX_s_1_2_2(mux_tmp_2218, or_2288_nl, fsm_output[7]);
  assign mux_2222_nl = MUX_s_1_2_2(mux_2221_nl, mux_2219_nl, fsm_output[5]);
  assign mux_2230_nl = MUX_s_1_2_2(mux_2229_nl, mux_2222_nl, fsm_output[2]);
  assign or_2285_nl = (~(and_574_cse | (fsm_output[3]))) | (fsm_output[10]);
  assign mux_2215_nl = MUX_s_1_2_2(or_tmp_14, or_2285_nl, fsm_output[7]);
  assign mux_2214_nl = MUX_s_1_2_2(or_tmp_2225, (fsm_output[10]), fsm_output[6]);
  assign or_2283_nl = (fsm_output[7]) | mux_2214_nl;
  assign mux_2216_nl = MUX_s_1_2_2(mux_2215_nl, or_2283_nl, fsm_output[5]);
  assign or_2279_nl = (~((fsm_output[3]) | (fsm_output[6]))) | (fsm_output[10]);
  assign mux_2212_nl = MUX_s_1_2_2(or_tmp_2223, or_2279_nl, fsm_output[7]);
  assign nand_90_nl = ~((fsm_output[6]) & (~ or_tmp_2220));
  assign mux_2211_nl = MUX_s_1_2_2((fsm_output[10]), nand_90_nl, fsm_output[7]);
  assign mux_2213_nl = MUX_s_1_2_2(mux_2212_nl, mux_2211_nl, fsm_output[5]);
  assign mux_2217_nl = MUX_s_1_2_2(mux_2216_nl, mux_2213_nl, fsm_output[2]);
  assign mux_2231_nl = MUX_s_1_2_2(mux_2230_nl, mux_2217_nl, fsm_output[8]);
  assign mux_2249_nl = MUX_s_1_2_2(mux_2248_nl, mux_2231_nl, fsm_output[4]);
  assign mux_2303_nl = MUX_s_1_2_2(mux_2302_nl, mux_2249_nl, fsm_output[9]);
  assign or_2355_nl = (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[10]);
  assign mux_2373_nl = MUX_s_1_2_2(or_2355_nl, or_tmp_2267, fsm_output[7]);
  assign mux_2372_nl = MUX_s_1_2_2(or_tmp_2281, (~ mux_tmp_2218), fsm_output[7]);
  assign mux_2374_nl = MUX_s_1_2_2(mux_2373_nl, mux_2372_nl, fsm_output[5]);
  assign mux_2369_nl = MUX_s_1_2_2((~ nor_tmp_300), or_tmp_2271, fsm_output[6]);
  assign or_2354_nl = (fsm_output[6]) | ((fsm_output[0]) & (fsm_output[1]) & (~ (fsm_output[3]))
      & (fsm_output[10]));
  assign mux_2370_nl = MUX_s_1_2_2(mux_2369_nl, or_2354_nl, fsm_output[7]);
  assign or_2351_nl = (fsm_output[6]) | and_dcpl_223;
  assign mux_2367_nl = MUX_s_1_2_2(or_tmp_21, mux_tmp_2362, fsm_output[6]);
  assign mux_2368_nl = MUX_s_1_2_2(or_2351_nl, mux_2367_nl, fsm_output[7]);
  assign mux_2371_nl = MUX_s_1_2_2(mux_2370_nl, mux_2368_nl, fsm_output[5]);
  assign mux_2375_nl = MUX_s_1_2_2(mux_2374_nl, mux_2371_nl, fsm_output[2]);
  assign mux_2364_nl = MUX_s_1_2_2(mux_tmp_2285, (fsm_output[6]), fsm_output[7]);
  assign nand_100_nl = ~((fsm_output[6]) & (~ mux_tmp_2362));
  assign mux_2363_nl = MUX_s_1_2_2(nand_100_nl, or_tmp_2293, fsm_output[7]);
  assign mux_2365_nl = MUX_s_1_2_2((~ mux_2364_nl), mux_2363_nl, fsm_output[5]);
  assign nand_99_nl = ~((fsm_output[6]) & (~ mux_tmp_2239));
  assign mux_2360_nl = MUX_s_1_2_2((~ mux_28_cse), nand_99_nl, fsm_output[7]);
  assign nand_98_nl = ~((fsm_output[6]) & (~ nor_tmp_295));
  assign mux_2359_nl = MUX_s_1_2_2(nand_98_nl, or_tmp_434, fsm_output[7]);
  assign mux_2361_nl = MUX_s_1_2_2(mux_2360_nl, mux_2359_nl, fsm_output[5]);
  assign mux_2366_nl = MUX_s_1_2_2(mux_2365_nl, mux_2361_nl, fsm_output[2]);
  assign mux_2376_nl = MUX_s_1_2_2(mux_2375_nl, mux_2366_nl, fsm_output[8]);
  assign mux_2354_nl = MUX_s_1_2_2((fsm_output[10]), (~ or_tmp_2248), fsm_output[6]);
  assign mux_2355_nl = MUX_s_1_2_2(mux_2354_nl, mux_tmp_2327, fsm_output[7]);
  assign mux_2352_nl = MUX_s_1_2_2(and_dcpl_109, nor_tmp_6, fsm_output[6]);
  assign mux_2353_nl = MUX_s_1_2_2(mux_2352_nl, and_tmp_16, fsm_output[7]);
  assign mux_2356_nl = MUX_s_1_2_2(mux_2355_nl, mux_2353_nl, fsm_output[5]);
  assign nand_261_nl = ~(or_2348_cse & mux_tmp_2239);
  assign mux_2348_nl = MUX_s_1_2_2(nand_261_nl, nor_tmp_6, fsm_output[6]);
  assign mux_2350_nl = MUX_s_1_2_2((~ mux_tmp_2349), mux_2348_nl, fsm_output[7]);
  assign and_275_nl = (fsm_output[6]) & ((fsm_output[1]) | (~ (fsm_output[3])) |
      (fsm_output[10]));
  assign mux_2347_nl = MUX_s_1_2_2(mux_tmp_2265, and_275_nl, fsm_output[7]);
  assign mux_2351_nl = MUX_s_1_2_2(mux_2350_nl, mux_2347_nl, fsm_output[5]);
  assign mux_2357_nl = MUX_s_1_2_2(mux_2356_nl, mux_2351_nl, fsm_output[2]);
  assign mux_2344_nl = MUX_s_1_2_2(not_tmp_463, nand_tmp_96, fsm_output[7]);
  assign or_2342_nl = (fsm_output[1]) | (~ nor_tmp_6);
  assign mux_2342_nl = MUX_s_1_2_2(or_tmp_2266, or_2342_nl, fsm_output[0]);
  assign or_2343_nl = (fsm_output[6]) | (~ mux_2342_nl);
  assign mux_2343_nl = MUX_s_1_2_2(or_tmp_3, or_2343_nl, fsm_output[7]);
  assign mux_2345_nl = MUX_s_1_2_2(mux_2344_nl, mux_2343_nl, fsm_output[5]);
  assign or_2341_nl = (fsm_output[1]) | (fsm_output[3]) | (~ (fsm_output[10]));
  assign mux_2339_nl = MUX_s_1_2_2(or_2341_nl, or_tmp_2282, fsm_output[0]);
  assign nand_262_nl = ~((fsm_output[6]) & mux_2339_nl);
  assign mux_2340_nl = MUX_s_1_2_2(nand_262_nl, or_tmp_3, fsm_output[7]);
  assign mux_2337_nl = MUX_s_1_2_2((~ and_dcpl_240), or_tmp_2238, fsm_output[6]);
  assign mux_2338_nl = MUX_s_1_2_2(mux_2337_nl, or_tmp_2281, fsm_output[7]);
  assign mux_2341_nl = MUX_s_1_2_2(mux_2340_nl, mux_2338_nl, fsm_output[5]);
  assign mux_2346_nl = MUX_s_1_2_2(mux_2345_nl, mux_2341_nl, fsm_output[2]);
  assign mux_2358_nl = MUX_s_1_2_2((~ mux_2357_nl), mux_2346_nl, fsm_output[8]);
  assign mux_2377_nl = MUX_s_1_2_2(mux_2376_nl, mux_2358_nl, fsm_output[4]);
  assign mux_2332_nl = MUX_s_1_2_2(or_36_cse, or_tmp_14, fsm_output[7]);
  assign mux_2331_nl = MUX_s_1_2_2(or_tmp_2280, or_15_cse, fsm_output[7]);
  assign mux_2333_nl = MUX_s_1_2_2(mux_2332_nl, mux_2331_nl, fsm_output[5]);
  assign mux_2329_nl = MUX_s_1_2_2(or_36_cse, or_tmp_2255, fsm_output[7]);
  assign mux_2328_nl = MUX_s_1_2_2((~ mux_tmp_2327), or_tmp_4, fsm_output[7]);
  assign mux_2330_nl = MUX_s_1_2_2(mux_2329_nl, mux_2328_nl, fsm_output[5]);
  assign mux_2334_nl = MUX_s_1_2_2(mux_2333_nl, mux_2330_nl, fsm_output[2]);
  assign mux_2323_nl = MUX_s_1_2_2(or_tmp_2248, or_tmp_237, fsm_output[6]);
  assign nand_97_nl = ~((fsm_output[6]) & (~ or_tmp_2275));
  assign mux_2324_nl = MUX_s_1_2_2(mux_2323_nl, nand_97_nl, fsm_output[7]);
  assign mux_2322_nl = MUX_s_1_2_2(or_tmp_4, or_tmp_2276, fsm_output[7]);
  assign mux_2325_nl = MUX_s_1_2_2(mux_2324_nl, mux_2322_nl, fsm_output[5]);
  assign mux_2319_nl = MUX_s_1_2_2(or_tmp_21, or_tmp_2275, fsm_output[6]);
  assign mux_2320_nl = MUX_s_1_2_2(mux_2319_nl, or_tmp_4, fsm_output[7]);
  assign mux_2318_nl = MUX_s_1_2_2(nand_tmp_96, or_tmp_2246, fsm_output[7]);
  assign mux_2321_nl = MUX_s_1_2_2(mux_2320_nl, mux_2318_nl, fsm_output[5]);
  assign mux_2326_nl = MUX_s_1_2_2(mux_2325_nl, mux_2321_nl, fsm_output[2]);
  assign mux_2335_nl = MUX_s_1_2_2(mux_2334_nl, mux_2326_nl, fsm_output[8]);
  assign or_2330_nl = (fsm_output[6]) | mux_tmp_2254;
  assign or_2329_nl = (fsm_output[6]) | or_tmp_2271;
  assign mux_2314_nl = MUX_s_1_2_2(or_2330_nl, or_2329_nl, fsm_output[7]);
  assign mux_2313_nl = MUX_s_1_2_2((~ mux_tmp_2223), nand_tmp_95, fsm_output[7]);
  assign mux_2315_nl = MUX_s_1_2_2(mux_2314_nl, mux_2313_nl, fsm_output[5]);
  assign mux_2311_nl = MUX_s_1_2_2(or_tmp_2267, or_tmp_14, fsm_output[7]);
  assign nand_94_nl = ~((fsm_output[6]) & (~ or_tmp_2225));
  assign mux_2308_nl = MUX_s_1_2_2((~ mux_tmp_2218), nand_94_nl, fsm_output[7]);
  assign mux_2312_nl = MUX_s_1_2_2(mux_2311_nl, mux_2308_nl, fsm_output[5]);
  assign mux_2316_nl = MUX_s_1_2_2(mux_2315_nl, mux_2312_nl, fsm_output[2]);
  assign mux_2305_nl = MUX_s_1_2_2(or_tmp_3, nand_tmp_93, fsm_output[7]);
  assign or_2321_nl = (~ (fsm_output[7])) | (fsm_output[6]) | (fsm_output[10]);
  assign mux_2306_nl = MUX_s_1_2_2(mux_2305_nl, or_2321_nl, fsm_output[5]);
  assign or_2319_nl = (fsm_output[7:6]!=2'b10) | or_tmp_2248;
  assign mux_2304_nl = MUX_s_1_2_2(or_tmp_2263, or_2319_nl, fsm_output[5]);
  assign mux_2307_nl = MUX_s_1_2_2(mux_2306_nl, mux_2304_nl, fsm_output[2]);
  assign mux_2317_nl = MUX_s_1_2_2(mux_2316_nl, mux_2307_nl, fsm_output[8]);
  assign mux_2336_nl = MUX_s_1_2_2(mux_2335_nl, mux_2317_nl, fsm_output[4]);
  assign mux_2378_nl = MUX_s_1_2_2(mux_2377_nl, mux_2336_nl, fsm_output[9]);
  assign nor_758_nl = ~((~ (fsm_output[7])) | (~ (fsm_output[8])) | (~ (fsm_output[2]))
      | (fsm_output[3]) | (~ (fsm_output[9])) | (fsm_output[5]) | (fsm_output[10]));
  assign nor_759_nl = ~((fsm_output[7]) | (~ (fsm_output[8])) | (fsm_output[2]) |
      (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[5]) | (~ (fsm_output[10])));
  assign mux_2391_nl = MUX_s_1_2_2(nor_758_nl, nor_759_nl, fsm_output[4]);
  assign nor_760_nl = ~((fsm_output[8]) | (~ (fsm_output[2])) | (~ (fsm_output[3]))
      | (fsm_output[9]) | (fsm_output[5]) | (fsm_output[10]));
  assign nor_761_nl = ~((~ (fsm_output[8])) | (fsm_output[2]) | (fsm_output[3]) |
      (fsm_output[9]) | (~ (fsm_output[5])) | (fsm_output[10]));
  assign mux_2390_nl = MUX_s_1_2_2(nor_760_nl, nor_761_nl, fsm_output[7]);
  assign and_568_nl = (fsm_output[4]) & mux_2390_nl;
  assign mux_2392_nl = MUX_s_1_2_2(mux_2391_nl, and_568_nl, fsm_output[6]);
  assign nor_762_nl = ~((fsm_output[7]) | (~ (fsm_output[8])) | (~ (fsm_output[2]))
      | (fsm_output[3]) | (fsm_output[9]) | (~ (fsm_output[5])) | (fsm_output[10]));
  assign nor_763_nl = ~((~ (fsm_output[7])) | (fsm_output[8]) | (fsm_output[2]) |
      (~ (fsm_output[3])) | (~ (fsm_output[9])) | (~ (fsm_output[5])) | (fsm_output[10]));
  assign mux_2388_nl = MUX_s_1_2_2(nor_762_nl, nor_763_nl, fsm_output[4]);
  assign or_2372_nl = (fsm_output[8]) | (~ (fsm_output[2])) | (~ (fsm_output[3]))
      | (fsm_output[9]) | (fsm_output[5]) | (~ (fsm_output[10]));
  assign or_2370_nl = (~ (fsm_output[8])) | (fsm_output[2]) | (fsm_output[3]) | (fsm_output[9])
      | not_tmp_45;
  assign mux_2387_nl = MUX_s_1_2_2(or_2372_nl, or_2370_nl, fsm_output[7]);
  assign nor_764_nl = ~((fsm_output[4]) | mux_2387_nl);
  assign mux_2389_nl = MUX_s_1_2_2(mux_2388_nl, nor_764_nl, fsm_output[6]);
  assign mux_2393_nl = MUX_s_1_2_2(mux_2392_nl, mux_2389_nl, fsm_output[1]);
  assign nor_765_nl = ~((fsm_output[2]) | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[5])
      | (fsm_output[10]));
  assign nor_766_nl = ~((fsm_output[2]) | (~ (fsm_output[3])) | (~ (fsm_output[9]))
      | (~ (fsm_output[5])) | (fsm_output[10]));
  assign mux_2384_nl = MUX_s_1_2_2(nor_765_nl, nor_766_nl, fsm_output[8]);
  assign and_570_nl = (fsm_output[7]) & mux_2384_nl;
  assign or_2365_nl = (~ (fsm_output[2])) | (fsm_output[3]) | (~ (fsm_output[9]))
      | (fsm_output[5]) | (fsm_output[10]);
  assign or_2364_nl = (~ (fsm_output[2])) | (~ (fsm_output[3])) | (fsm_output[9])
      | not_tmp_45;
  assign mux_2383_nl = MUX_s_1_2_2(or_2365_nl, or_2364_nl, fsm_output[8]);
  assign nor_767_nl = ~((fsm_output[7]) | mux_2383_nl);
  assign mux_2385_nl = MUX_s_1_2_2(and_570_nl, nor_767_nl, fsm_output[4]);
  assign and_569_nl = (fsm_output[6]) & mux_2385_nl;
  assign nor_768_nl = ~((~ (fsm_output[7])) | (~ (fsm_output[8])) | (fsm_output[2])
      | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[5]) | (fsm_output[10]));
  assign nor_769_nl = ~((fsm_output[2]) | (fsm_output[3]) | (fsm_output[9]) | (~
      (fsm_output[5])) | (fsm_output[10]));
  assign nor_770_nl = ~((~ (fsm_output[2])) | (~ (fsm_output[3])) | (~ (fsm_output[9]))
      | (fsm_output[5]) | (fsm_output[10]));
  assign mux_2379_nl = MUX_s_1_2_2(nor_769_nl, nor_770_nl, fsm_output[8]);
  assign nor_771_nl = ~((fsm_output[8]) | (fsm_output[2]) | (fsm_output[3]) | (fsm_output[9])
      | not_tmp_45);
  assign mux_2380_nl = MUX_s_1_2_2(mux_2379_nl, nor_771_nl, fsm_output[7]);
  assign mux_2381_nl = MUX_s_1_2_2(nor_768_nl, mux_2380_nl, fsm_output[4]);
  assign nor_772_nl = ~((fsm_output[4]) | (fsm_output[7]) | (fsm_output[8]) | (~
      (fsm_output[2])) | (fsm_output[3]) | (~ (fsm_output[9])) | (fsm_output[5])
      | (~ (fsm_output[10])));
  assign mux_2382_nl = MUX_s_1_2_2(mux_2381_nl, nor_772_nl, fsm_output[6]);
  assign mux_2386_nl = MUX_s_1_2_2(and_569_nl, mux_2382_nl, fsm_output[1]);
  assign mux_2394_nl = MUX_s_1_2_2(mux_2393_nl, mux_2386_nl, fsm_output[0]);
  assign nand_109_nl = ~((fsm_output[5]) & (~ mux_tmp_2425));
  assign mux_2456_nl = MUX_s_1_2_2(nand_109_nl, nand_tmp_108, or_2348_cse);
  assign mux_2455_nl = MUX_s_1_2_2(nand_tmp_108, nand_tmp_107, and_573_cse);
  assign mux_2457_nl = MUX_s_1_2_2(mux_2456_nl, mux_2455_nl, fsm_output[2]);
  assign mux_2452_nl = MUX_s_1_2_2((~ or_tmp_2342), mux_tmp_2426, fsm_output[0]);
  assign mux_2453_nl = MUX_s_1_2_2((~ or_tmp_2343), mux_2452_nl, fsm_output[1]);
  assign mux_2451_nl = MUX_s_1_2_2(mux_tmp_2426, mux_tmp_2436, fsm_output[1]);
  assign mux_2454_nl = MUX_s_1_2_2(mux_2453_nl, mux_2451_nl, fsm_output[2]);
  assign mux_2458_nl = MUX_s_1_2_2(mux_2457_nl, (~ mux_2454_nl), fsm_output[7]);
  assign mux_2447_nl = MUX_s_1_2_2(mux_tmp_2401, (~ nor_tmp_307), fsm_output[5]);
  assign mux_2446_nl = MUX_s_1_2_2(mux_tmp_2401, nand_257_cse, fsm_output[5]);
  assign mux_2448_nl = MUX_s_1_2_2(mux_2447_nl, mux_2446_nl, or_2348_cse);
  assign mux_2443_nl = MUX_s_1_2_2(or_tmp_434, (~ (fsm_output[6])), fsm_output[8]);
  assign mux_2444_nl = MUX_s_1_2_2(or_tmp_2334, mux_2443_nl, fsm_output[5]);
  assign mux_2445_nl = MUX_s_1_2_2(mux_2444_nl, mux_tmp_2423, or_2348_cse);
  assign mux_2449_nl = MUX_s_1_2_2(mux_2448_nl, mux_2445_nl, fsm_output[2]);
  assign mux_2450_nl = MUX_s_1_2_2(mux_tmp_2406, mux_2449_nl, fsm_output[7]);
  assign mux_2459_nl = MUX_s_1_2_2(mux_2458_nl, mux_2450_nl, fsm_output[4]);
  assign mux_2439_nl = MUX_s_1_2_2(nand_tmp_107, nand_tmp_105, and_573_cse);
  assign mux_2438_nl = MUX_s_1_2_2(nand_tmp_105, mux_tmp_2406, and_573_cse);
  assign mux_2440_nl = MUX_s_1_2_2(mux_2439_nl, mux_2438_nl, fsm_output[2]);
  assign mux_2434_nl = MUX_s_1_2_2((~ mux_2433_itm), nor_tmp_307, fsm_output[5]);
  assign mux_2437_nl = MUX_s_1_2_2(mux_tmp_2436, mux_2434_nl, fsm_output[2]);
  assign mux_2441_nl = MUX_s_1_2_2(mux_2440_nl, (~ mux_2437_nl), fsm_output[7]);
  assign mux_2430_nl = MUX_s_1_2_2(mux_tmp_2406, or_tmp_2343, or_2348_cse);
  assign mux_2428_nl = MUX_s_1_2_2(or_tmp_2343, or_tmp_2342, fsm_output[0]);
  assign mux_2429_nl = MUX_s_1_2_2(mux_2428_nl, (~ mux_tmp_2426), fsm_output[1]);
  assign mux_2431_nl = MUX_s_1_2_2(mux_2430_nl, mux_2429_nl, fsm_output[2]);
  assign nand_106_nl = ~((fsm_output[5]) & (~ mux_tmp_917));
  assign mux_2424_nl = MUX_s_1_2_2(mux_tmp_2423, nand_106_nl, and_563_cse);
  assign mux_2432_nl = MUX_s_1_2_2(mux_2431_nl, mux_2424_nl, fsm_output[7]);
  assign mux_2442_nl = MUX_s_1_2_2(mux_2441_nl, mux_2432_nl, fsm_output[4]);
  assign mux_2460_nl = MUX_s_1_2_2(mux_2459_nl, mux_2442_nl, fsm_output[3]);
  assign or_2397_nl = (fsm_output[8]) | (fsm_output[6]) | (fsm_output[10]);
  assign mux_2416_nl = MUX_s_1_2_2(or_2397_nl, mux_tmp_2401, fsm_output[5]);
  assign mux_2417_nl = MUX_s_1_2_2(mux_2416_nl, nand_tmp_105, and_573_cse);
  assign mux_2418_nl = MUX_s_1_2_2(mux_2417_nl, nand_tmp_105, fsm_output[2]);
  assign mux_2414_nl = MUX_s_1_2_2(or_tmp_2329, or_tmp_2335, or_2348_cse);
  assign mux_2415_nl = MUX_s_1_2_2(or_tmp_2329, mux_2414_nl, fsm_output[2]);
  assign mux_2419_nl = MUX_s_1_2_2(mux_2418_nl, mux_2415_nl, fsm_output[7]);
  assign mux_2411_nl = MUX_s_1_2_2(mux_tmp_2406, or_tmp_2338, fsm_output[1]);
  assign mux_2410_nl = MUX_s_1_2_2(or_tmp_2338, or_tmp_2331, fsm_output[1]);
  assign mux_2412_nl = MUX_s_1_2_2(mux_2411_nl, mux_2410_nl, fsm_output[2]);
  assign mux_2409_nl = MUX_s_1_2_2(mux_tmp_2400, or_tmp_2327, and_565_cse);
  assign mux_2413_nl = MUX_s_1_2_2(mux_2412_nl, mux_2409_nl, fsm_output[7]);
  assign mux_2420_nl = MUX_s_1_2_2(mux_2419_nl, mux_2413_nl, fsm_output[4]);
  assign mux_2404_nl = MUX_s_1_2_2(or_tmp_2335, mux_tmp_2402, fsm_output[1]);
  assign mux_2403_nl = MUX_s_1_2_2(mux_tmp_2402, mux_tmp_2400, or_2348_cse);
  assign mux_2405_nl = MUX_s_1_2_2(mux_2404_nl, mux_2403_nl, fsm_output[2]);
  assign mux_2407_nl = MUX_s_1_2_2(mux_tmp_2406, mux_2405_nl, fsm_output[7]);
  assign mux_2398_nl = MUX_s_1_2_2(or_tmp_2331, or_tmp_2329, or_2385_cse);
  assign mux_2395_nl = MUX_s_1_2_2(or_tmp_14, or_tmp_4, fsm_output[8]);
  assign nand_104_nl = ~((fsm_output[5]) & (~ mux_2395_nl));
  assign mux_2396_nl = MUX_s_1_2_2(or_tmp_2327, nand_104_nl, and_573_cse);
  assign or_2381_nl = (~ (fsm_output[5])) | (fsm_output[8]) | (fsm_output[6]) | (fsm_output[10]);
  assign mux_2397_nl = MUX_s_1_2_2(mux_2396_nl, or_2381_nl, fsm_output[2]);
  assign mux_2399_nl = MUX_s_1_2_2(mux_2398_nl, mux_2397_nl, fsm_output[7]);
  assign mux_2408_nl = MUX_s_1_2_2(mux_2407_nl, mux_2399_nl, fsm_output[4]);
  assign mux_2421_nl = MUX_s_1_2_2(mux_2420_nl, mux_2408_nl, fsm_output[3]);
  assign mux_2461_nl = MUX_s_1_2_2(mux_2460_nl, mux_2421_nl, fsm_output[9]);
  assign COMP_LOOP_nor_11_nl = ~((z_out_7[4:2]!=3'b000));
  assign COMP_LOOP_and_274_nl = (~ and_dcpl_281) & and_dcpl_273;
  assign or_2728_nl = (fsm_output[8]) | ((fsm_output[4]) & or_tmp_187);
  assign mux_2971_nl = MUX_s_1_2_2(or_2729_cse, or_2728_nl, fsm_output[1]);
  assign mux_2972_nl = MUX_s_1_2_2(mux_tmp_413, mux_2971_nl, fsm_output[6]);
  assign mux_2969_nl = MUX_s_1_2_2(mux_tmp_2930, mux_tmp_2907, or_2348_cse);
  assign mux_2970_nl = MUX_s_1_2_2(mux_2969_nl, nand_tmp_140, fsm_output[6]);
  assign mux_2973_nl = MUX_s_1_2_2(mux_2972_nl, mux_2970_nl, fsm_output[7]);
  assign mux_2965_nl = MUX_s_1_2_2((~ mux_tmp_2911), or_tmp_182, fsm_output[8]);
  assign mux_2966_nl = MUX_s_1_2_2(mux_2965_nl, or_tmp_2663, and_573_cse);
  assign mux_2964_nl = MUX_s_1_2_2(nand_tmp_140, nand_tmp_13, fsm_output[1]);
  assign mux_2967_nl = MUX_s_1_2_2(mux_2966_nl, mux_2964_nl, fsm_output[6]);
  assign mux_2963_nl = MUX_s_1_2_2(or_tmp_189, mux_tmp_2930, fsm_output[6]);
  assign mux_2968_nl = MUX_s_1_2_2(mux_2967_nl, mux_2963_nl, fsm_output[7]);
  assign mux_2974_nl = MUX_s_1_2_2(mux_2973_nl, mux_2968_nl, fsm_output[5]);
  assign mux_426_nl = MUX_s_1_2_2(or_tmp_187, nor_tmp_46, fsm_output[8]);
  assign mux_427_nl = MUX_s_1_2_2(mux_tmp_412, mux_426_nl, fsm_output[1]);
  assign mux_2956_nl = MUX_s_1_2_2(mux_tmp_2912, mux_tmp_2919, fsm_output[1]);
  assign mux_2957_nl = MUX_s_1_2_2(mux_tmp_2913, mux_2956_nl, fsm_output[0]);
  assign mux_2960_nl = MUX_s_1_2_2(mux_427_nl, mux_2957_nl, fsm_output[6]);
  assign mux_2955_nl = MUX_s_1_2_2(mux_tmp_2905, nand_tmp_13, fsm_output[6]);
  assign mux_2961_nl = MUX_s_1_2_2(mux_2960_nl, mux_2955_nl, fsm_output[7]);
  assign mux_421_nl = MUX_s_1_2_2(nand_tmp_13, nand_tmp_12, fsm_output[1]);
  assign mux_422_nl = MUX_s_1_2_2(or_tmp_191, mux_421_nl, fsm_output[6]);
  assign mux_2950_nl = MUX_s_1_2_2(or_tmp_2659, mux_tmp_2912, or_2348_cse);
  assign mux_2951_nl = MUX_s_1_2_2(mux_2950_nl, mux_tmp_2907, fsm_output[6]);
  assign mux_2954_nl = MUX_s_1_2_2(mux_422_nl, mux_2951_nl, fsm_output[7]);
  assign mux_2962_nl = MUX_s_1_2_2(mux_2961_nl, mux_2954_nl, fsm_output[5]);
  assign mux_2975_nl = MUX_s_1_2_2(mux_2974_nl, mux_2962_nl, fsm_output[3]);
  assign mux_414_nl = MUX_s_1_2_2(mux_tmp_413, mux_tmp_412, or_2348_cse);
  assign mux_2940_nl = MUX_s_1_2_2(mux_726_cse, or_tmp_187, fsm_output[4]);
  assign mux_2941_nl = MUX_s_1_2_2(mux_2940_nl, or_tmp_2652, fsm_output[8]);
  assign mux_2942_nl = MUX_s_1_2_2(mux_tmp_2912, mux_2941_nl, nor_412_cse);
  assign mux_2946_nl = MUX_s_1_2_2(mux_414_nl, mux_2942_nl, fsm_output[6]);
  assign mux_2938_nl = MUX_s_1_2_2(nand_tmp_140, nand_tmp_13, and_573_cse);
  assign mux_2939_nl = MUX_s_1_2_2(mux_tmp_2907, mux_2938_nl, fsm_output[6]);
  assign mux_2947_nl = MUX_s_1_2_2(mux_2946_nl, mux_2939_nl, fsm_output[7]);
  assign mux_2934_nl = MUX_s_1_2_2(or_tmp_2663, or_tmp_191, or_2348_cse);
  assign mux_2935_nl = MUX_s_1_2_2(mux_2934_nl, nand_tmp_13, fsm_output[6]);
  assign mux_2932_nl = MUX_s_1_2_2(or_tmp_189, or_tmp_2659, and_573_cse);
  assign mux_2931_nl = MUX_s_1_2_2(mux_tmp_2930, mux_tmp_2907, fsm_output[1]);
  assign mux_2933_nl = MUX_s_1_2_2(mux_2932_nl, mux_2931_nl, fsm_output[6]);
  assign mux_2936_nl = MUX_s_1_2_2(mux_2935_nl, mux_2933_nl, fsm_output[7]);
  assign mux_2948_nl = MUX_s_1_2_2(mux_2947_nl, mux_2936_nl, fsm_output[5]);
  assign or_2718_nl = (~ (fsm_output[8])) | (fsm_output[4]);
  assign mux_2924_nl = MUX_s_1_2_2(and_816_cse, or_tmp_187, or_2718_nl);
  assign mux_2925_nl = MUX_s_1_2_2(mux_2924_nl, mux_tmp_2921, fsm_output[1]);
  assign mux_2922_nl = MUX_s_1_2_2(or_tmp_182, mux_tmp_2911, fsm_output[8]);
  assign mux_2923_nl = MUX_s_1_2_2(mux_2922_nl, mux_tmp_2921, fsm_output[1]);
  assign mux_2926_nl = MUX_s_1_2_2(mux_2925_nl, mux_2923_nl, fsm_output[0]);
  assign mux_2927_nl = MUX_s_1_2_2(mux_2926_nl, mux_tmp_2919, fsm_output[6]);
  assign mux_386_nl = MUX_s_1_2_2(nand_tmp_13, nand_tmp_12, and_573_cse);
  assign mux_2918_nl = MUX_s_1_2_2(or_tmp_2649, mux_386_nl, fsm_output[6]);
  assign mux_2928_nl = MUX_s_1_2_2(mux_2927_nl, mux_2918_nl, fsm_output[7]);
  assign mux_2908_nl = MUX_s_1_2_2(mux_tmp_2907, nand_tmp_136, fsm_output[1]);
  assign mux_2909_nl = MUX_s_1_2_2(mux_2908_nl, mux_tmp_2905, fsm_output[0]);
  assign mux_2914_nl = MUX_s_1_2_2(mux_tmp_2913, mux_2909_nl, fsm_output[6]);
  assign mux_2916_nl = MUX_s_1_2_2(mux_384_cse, mux_2914_nl, fsm_output[7]);
  assign mux_2929_nl = MUX_s_1_2_2(mux_2928_nl, mux_2916_nl, fsm_output[5]);
  assign mux_2949_nl = MUX_s_1_2_2(mux_2948_nl, mux_2929_nl, fsm_output[3]);
  assign mux_2976_nl = MUX_s_1_2_2(mux_2975_nl, mux_2949_nl, fsm_output[2]);
  assign COMP_LOOP_mux1h_428_nl = MUX1HOT_s_1_6_2((operator_66_true_div_cmp_z[0]),
      (tmp_10_lpi_4_dfm[0]), (z_out_6[5]), COMP_LOOP_nor_12_itm, COMP_LOOP_nor_11_itm,
      COMP_LOOP_nor_11_nl, {COMP_LOOP_and_274_nl , and_dcpl_281 , and_dcpl_119 ,
      not_tmp_646 , (~ mux_2976_nl) , COMP_LOOP_or_32_cse});
  assign or_3351_nl = (fsm_output[4]) | (~ (fsm_output[2])) | (fsm_output[6]) | (fsm_output[3])
      | (fsm_output[8]) | (fsm_output[9]) | not_tmp_45;
  assign or_2678_nl = (fsm_output[9:8]!=2'b01) | not_tmp_45;
  assign mux_2885_nl = MUX_s_1_2_2(or_2679_cse, or_2678_nl, fsm_output[3]);
  assign nor_667_nl = ~((fsm_output[6]) | mux_2885_nl);
  assign nor_668_nl = ~((~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[8])
      | (fsm_output[9]) | (~ (fsm_output[5])) | (fsm_output[10]));
  assign mux_2886_nl = MUX_s_1_2_2(nor_667_nl, nor_668_nl, fsm_output[2]);
  assign nand_421_nl = ~((fsm_output[4]) & mux_2886_nl);
  assign mux_2887_nl = MUX_s_1_2_2(or_3351_nl, nand_421_nl, fsm_output[7]);
  assign or_2674_nl = (fsm_output[3]) | (fsm_output[8]) | (fsm_output[9]) | (~ (fsm_output[5]))
      | (fsm_output[10]);
  assign or_2673_nl = (~ (fsm_output[3])) | (~ (fsm_output[8])) | (~ (fsm_output[9]))
      | (fsm_output[5]) | (fsm_output[10]);
  assign mux_2883_nl = MUX_s_1_2_2(or_2674_nl, or_2673_nl, fsm_output[6]);
  assign or_3352_nl = (~ (fsm_output[4])) | (fsm_output[2]) | mux_2883_nl;
  assign nor_671_nl = ~((fsm_output[9:8]!=2'b00) | not_tmp_45);
  assign mux_2882_nl = MUX_s_1_2_2(nor_670_cse, nor_671_nl, fsm_output[3]);
  assign nand_422_nl = ~(nor_381_cse & mux_2882_nl);
  assign mux_2884_nl = MUX_s_1_2_2(or_3352_nl, nand_422_nl, fsm_output[7]);
  assign mux_2888_nl = MUX_s_1_2_2(mux_2887_nl, mux_2884_nl, fsm_output[1]);
  assign nor_646_nl = ~((~ (fsm_output[7])) | (fsm_output[1]) | (~ (fsm_output[3]))
      | (fsm_output[6]) | (fsm_output[5]) | (~ (fsm_output[10])));
  assign nor_647_nl = ~((fsm_output[7]) | (fsm_output[1]) | (fsm_output[3]) | (~
      (fsm_output[6])) | (~ (fsm_output[5])) | (fsm_output[10]));
  assign mux_2980_nl = MUX_s_1_2_2(nor_646_nl, nor_647_nl, fsm_output[8]);
  assign nor_648_nl = ~((~ (fsm_output[8])) | (fsm_output[7]) | (~ (fsm_output[1]))
      | (fsm_output[3]) | (~ (fsm_output[6])) | (fsm_output[5]) | (~ (fsm_output[10])));
  assign mux_2981_nl = MUX_s_1_2_2(mux_2980_nl, nor_648_nl, fsm_output[4]);
  assign nor_649_nl = ~((fsm_output[4]) | (fsm_output[8]) | (fsm_output[7]) | (~
      (fsm_output[1])) | (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5]))
      | (fsm_output[10]));
  assign mux_2982_nl = MUX_s_1_2_2(mux_2981_nl, nor_649_nl, fsm_output[9]);
  assign nor_650_nl = ~((~ (fsm_output[4])) | (fsm_output[8]) | (~ (fsm_output[7]))
      | (~ (fsm_output[1])) | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[5])
      | (fsm_output[10]));
  assign nor_651_nl = ~((fsm_output[1]) | (~ (fsm_output[3])) | (fsm_output[6]) |
      (fsm_output[5]) | (~ (fsm_output[10])));
  assign nor_652_nl = ~((fsm_output[1]) | (fsm_output[3]) | (~ (fsm_output[6])) |
      (~ (fsm_output[5])) | (fsm_output[10]));
  assign mux_2977_nl = MUX_s_1_2_2(nor_651_nl, nor_652_nl, fsm_output[7]);
  assign nor_653_nl = ~((~ (fsm_output[7])) | (~ (fsm_output[1])) | (~ (fsm_output[3]))
      | (fsm_output[6]) | (~ (fsm_output[5])) | (fsm_output[10]));
  assign mux_2978_nl = MUX_s_1_2_2(mux_2977_nl, nor_653_nl, fsm_output[8]);
  assign and_490_nl = (fsm_output[4]) & mux_2978_nl;
  assign mux_2979_nl = MUX_s_1_2_2(nor_650_nl, and_490_nl, fsm_output[9]);
  assign mux_2983_nl = MUX_s_1_2_2(mux_2982_nl, mux_2979_nl, fsm_output[2]);
  assign COMP_LOOP_mux1h_464_nl = MUX1HOT_s_1_4_2((COMP_LOOP_k_9_4_sva_4_0[3]), COMP_LOOP_nor_134_itm,
      modExp_exp_1_7_1_sva, (COMP_LOOP_k_9_4_sva_4_0[4]), {and_dcpl_283 , and_dcpl_332
      , (~ mux_3369_itm) , not_tmp_762});
  assign nor_580_nl = ~((fsm_output[6]) | mux_3394_cse);
  assign mux_3395_nl = MUX_s_1_2_2(nor_580_nl, mux_3392_cse, fsm_output[3]);
  assign mux_3396_nl = MUX_s_1_2_2(mux_3395_nl, mux_3388_cse, fsm_output[9]);
  assign COMP_LOOP_nor_12_nl = ~((z_out_7[4]) | (z_out_7[3]) | (z_out_7[1]));
  assign mux_3487_nl = MUX_s_1_2_2(mux_tmp_3452, mux_tmp_3450, and_573_cse);
  assign mux_3486_nl = MUX_s_1_2_2(mux_tmp_3450, mux_tmp_3449, or_2348_cse);
  assign mux_3488_nl = MUX_s_1_2_2(mux_3487_nl, mux_3486_nl, fsm_output[2]);
  assign mux_3483_nl = MUX_s_1_2_2((~ or_212_cse), and_tmp_36, fsm_output[5]);
  assign mux_3482_nl = MUX_s_1_2_2((~ or_212_cse), (fsm_output[8]), fsm_output[5]);
  assign mux_3484_nl = MUX_s_1_2_2(mux_3483_nl, mux_3482_nl, fsm_output[1]);
  assign mux_3480_nl = MUX_s_1_2_2(mux_tmp_3456, (fsm_output[8]), fsm_output[5]);
  assign mux_3481_nl = MUX_s_1_2_2(mux_3480_nl, mux_tmp_3471, fsm_output[1]);
  assign mux_3485_nl = MUX_s_1_2_2(mux_3484_nl, mux_3481_nl, fsm_output[2]);
  assign mux_3489_nl = MUX_s_1_2_2(mux_3488_nl, (~ mux_3485_nl), fsm_output[6]);
  assign mux_3478_nl = MUX_s_1_2_2(mux_tmp_3426, or_2729_cse, fsm_output[5]);
  assign mux_3476_nl = MUX_s_1_2_2((~ and_tmp_36), mux_tmp_3426, fsm_output[5]);
  assign mux_3477_nl = MUX_s_1_2_2(mux_3476_nl, mux_tmp_3452, and_565_cse);
  assign mux_3479_nl = MUX_s_1_2_2(mux_3478_nl, mux_3477_nl, fsm_output[6]);
  assign mux_3490_nl = MUX_s_1_2_2(mux_3489_nl, mux_3479_nl, fsm_output[7]);
  assign mux_3469_nl = MUX_s_1_2_2((~ mux_tmp_3468), nand_tmp_167, fsm_output[5]);
  assign mux_3470_nl = MUX_s_1_2_2(mux_3469_nl, mux_tmp_3467, fsm_output[0]);
  assign mux_3472_nl = MUX_s_1_2_2((~ mux_tmp_3471), mux_3470_nl, fsm_output[1]);
  assign mux_3473_nl = MUX_s_1_2_2(mux_3472_nl, mux_tmp_3467, fsm_output[2]);
  assign mux_3474_nl = MUX_s_1_2_2(mux_tmp_3449, mux_3473_nl, fsm_output[6]);
  assign mux_3462_nl = MUX_s_1_2_2(or_tmp_150, or_2729_cse, fsm_output[5]);
  assign mux_3461_nl = MUX_s_1_2_2((~ or_tmp_150), mux_tmp_3458, fsm_output[5]);
  assign mux_3463_nl = MUX_s_1_2_2((~ mux_3462_nl), mux_3461_nl, fsm_output[0]);
  assign mux_3464_nl = MUX_s_1_2_2(mux_3463_nl, mux_tmp_3459, fsm_output[1]);
  assign mux_3457_nl = MUX_s_1_2_2((~ or_tmp_191), mux_tmp_3456, fsm_output[5]);
  assign mux_3460_nl = MUX_s_1_2_2(mux_tmp_3459, mux_3457_nl, fsm_output[1]);
  assign mux_3465_nl = MUX_s_1_2_2(mux_3464_nl, mux_3460_nl, fsm_output[2]);
  assign mux_3453_nl = MUX_s_1_2_2(mux_tmp_3452, mux_tmp_3450, fsm_output[0]);
  assign mux_3451_nl = MUX_s_1_2_2(mux_tmp_3450, mux_tmp_3449, fsm_output[0]);
  assign mux_3454_nl = MUX_s_1_2_2(mux_3453_nl, mux_3451_nl, fsm_output[1]);
  assign mux_3455_nl = MUX_s_1_2_2(mux_tmp_3452, mux_3454_nl, fsm_output[2]);
  assign mux_3466_nl = MUX_s_1_2_2((~ mux_3465_nl), mux_3455_nl, fsm_output[6]);
  assign mux_3475_nl = MUX_s_1_2_2(mux_3474_nl, mux_3466_nl, fsm_output[7]);
  assign mux_3491_nl = MUX_s_1_2_2(mux_3490_nl, mux_3475_nl, fsm_output[3]);
  assign mux_3443_nl = MUX_s_1_2_2(or_2729_cse, or_tmp_118, fsm_output[5]);
  assign mux_3442_nl = MUX_s_1_2_2(or_212_cse, or_tmp_118, fsm_output[5]);
  assign mux_3444_nl = MUX_s_1_2_2(mux_3443_nl, mux_3442_nl, fsm_output[1]);
  assign mux_3445_nl = MUX_s_1_2_2(mux_3444_nl, mux_tmp_226, fsm_output[2]);
  assign mux_3446_nl = MUX_s_1_2_2(mux_tmp_3430, mux_3445_nl, fsm_output[6]);
  assign mux_3438_nl = MUX_s_1_2_2(or_163_cse, or_tmp_110, fsm_output[5]);
  assign mux_3439_nl = MUX_s_1_2_2(mux_3438_nl, mux_tmp_3436, or_2348_cse);
  assign mux_3437_nl = MUX_s_1_2_2(mux_tmp_3436, mux_tmp_207, and_573_cse);
  assign mux_3440_nl = MUX_s_1_2_2(mux_3439_nl, mux_3437_nl, fsm_output[2]);
  assign mux_3434_nl = MUX_s_1_2_2(or_tmp_118, or_163_cse, fsm_output[5]);
  assign mux_3435_nl = MUX_s_1_2_2(mux_3434_nl, mux_tmp_3418, and_563_cse);
  assign mux_3441_nl = MUX_s_1_2_2(mux_3440_nl, mux_3435_nl, fsm_output[6]);
  assign mux_3447_nl = MUX_s_1_2_2(mux_3446_nl, mux_3441_nl, fsm_output[7]);
  assign mux_3428_nl = MUX_s_1_2_2(or_163_cse, (fsm_output[8]), fsm_output[5]);
  assign mux_3427_nl = MUX_s_1_2_2(mux_tmp_3426, (fsm_output[8]), fsm_output[5]);
  assign mux_3429_nl = MUX_s_1_2_2(mux_3428_nl, mux_3427_nl, fsm_output[1]);
  assign mux_3431_nl = MUX_s_1_2_2(mux_tmp_3430, mux_3429_nl, fsm_output[2]);
  assign mux_3424_nl = MUX_s_1_2_2(mux_tmp_226, mux_tmp_3422, and_573_cse);
  assign mux_3425_nl = MUX_s_1_2_2(mux_3424_nl, mux_tmp_3422, fsm_output[2]);
  assign mux_3432_nl = MUX_s_1_2_2(mux_3431_nl, mux_3425_nl, fsm_output[6]);
  assign mux_3420_nl = MUX_s_1_2_2(mux_tmp_207, mux_tmp_3418, fsm_output[6]);
  assign mux_3433_nl = MUX_s_1_2_2(mux_3432_nl, mux_3420_nl, fsm_output[7]);
  assign mux_3448_nl = MUX_s_1_2_2(mux_3447_nl, mux_3433_nl, fsm_output[3]);
  assign mux_3492_nl = MUX_s_1_2_2(mux_3491_nl, mux_3448_nl, fsm_output[9]);
  assign or_3090_nl = (fsm_output[6]) | mux_3394_cse;
  assign or_3084_nl = (fsm_output[0]) | mux_tmp_3386;
  assign or_3083_nl = (~ (fsm_output[5])) | (~ (fsm_output[1])) | (fsm_output[2])
      | (fsm_output[7]) | not_tmp_34;
  assign mux_3499_nl = MUX_s_1_2_2(or_3002_cse, mux_3498_cse, fsm_output[1]);
  assign or_3079_nl = (fsm_output[1]) | (~ (fsm_output[2])) | (~ (fsm_output[7]))
      | (~ (fsm_output[8])) | (fsm_output[4]) | (fsm_output[10]);
  assign mux_3500_nl = MUX_s_1_2_2(mux_3499_nl, or_3079_nl, fsm_output[5]);
  assign mux_3501_nl = MUX_s_1_2_2(or_3083_nl, mux_3500_nl, fsm_output[0]);
  assign mux_3502_nl = MUX_s_1_2_2(or_3084_nl, mux_3501_nl, fsm_output[6]);
  assign mux_3505_nl = MUX_s_1_2_2(or_3090_nl, mux_3502_nl, fsm_output[3]);
  assign nand_168_nl = ~((fsm_output[0]) & (~ mux_tmp_3386));
  assign or_3076_nl = (fsm_output[0]) | mux_3385_cse;
  assign mux_3496_nl = MUX_s_1_2_2(nand_168_nl, or_3076_nl, fsm_output[6]);
  assign or_3071_nl = (fsm_output[6]) | (fsm_output[0]) | (fsm_output[5]) | (fsm_output[1])
      | (~ (fsm_output[2])) | (fsm_output[7]) | (~ (fsm_output[8])) | (~ (fsm_output[4]))
      | (fsm_output[10]);
  assign mux_3497_nl = MUX_s_1_2_2(mux_3496_nl, or_3071_nl, fsm_output[3]);
  assign mux_3506_nl = MUX_s_1_2_2(mux_3505_nl, mux_3497_nl, fsm_output[9]);
  assign COMP_LOOP_mux1h_474_nl = MUX1HOT_s_1_3_2(COMP_LOOP_nor_12_itm, COMP_LOOP_nor_134_itm,
      COMP_LOOP_nor_12_nl, {(~ mux_3492_nl) , (~ mux_3506_nl) , COMP_LOOP_or_32_cse});
  assign or_3055_nl = (fsm_output[6]) | (fsm_output[8]) | (~ (fsm_output[5])) | (~
      (fsm_output[0])) | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[10]);
  assign or_3054_nl = (fsm_output[8]) | (~ (fsm_output[5])) | (fsm_output[0]) | (fsm_output[3])
      | (fsm_output[9]) | (fsm_output[10]);
  assign or_3052_nl = (~ (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[10]);
  assign or_3051_nl = (fsm_output[3]) | (fsm_output[9]) | (~ (fsm_output[10]));
  assign mux_3414_nl = MUX_s_1_2_2(or_3052_nl, or_3051_nl, fsm_output[0]);
  assign or_3053_nl = (~ (fsm_output[8])) | (fsm_output[5]) | mux_3414_nl;
  assign mux_3415_nl = MUX_s_1_2_2(or_3054_nl, or_3053_nl, fsm_output[6]);
  assign mux_3416_nl = MUX_s_1_2_2(or_3055_nl, mux_3415_nl, fsm_output[4]);
  assign nor_569_nl = ~((fsm_output[7]) | mux_3416_nl);
  assign nor_570_nl = ~((~ (fsm_output[5])) | (fsm_output[0]) | (~ (fsm_output[3]))
      | (fsm_output[9]) | (~ (fsm_output[10])));
  assign nor_571_nl = ~((fsm_output[5]) | (fsm_output[0]) | (fsm_output[3]) | (fsm_output[9])
      | (fsm_output[10]));
  assign mux_3412_nl = MUX_s_1_2_2(nor_570_nl, nor_571_nl, fsm_output[8]);
  assign and_410_nl = (fsm_output[6]) & mux_3412_nl;
  assign or_3044_nl = (fsm_output[5]) | (~ (fsm_output[0])) | (fsm_output[3]) | (fsm_output[9])
      | (fsm_output[10]);
  assign nand_208_nl = ~((fsm_output[5]) & (fsm_output[0]) & (fsm_output[3]) & (fsm_output[9])
      & (~ (fsm_output[10])));
  assign mux_3411_nl = MUX_s_1_2_2(or_3044_nl, nand_208_nl, fsm_output[8]);
  assign nor_572_nl = ~((fsm_output[6]) | mux_3411_nl);
  assign mux_3413_nl = MUX_s_1_2_2(and_410_nl, nor_572_nl, fsm_output[4]);
  assign and_409_nl = (fsm_output[7]) & mux_3413_nl;
  assign mux_3417_nl = MUX_s_1_2_2(nor_569_nl, and_409_nl, fsm_output[2]);
  assign or_3348_nl = (~ (fsm_output[2])) | (fsm_output[7]) | (fsm_output[6]) | (~
      (fsm_output[5])) | (fsm_output[3]) | (fsm_output[8]) | (~ (fsm_output[10]));
  assign or_3099_nl = (~ (fsm_output[6])) | (~ (fsm_output[5])) | (fsm_output[3])
      | (~ (fsm_output[8])) | (fsm_output[10]);
  assign mux_3510_nl = MUX_s_1_2_2(or_3099_nl, or_tmp_3025, fsm_output[7]);
  assign or_3349_nl = (fsm_output[2]) | mux_3510_nl;
  assign mux_3511_nl = MUX_s_1_2_2(or_3348_nl, or_3349_nl, fsm_output[0]);
  assign or_3097_nl = (~ (fsm_output[7])) | (fsm_output[6]) | (~((fsm_output[5])
      & (fsm_output[3]) & (fsm_output[8]) & (fsm_output[10])));
  assign or_3095_nl = (~ (fsm_output[7])) | (~ (fsm_output[6])) | (~ (fsm_output[5]))
      | (~ (fsm_output[3])) | (fsm_output[8]) | (fsm_output[10]);
  assign mux_3509_nl = MUX_s_1_2_2(or_3097_nl, or_3095_nl, fsm_output[2]);
  assign or_3350_nl = (fsm_output[0]) | mux_3509_nl;
  assign mux_3512_nl = MUX_s_1_2_2(mux_3511_nl, or_3350_nl, fsm_output[4]);
  assign nor_567_nl = ~((fsm_output[2]) | (~ (fsm_output[7])) | (fsm_output[6]) |
      (fsm_output[5]) | (fsm_output[3]) | (fsm_output[8]) | (fsm_output[10]));
  assign or_3091_nl = (~ (fsm_output[6])) | (~ (fsm_output[5])) | (fsm_output[3])
      | (fsm_output[8]) | (fsm_output[10]);
  assign mux_3507_nl = MUX_s_1_2_2(or_tmp_3025, or_3091_nl, fsm_output[7]);
  assign and_402_nl = (fsm_output[2]) & (~ mux_3507_nl);
  assign mux_3508_nl = MUX_s_1_2_2(nor_567_nl, and_402_nl, fsm_output[0]);
  assign nand_420_nl = ~((fsm_output[4]) & mux_3508_nl);
  assign mux_3513_nl = MUX_s_1_2_2(mux_3512_nl, nand_420_nl, fsm_output[9]);
  assign COMP_LOOP_nor_14_nl = ~((z_out_7[4]) | (z_out_7[2]) | (z_out_7[1]));
  assign mux_3558_nl = MUX_s_1_2_2(mux_tmp_379, mux_tmp_3323, fsm_output[1]);
  assign mux_3559_nl = MUX_s_1_2_2(mux_382_cse, mux_3558_nl, fsm_output[0]);
  assign mux_3560_nl = MUX_s_1_2_2(nand_tmp_12, mux_3559_nl, fsm_output[6]);
  assign mux_3561_nl = MUX_s_1_2_2(mux_3560_nl, mux_3557_cse, fsm_output[5]);
  assign mux_3562_nl = MUX_s_1_2_2(mux_3561_nl, mux_3555_cse, fsm_output[7]);
  assign mux_3576_nl = MUX_s_1_2_2(mux_3575_cse, mux_3562_nl, fsm_output[3]);
  assign mux_3577_nl = MUX_s_1_2_2(mux_3576_nl, mux_3551_cse, fsm_output[2]);
  assign COMP_LOOP_mux1h_477_nl = MUX1HOT_s_1_4_2((COMP_LOOP_k_9_4_sva_4_0[4]), COMP_LOOP_nor_137_itm,
      COMP_LOOP_nor_134_itm, COMP_LOOP_nor_14_nl, {and_dcpl_283 , not_tmp_776 , (~
      mux_3577_nl) , COMP_LOOP_or_32_cse});
  assign nor_558_nl = ~((~ (fsm_output[5])) | (fsm_output[3]) | (fsm_output[6]) |
      (fsm_output[9]) | (fsm_output[8]) | (fsm_output[4]) | (~ (fsm_output[10])));
  assign nor_559_nl = ~((~ (fsm_output[5])) | (~ (fsm_output[3])) | (~ (fsm_output[6]))
      | (fsm_output[9]) | (fsm_output[8]) | (~ (fsm_output[4])) | (fsm_output[10]));
  assign mux_3582_nl = MUX_s_1_2_2(nor_558_nl, nor_559_nl, fsm_output[7]);
  assign nand_452_nl = ~((fsm_output[2]) & mux_3582_nl);
  assign or_3474_nl = (fsm_output[10:2]!=9'b011010110);
  assign mux_3583_nl = MUX_s_1_2_2(nand_452_nl, or_3474_nl, fsm_output[1]);
  assign or_3127_nl = (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[9])
      | (fsm_output[8]) | (~ (fsm_output[4])) | (fsm_output[10]);
  assign or_3126_nl = (fsm_output[3]) | (~ (fsm_output[6])) | (fsm_output[9]) | (~
      (fsm_output[8])) | (fsm_output[4]) | (fsm_output[10]);
  assign mux_3579_nl = MUX_s_1_2_2(or_3127_nl, or_3126_nl, fsm_output[5]);
  assign or_3125_nl = (fsm_output[5]) | (~ (fsm_output[3])) | (fsm_output[6]) | (fsm_output[9])
      | (fsm_output[8]) | (fsm_output[4]) | (~ (fsm_output[10]));
  assign mux_3580_nl = MUX_s_1_2_2(mux_3579_nl, or_3125_nl, fsm_output[7]);
  assign or_3475_nl = (fsm_output[2]) | mux_3580_nl;
  assign nor_562_nl = ~((fsm_output[3]) | (fsm_output[6]) | (fsm_output[9]) | (fsm_output[8])
      | (~ (fsm_output[4])) | (fsm_output[10]));
  assign nor_563_nl = ~((~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[9]))
      | (~ (fsm_output[8])) | (~ (fsm_output[4])) | (fsm_output[10]));
  assign mux_3578_nl = MUX_s_1_2_2(nor_562_nl, nor_563_nl, fsm_output[5]);
  assign nand_453_nl = ~((fsm_output[2]) & (fsm_output[7]) & mux_3578_nl);
  assign mux_3581_nl = MUX_s_1_2_2(or_3475_nl, nand_453_nl, fsm_output[1]);
  assign mux_3584_nl = MUX_s_1_2_2(mux_3583_nl, mux_3581_nl, fsm_output[0]);
  assign or_3145_nl = (~ (fsm_output[5])) | (fsm_output[9]) | not_tmp_51;
  assign mux_3589_nl = MUX_s_1_2_2(or_2679_cse, or_3145_nl, fsm_output[3]);
  assign nor_552_nl = ~((fsm_output[2]) | (~ (fsm_output[4])) | (fsm_output[6]) |
      mux_3589_nl);
  assign nor_554_nl = ~((~ (fsm_output[5])) | (fsm_output[9]) | (fsm_output[8]) |
      (~ (fsm_output[10])));
  assign mux_3588_nl = MUX_s_1_2_2(nor_670_cse, nor_554_nl, fsm_output[3]);
  assign and_392_nl = nor_381_cse & mux_3588_nl;
  assign mux_3590_nl = MUX_s_1_2_2(nor_552_nl, and_392_nl, fsm_output[1]);
  assign and_391_nl = (fsm_output[7]) & mux_3590_nl;
  assign nor_555_nl = ~((~ (fsm_output[2])) | (~ (fsm_output[4])) | (fsm_output[6])
      | (~ (fsm_output[3])) | (fsm_output[5]) | (~ (fsm_output[9])) | (fsm_output[8])
      | (~ (fsm_output[10])));
  assign or_3136_nl = (fsm_output[6]) | (~ (fsm_output[3])) | (~ (fsm_output[5]))
      | (~ (fsm_output[9])) | (fsm_output[8]) | (fsm_output[10]);
  assign or_3135_nl = (~ (fsm_output[6])) | (fsm_output[3]) | (fsm_output[5]) | (fsm_output[9])
      | not_tmp_51;
  assign mux_3585_nl = MUX_s_1_2_2(or_3136_nl, or_3135_nl, fsm_output[4]);
  assign nor_556_nl = ~((fsm_output[2]) | mux_3585_nl);
  assign mux_3586_nl = MUX_s_1_2_2(nor_555_nl, nor_556_nl, fsm_output[1]);
  assign nor_557_nl = ~((fsm_output[1]) | (~ (fsm_output[2])) | (~ (fsm_output[4]))
      | (~ (fsm_output[6])) | (fsm_output[3]) | (~ (fsm_output[5])) | (~ (fsm_output[9]))
      | (fsm_output[8]) | (fsm_output[10]));
  assign mux_3587_nl = MUX_s_1_2_2(mux_3586_nl, nor_557_nl, fsm_output[7]);
  assign mux_3591_nl = MUX_s_1_2_2(and_391_nl, mux_3587_nl, fsm_output[0]);
  assign COMP_LOOP_nor_17_nl = ~((z_out_7[3:1]!=3'b000));
  assign COMP_LOOP_mux1h_479_nl = MUX1HOT_s_1_3_2(COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm,
      COMP_LOOP_nor_137_itm, COMP_LOOP_nor_17_nl, {not_tmp_776 , (~ mux_3369_itm)
      , COMP_LOOP_or_32_cse});
  assign or_3158_nl = (fsm_output[6]) | (fsm_output[2]) | (~ (fsm_output[7])) | (~
      (fsm_output[4])) | (fsm_output[8]) | (~ (fsm_output[9]));
  assign or_3156_nl = (~ (fsm_output[6])) | (~ (fsm_output[2])) | (~ (fsm_output[7]))
      | (fsm_output[4]) | (~ (fsm_output[8])) | (fsm_output[9]);
  assign mux_3596_nl = MUX_s_1_2_2(or_3158_nl, or_3156_nl, fsm_output[1]);
  assign or_3155_nl = (~ (fsm_output[1])) | (fsm_output[6]) | (~ (fsm_output[2]))
      | (~ (fsm_output[7])) | (~ (fsm_output[4])) | (fsm_output[8]) | (fsm_output[9]);
  assign mux_3597_nl = MUX_s_1_2_2(mux_3596_nl, or_3155_nl, fsm_output[0]);
  assign or_3342_nl = (fsm_output[3]) | mux_3597_nl;
  assign or_3343_nl = (~ (fsm_output[1])) | (fsm_output[6]) | (fsm_output[2]) | (fsm_output[7])
      | (~ (fsm_output[4])) | (fsm_output[8]) | (fsm_output[9]);
  assign nor_548_nl = ~((fsm_output[7]) | (fsm_output[4]) | (~ (fsm_output[8])) |
      (fsm_output[9]));
  assign and_820_nl = (fsm_output[7]) & (fsm_output[4]) & (~ (fsm_output[8])) & (fsm_output[9]);
  assign mux_3593_nl = MUX_s_1_2_2(nor_548_nl, and_820_nl, fsm_output[2]);
  assign nand_419_nl = ~((~((fsm_output[1]) | (~ (fsm_output[6])))) & mux_3593_nl);
  assign mux_3594_nl = MUX_s_1_2_2(or_3343_nl, nand_419_nl, fsm_output[0]);
  assign or_3344_nl = (fsm_output[1]) | (~ (fsm_output[6])) | (~ (fsm_output[2]))
      | (~ (fsm_output[7])) | (~ (fsm_output[4])) | (fsm_output[8]) | (fsm_output[9]);
  assign or_3345_nl = (~ (fsm_output[1])) | (fsm_output[6]) | (fsm_output[2]) | (fsm_output[7])
      | (fsm_output[4]) | (fsm_output[8]) | (~ (fsm_output[9]));
  assign mux_3592_nl = MUX_s_1_2_2(or_3344_nl, or_3345_nl, fsm_output[0]);
  assign mux_3595_nl = MUX_s_1_2_2(mux_3594_nl, mux_3592_nl, fsm_output[3]);
  assign mux_3598_nl = MUX_s_1_2_2(or_3342_nl, mux_3595_nl, fsm_output[5]);
  assign nand_181_nl = ~((fsm_output[5]) & mux_3603_cse);
  assign nor_541_nl = ~((~ (fsm_output[2])) | (~ (fsm_output[9])) | (fsm_output[8])
      | nand_398_cse);
  assign nor_542_nl = ~((fsm_output[2]) | (fsm_output[9]) | (fsm_output[8]) | (fsm_output[4])
      | (~ (fsm_output[10])));
  assign mux_3602_nl = MUX_s_1_2_2(nor_541_nl, nor_542_nl, fsm_output[7]);
  assign nand_180_nl = ~(nor_515_cse & mux_3602_nl);
  assign mux_3604_nl = MUX_s_1_2_2(nand_181_nl, nand_180_nl, fsm_output[0]);
  assign nor_538_nl = ~((fsm_output[6]) | mux_3604_nl);
  assign and_389_nl = (fsm_output[0]) & (fsm_output[5]) & (fsm_output[3]) & (fsm_output[7])
      & (fsm_output[2]) & (fsm_output[9]) & (fsm_output[8]) & (fsm_output[4]) & (~
      (fsm_output[10]));
  assign nor_543_nl = ~((~ (fsm_output[3])) | (fsm_output[7]) | (fsm_output[2]) |
      (~ (fsm_output[9])) | (~ (fsm_output[8])) | (~ (fsm_output[4])) | (fsm_output[10]));
  assign mux_3599_nl = MUX_s_1_2_2(nor_543_nl, nor_544_cse, fsm_output[5]);
  assign mux_3600_nl = MUX_s_1_2_2(mux_3599_nl, nor_545_cse, fsm_output[0]);
  assign mux_3601_nl = MUX_s_1_2_2(and_389_nl, mux_3600_nl, fsm_output[6]);
  assign mux_3605_nl = MUX_s_1_2_2(nor_538_nl, mux_3601_nl, fsm_output[1]);
  assign mux_3668_nl = MUX_s_1_2_2(nand_tmp_119, or_tmp_3107, fsm_output[7]);
  assign mux_3667_nl = MUX_s_1_2_2((~ nor_tmp_286), (fsm_output[6]), fsm_output[7]);
  assign mux_3669_nl = MUX_s_1_2_2(mux_3668_nl, mux_3667_nl, fsm_output[5]);
  assign nand_195_nl = ~((fsm_output[6]) & ((fsm_output[1:0]!=2'b00) | (~ nor_tmp_6)));
  assign mux_3665_nl = MUX_s_1_2_2(nand_195_nl, or_tmp_434, fsm_output[7]);
  assign and_388_nl = ((fsm_output[6]) | (fsm_output[0]) | (fsm_output[1]) | (fsm_output[3]))
      & (fsm_output[10]);
  assign mux_3664_nl = MUX_s_1_2_2(and_388_nl, nand_tmp_119, fsm_output[7]);
  assign mux_3666_nl = MUX_s_1_2_2((~ mux_3665_nl), mux_3664_nl, fsm_output[5]);
  assign mux_3670_nl = MUX_s_1_2_2((~ mux_3669_nl), mux_3666_nl, fsm_output[2]);
  assign mux_3661_nl = MUX_s_1_2_2(not_tmp_378, mux_tmp_2696, fsm_output[7]);
  assign mux_3659_nl = MUX_s_1_2_2((~ or_tmp_2269), or_tmp_9, fsm_output[6]);
  assign and_386_nl = (fsm_output[6]) & or_tmp_2483;
  assign mux_3660_nl = MUX_s_1_2_2(mux_3659_nl, and_386_nl, fsm_output[7]);
  assign mux_3662_nl = MUX_s_1_2_2(mux_3661_nl, mux_3660_nl, fsm_output[5]);
  assign or_3182_nl = (fsm_output[6]) | (~ or_tmp_2275);
  assign and_385_nl = (fsm_output[6]) & or_tmp_2220;
  assign mux_3657_nl = MUX_s_1_2_2(or_3182_nl, and_385_nl, fsm_output[7]);
  assign mux_3658_nl = MUX_s_1_2_2(mux_tmp_2290, mux_3657_nl, fsm_output[5]);
  assign mux_3663_nl = MUX_s_1_2_2(mux_3662_nl, mux_3658_nl, fsm_output[2]);
  assign mux_3671_nl = MUX_s_1_2_2(mux_3670_nl, mux_3663_nl, fsm_output[8]);
  assign mux_3653_nl = MUX_s_1_2_2(and_tmp_16, (~ or_tmp_2479), fsm_output[7]);
  assign mux_3652_nl = MUX_s_1_2_2(or_15_cse, mux_tmp_893, fsm_output[7]);
  assign mux_3654_nl = MUX_s_1_2_2(mux_3653_nl, mux_3652_nl, fsm_output[5]);
  assign nand_196_nl = ~((fsm_output[6]) & or_tmp_237);
  assign mux_3650_nl = MUX_s_1_2_2(nand_196_nl, or_tmp_2479, fsm_output[7]);
  assign mux_3648_nl = MUX_s_1_2_2((~ or_tmp_2253), or_tmp_2248, fsm_output[6]);
  assign mux_3649_nl = MUX_s_1_2_2(or_tmp_4, mux_3648_nl, fsm_output[7]);
  assign mux_3651_nl = MUX_s_1_2_2((~ mux_3650_nl), mux_3649_nl, fsm_output[5]);
  assign mux_3655_nl = MUX_s_1_2_2(mux_3654_nl, mux_3651_nl, fsm_output[2]);
  assign mux_3644_nl = MUX_s_1_2_2((~ nor_tmp_6), or_tmp_2260, fsm_output[6]);
  assign mux_3645_nl = MUX_s_1_2_2(mux_3644_nl, (fsm_output[6]), fsm_output[7]);
  assign mux_3642_nl = MUX_s_1_2_2((fsm_output[10]), and_dcpl_240, fsm_output[6]);
  assign mux_3641_nl = MUX_s_1_2_2(nor_tmp_291, (fsm_output[10]), fsm_output[6]);
  assign mux_3643_nl = MUX_s_1_2_2((~ mux_3642_nl), mux_3641_nl, fsm_output[7]);
  assign mux_3646_nl = MUX_s_1_2_2(mux_3645_nl, mux_3643_nl, fsm_output[5]);
  assign nor_536_nl = ~((fsm_output[6]) | (~ nor_tmp_9));
  assign mux_3639_nl = MUX_s_1_2_2(nor_536_nl, nand_tmp_119, fsm_output[7]);
  assign nand_197_nl = ~(((~ (fsm_output[6])) | (fsm_output[3])) & (fsm_output[10]));
  assign mux_3638_nl = MUX_s_1_2_2(nand_197_nl, nor_tmp_286, fsm_output[7]);
  assign mux_3640_nl = MUX_s_1_2_2((~ mux_3639_nl), mux_3638_nl, fsm_output[5]);
  assign mux_3647_nl = MUX_s_1_2_2(mux_3646_nl, mux_3640_nl, fsm_output[2]);
  assign mux_3656_nl = MUX_s_1_2_2(mux_3655_nl, mux_3647_nl, fsm_output[8]);
  assign mux_3672_nl = MUX_s_1_2_2(mux_3671_nl, mux_3656_nl, fsm_output[4]);
  assign mux_3632_nl = MUX_s_1_2_2((~ (fsm_output[10])), nor_tmp_6, fsm_output[6]);
  assign mux_3633_nl = MUX_s_1_2_2(mux_3632_nl, or_tmp_4, fsm_output[7]);
  assign mux_3631_nl = MUX_s_1_2_2(or_tmp_434, (fsm_output[10]), fsm_output[7]);
  assign mux_3634_nl = MUX_s_1_2_2(mux_3633_nl, mux_3631_nl, fsm_output[5]);
  assign mux_3629_nl = MUX_s_1_2_2(mux_tmp_893, or_tmp_4, fsm_output[7]);
  assign mux_3627_nl = MUX_s_1_2_2(or_tmp_2479, (fsm_output[10]), fsm_output[7]);
  assign mux_3630_nl = MUX_s_1_2_2(mux_3629_nl, mux_3627_nl, fsm_output[5]);
  assign mux_3635_nl = MUX_s_1_2_2(mux_3634_nl, mux_3630_nl, fsm_output[2]);
  assign mux_3624_nl = MUX_s_1_2_2(or_tmp_14, mux_tmp_2788, fsm_output[7]);
  assign mux_3625_nl = MUX_s_1_2_2(mux_3624_nl, mux_3_cse, fsm_output[5]);
  assign mux_2589_nl = MUX_s_1_2_2(or_tmp_14, or_tmp_4, fsm_output[7]);
  assign or_3179_nl = (~ (fsm_output[6])) | (fsm_output[1]) | (fsm_output[3]) | (fsm_output[10]);
  assign mux_3622_nl = MUX_s_1_2_2(or_tmp_4, or_3179_nl, fsm_output[7]);
  assign mux_3623_nl = MUX_s_1_2_2(mux_2589_nl, mux_3622_nl, fsm_output[5]);
  assign mux_3626_nl = MUX_s_1_2_2(mux_3625_nl, mux_3623_nl, fsm_output[2]);
  assign mux_3636_nl = MUX_s_1_2_2(mux_3635_nl, mux_3626_nl, fsm_output[8]);
  assign mux_3617_nl = MUX_s_1_2_2((~ (fsm_output[10])), or_tmp_9, fsm_output[6]);
  assign or_3178_nl = (~((fsm_output[6]) | (fsm_output[0]) | (fsm_output[1]) | (fsm_output[3])))
      | (fsm_output[10]);
  assign mux_3618_nl = MUX_s_1_2_2(mux_3617_nl, or_3178_nl, fsm_output[7]);
  assign or_3176_nl = (~((fsm_output[6]) | (fsm_output[0]) | (fsm_output[1]) | (~
      (fsm_output[3])))) | (fsm_output[10]);
  assign mux_3616_nl = MUX_s_1_2_2((fsm_output[6]), or_3176_nl, fsm_output[7]);
  assign mux_3619_nl = MUX_s_1_2_2(mux_3618_nl, mux_3616_nl, fsm_output[5]);
  assign mux_3614_nl = MUX_s_1_2_2(or_tmp_3107, (fsm_output[10]), fsm_output[7]);
  assign mux_3611_nl = MUX_s_1_2_2(or_tmp_2269, or_tmp_2271, fsm_output[6]);
  assign mux_3612_nl = MUX_s_1_2_2((fsm_output[6]), mux_3611_nl, fsm_output[7]);
  assign mux_3615_nl = MUX_s_1_2_2(mux_3614_nl, mux_3612_nl, fsm_output[5]);
  assign mux_3620_nl = MUX_s_1_2_2(mux_3619_nl, mux_3615_nl, fsm_output[2]);
  assign mux_3608_nl = MUX_s_1_2_2(mux_9_cse, or_tmp_4, fsm_output[7]);
  assign mux_3609_nl = MUX_s_1_2_2(mux_3608_nl, or_tmp_2263, fsm_output[5]);
  assign mux_3606_nl = MUX_s_1_2_2(mux_tmp_2790, or_tmp_4, fsm_output[7]);
  assign mux_3607_nl = MUX_s_1_2_2(mux_3606_nl, or_tmp_2263, fsm_output[5]);
  assign mux_3610_nl = MUX_s_1_2_2(mux_3609_nl, mux_3607_nl, fsm_output[2]);
  assign mux_3621_nl = MUX_s_1_2_2(mux_3620_nl, mux_3610_nl, fsm_output[8]);
  assign mux_3637_nl = MUX_s_1_2_2(mux_3636_nl, mux_3621_nl, fsm_output[4]);
  assign mux_3673_nl = MUX_s_1_2_2(mux_3672_nl, (~ mux_3637_nl), fsm_output[9]);
  assign COMP_LOOP_or_28_nl = and_dcpl_147 | and_dcpl_217;
  assign COMP_LOOP_mux1h_480_nl = MUX1HOT_s_1_6_2(modExp_exp_1_4_1_sva, COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm,
      (COMP_LOOP_k_9_4_sva_4_0[0]), (z_out_8_8_7[0]), (z_out_9[6]), (z_out_9[5]),
      {not_tmp_776 , mux_3673_nl , not_tmp_762 , COMP_LOOP_or_28_nl , and_dcpl_182
      , and_dcpl_247});
  assign or_3297_nl = (fsm_output[7]) | (fsm_output[9]) | (fsm_output[10]);
  assign nand_250_nl = ~((fsm_output[0]) & (fsm_output[7]) & (fsm_output[9]) & (fsm_output[10]));
  assign mux_2493_nl = MUX_s_1_2_2(or_3297_nl, nand_250_nl, fsm_output[1]);
  assign mux_2494_nl = MUX_s_1_2_2(mux_2493_nl, nand_375_cse, or_495_cse);
  assign mux_2495_nl = MUX_s_1_2_2(mux_2494_nl, nand_376_cse, fsm_output[8]);
  assign nor_1453_nl = ~((~((fsm_output[2:0]!=3'b001))) | (fsm_output[4]));
  assign mux_3890_nl = MUX_s_1_2_2(nor_1453_nl, mux_tmp_3878, fsm_output[9]);
  assign mux_3891_nl = MUX_s_1_2_2(mux_3890_nl, mux_tmp_3834, fsm_output[3]);
  assign mux_3889_nl = MUX_s_1_2_2(not_tmp_1021, mux_tmp_3828, fsm_output[3]);
  assign mux_3892_nl = MUX_s_1_2_2((~ mux_3891_nl), mux_3889_nl, fsm_output[10]);
  assign and_1258_nl = ((fsm_output[9]) | (fsm_output[1]) | (~ (fsm_output[0])) |
      (fsm_output[2])) & (fsm_output[4]);
  assign mux_3886_nl = MUX_s_1_2_2((fsm_output[4]), or_tmp_3303, fsm_output[9]);
  assign mux_3887_nl = MUX_s_1_2_2(and_1258_nl, mux_3886_nl, fsm_output[3]);
  assign or_3508_nl = (fsm_output[3]) | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[4]);
  assign mux_3888_nl = MUX_s_1_2_2(mux_3887_nl, or_3508_nl, fsm_output[10]);
  assign mux_3893_nl = MUX_s_1_2_2(mux_3892_nl, mux_3888_nl, fsm_output[5]);
  assign and_1259_nl = (fsm_output[3]) & (fsm_output[9]) & (fsm_output[1]) & (fsm_output[0])
      & (fsm_output[2]) & (fsm_output[4]);
  assign mux_3883_nl = MUX_s_1_2_2((fsm_output[9]), or_2747_cse, fsm_output[3]);
  assign mux_3884_nl = MUX_s_1_2_2(and_1259_nl, mux_3883_nl, fsm_output[10]);
  assign and_1260_nl = ((fsm_output[9]) | (fsm_output[1]) | (fsm_output[0]) | (fsm_output[2]))
      & (fsm_output[4]);
  assign mux_3881_nl = MUX_s_1_2_2(mux_tmp_3853, and_1260_nl, fsm_output[3]);
  assign or_3506_nl = (fsm_output[9]) | mux_tmp_3878;
  assign mux_3880_nl = MUX_s_1_2_2(or_tmp, or_3506_nl, fsm_output[3]);
  assign mux_3882_nl = MUX_s_1_2_2((~ mux_3881_nl), mux_3880_nl, fsm_output[10]);
  assign mux_3885_nl = MUX_s_1_2_2(mux_3884_nl, mux_3882_nl, fsm_output[5]);
  assign mux_3894_nl = MUX_s_1_2_2((~ mux_3893_nl), mux_3885_nl, fsm_output[8]);
  assign or_3505_nl = (fsm_output[3]) | (fsm_output[9]);
  assign mux_3875_nl = MUX_s_1_2_2(mux_tmp_3861, (fsm_output[4]), or_3505_nl);
  assign or_3504_nl = (fsm_output[9]) | (~((fsm_output[1]) | (fsm_output[0]) | (fsm_output[2])
      | (fsm_output[4])));
  assign mux_3874_nl = MUX_s_1_2_2(or_tmp, or_3504_nl, fsm_output[3]);
  assign mux_3876_nl = MUX_s_1_2_2((~ mux_3875_nl), mux_3874_nl, fsm_output[10]);
  assign and_1256_nl = (fsm_output[3]) & (fsm_output[9]) & nor_tmp_540;
  assign or_3502_nl = (fsm_output[9]) | nor_tmp_539;
  assign mux_3872_nl = MUX_s_1_2_2(or_3502_nl, or_2747_cse, fsm_output[3]);
  assign mux_3873_nl = MUX_s_1_2_2(and_1256_nl, mux_3872_nl, fsm_output[10]);
  assign mux_3877_nl = MUX_s_1_2_2(mux_3876_nl, mux_3873_nl, fsm_output[5]);
  assign mux_3867_nl = MUX_s_1_2_2(not_tmp_1007, mux_tmp_3818, and_573_cse);
  assign mux_3868_nl = MUX_s_1_2_2((~ (fsm_output[4])), mux_3867_nl, fsm_output[9]);
  assign mux_3865_nl = MUX_s_1_2_2(not_tmp_1007, mux_tmp_3846, fsm_output[1]);
  assign mux_3866_nl = MUX_s_1_2_2(mux_3865_nl, (fsm_output[4]), fsm_output[9]);
  assign mux_3869_nl = MUX_s_1_2_2(mux_3868_nl, mux_3866_nl, fsm_output[3]);
  assign mux_3870_nl = MUX_s_1_2_2((~ mux_3869_nl), or_tmp, fsm_output[10]);
  assign mux_3863_nl = MUX_s_1_2_2((fsm_output[4]), (~ mux_tmp_3861), and_1262_cse);
  assign or_3500_nl = (fsm_output[9]) | (fsm_output[1]) | (fsm_output[2]) | (fsm_output[4]);
  assign mux_3861_nl = MUX_s_1_2_2(or_3500_nl, or_tmp, fsm_output[3]);
  assign mux_3864_nl = MUX_s_1_2_2(mux_3863_nl, mux_3861_nl, fsm_output[10]);
  assign mux_3871_nl = MUX_s_1_2_2(mux_3870_nl, mux_3864_nl, fsm_output[5]);
  assign mux_3878_nl = MUX_s_1_2_2(mux_3877_nl, mux_3871_nl, fsm_output[8]);
  assign mux_3895_nl = MUX_s_1_2_2(mux_3894_nl, mux_3878_nl, fsm_output[7]);
  assign and_1255_nl = (fsm_output[9]) & nor_tmp_536;
  assign mux_3856_nl = MUX_s_1_2_2(and_1255_nl, nor_tmp_535, fsm_output[3]);
  assign mux_3855_nl = MUX_s_1_2_2(not_tmp_1021, mux_tmp_3853, fsm_output[3]);
  assign mux_3857_nl = MUX_s_1_2_2(mux_3856_nl, (~ mux_3855_nl), fsm_output[10]);
  assign nor_1456_nl = ~(and_565_cse | (fsm_output[4]));
  assign mux_3851_nl = MUX_s_1_2_2(nor_1456_nl, nor_tmp_540, fsm_output[9]);
  assign mux_3852_nl = MUX_s_1_2_2((~ (fsm_output[4])), mux_3851_nl, fsm_output[3]);
  assign and_1264_nl = ((fsm_output[0]) | (fsm_output[2])) & (fsm_output[4]);
  assign mux_3848_nl = MUX_s_1_2_2(mux_tmp_3846, and_1264_nl, fsm_output[1]);
  assign mux_3849_nl = MUX_s_1_2_2(mux_3848_nl, (fsm_output[4]), fsm_output[9]);
  assign mux_3850_nl = MUX_s_1_2_2(mux_3849_nl, or_tmp_3304, fsm_output[3]);
  assign mux_3853_nl = MUX_s_1_2_2(mux_3852_nl, mux_3850_nl, fsm_output[10]);
  assign mux_3858_nl = MUX_s_1_2_2(mux_3857_nl, mux_3853_nl, fsm_output[5]);
  assign mux_3843_nl = MUX_s_1_2_2(or_tmp_3303, (~ nor_tmp_540), fsm_output[9]);
  assign mux_3844_nl = MUX_s_1_2_2(or_tmp_3304, mux_3843_nl, fsm_output[3]);
  assign or_3493_nl = (fsm_output[9]) | (~ nor_tmp_539);
  assign mux_3842_nl = MUX_s_1_2_2(or_3493_nl, or_tmp, fsm_output[3]);
  assign mux_3845_nl = MUX_s_1_2_2(mux_3844_nl, mux_3842_nl, fsm_output[10]);
  assign nor_1457_nl = ~((fsm_output[3]) | (fsm_output[9]) | (fsm_output[1]) | (fsm_output[0])
      | (fsm_output[2]) | (fsm_output[4]));
  assign or_3490_nl = (fsm_output[9]) | nor_tmp_536;
  assign mux_3840_nl = MUX_s_1_2_2((fsm_output[9]), or_3490_nl, fsm_output[3]);
  assign mux_3841_nl = MUX_s_1_2_2(nor_1457_nl, mux_3840_nl, fsm_output[10]);
  assign mux_3846_nl = MUX_s_1_2_2(mux_3845_nl, mux_3841_nl, fsm_output[5]);
  assign mux_3859_nl = MUX_s_1_2_2(mux_3858_nl, mux_3846_nl, fsm_output[8]);
  assign nor_1458_nl = ~(((fsm_output[0]) & (fsm_output[2])) | (fsm_output[4]));
  assign mux_3833_nl = MUX_s_1_2_2(nor_1458_nl, mux_tmp_3819, fsm_output[1]);
  assign mux_3834_nl = MUX_s_1_2_2((~ (fsm_output[4])), mux_3833_nl, fsm_output[9]);
  assign mux_3836_nl = MUX_s_1_2_2((~ mux_tmp_3834), mux_3834_nl, fsm_output[3]);
  assign mux_3832_nl = MUX_s_1_2_2(or_tmp_3293, or_2747_cse, fsm_output[3]);
  assign mux_3837_nl = MUX_s_1_2_2(mux_3836_nl, mux_3832_nl, fsm_output[10]);
  assign mux_3830_nl = MUX_s_1_2_2(mux_tmp_3828, nor_tmp_535, fsm_output[3]);
  assign mux_3828_nl = MUX_s_1_2_2(or_tmp, or_tmp_3293, fsm_output[3]);
  assign mux_3831_nl = MUX_s_1_2_2((~ mux_3830_nl), mux_3828_nl, fsm_output[10]);
  assign mux_3838_nl = MUX_s_1_2_2(mux_3837_nl, mux_3831_nl, fsm_output[5]);
  assign nor_1459_nl = ~((fsm_output[3]) | (fsm_output[9]) | or_tmp_3291);
  assign mux_3826_nl = MUX_s_1_2_2(nor_1459_nl, (fsm_output[9]), fsm_output[10]);
  assign mux_3824_nl = MUX_s_1_2_2((fsm_output[4]), (~ mux_tmp_3822), and_1262_cse);
  assign mux_3821_nl = MUX_s_1_2_2(mux_tmp_3819, nor_tmp, fsm_output[1]);
  assign or_3480_nl = (fsm_output[9]) | (~ mux_3821_nl);
  assign mux_3822_nl = MUX_s_1_2_2(or_3480_nl, or_tmp, fsm_output[3]);
  assign mux_3825_nl = MUX_s_1_2_2(mux_3824_nl, mux_3822_nl, fsm_output[10]);
  assign mux_3827_nl = MUX_s_1_2_2(mux_3826_nl, mux_3825_nl, fsm_output[5]);
  assign mux_3839_nl = MUX_s_1_2_2(mux_3838_nl, mux_3827_nl, fsm_output[8]);
  assign mux_3860_nl = MUX_s_1_2_2(mux_3859_nl, mux_3839_nl, fsm_output[7]);
  assign mux_3896_nl = MUX_s_1_2_2(mux_3895_nl, mux_3860_nl, fsm_output[6]);
  assign or_3579_nl = (~ (fsm_output[6])) | (~ (fsm_output[1])) | (~ COMP_LOOP_nor_11_itm)
      | (fsm_output[8]) | (fsm_output[10]) | not_tmp_1034;
  assign mux_3943_nl = MUX_s_1_2_2(nand_201_cse, or_tmp_3327, fsm_output[8]);
  assign nand_463_nl = ~((fsm_output[1]) & (~ mux_3943_nl));
  assign mux_3944_nl = MUX_s_1_2_2(or_tmp_3343, nand_463_nl, fsm_output[6]);
  assign mux_3945_nl = MUX_s_1_2_2(or_3579_nl, mux_3944_nl, fsm_output[3]);
  assign mux_3941_nl = MUX_s_1_2_2(or_tmp_3369, mux_tmp_3902, fsm_output[1]);
  assign or_3577_nl = (fsm_output[6]) | mux_3941_nl;
  assign mux_3942_nl = MUX_s_1_2_2(or_3577_nl, nand_tmp, fsm_output[3]);
  assign mux_3946_nl = MUX_s_1_2_2(mux_3945_nl, mux_3942_nl, fsm_output[5]);
  assign nor_1448_nl = ~((~ COMP_LOOP_nor_11_itm) | (fsm_output[8]) | (~ (fsm_output[10]))
      | (~ (fsm_output[9])) | (fsm_output[4]));
  assign nor_1449_nl = ~((~ COMP_LOOP_nor_11_itm) | (fsm_output[8]) | (fsm_output[10])
      | (fsm_output[9]) | (fsm_output[4]));
  assign mux_3938_nl = MUX_s_1_2_2(nor_1448_nl, nor_1449_nl, fsm_output[1]);
  assign nand_462_nl = ~((fsm_output[6]) & mux_3938_nl);
  assign or_3574_nl = (fsm_output[1]) | (~ COMP_LOOP_nor_11_itm) | (~ (fsm_output[8]))
      | (fsm_output[10]) | not_tmp_1034;
  assign mux_3939_nl = MUX_s_1_2_2(nand_462_nl, or_3574_nl, fsm_output[3]);
  assign or_3572_nl = (fsm_output[3]) | (fsm_output[6]) | nor_1450_cse | (fsm_output[8])
      | (~ (fsm_output[10])) | (fsm_output[9]) | (fsm_output[4]);
  assign mux_3940_nl = MUX_s_1_2_2(mux_3939_nl, or_3572_nl, fsm_output[5]);
  assign mux_3947_nl = MUX_s_1_2_2(mux_3946_nl, mux_3940_nl, fsm_output[2]);
  assign or_3568_nl = (fsm_output[6]) | mux_tmp_3898;
  assign mux_3935_nl = MUX_s_1_2_2(or_3568_nl, or_tmp_3320, fsm_output[3]);
  assign or_3567_nl = (fsm_output[1]) | (~ COMP_LOOP_nor_11_itm) | (fsm_output[8])
      | (~ (fsm_output[10])) | (fsm_output[9]) | (~ (fsm_output[4]));
  assign or_3565_nl = (fsm_output[6]) | nor_1450_cse | (~ (fsm_output[8])) | (~ (fsm_output[10]))
      | (fsm_output[9]) | (~ (fsm_output[4]));
  assign mux_3934_nl = MUX_s_1_2_2(or_3567_nl, or_3565_nl, fsm_output[3]);
  assign mux_3936_nl = MUX_s_1_2_2(mux_3935_nl, mux_3934_nl, fsm_output[5]);
  assign mux_3931_nl = MUX_s_1_2_2(or_tmp_3369, mux_tmp_3915, fsm_output[1]);
  assign nand_461_nl = ~((fsm_output[6]) & (~ mux_3931_nl));
  assign or_3559_nl = (fsm_output[6]) | (~ (fsm_output[1])) | (~ (fsm_output[8]))
      | (fsm_output[10]) | (fsm_output[9]) | (~ (fsm_output[4]));
  assign mux_3932_nl = MUX_s_1_2_2(nand_461_nl, or_3559_nl, fsm_output[3]);
  assign nand_465_nl = ~((fsm_output[6]) & (fsm_output[1]) & COMP_LOOP_nor_11_itm
      & (fsm_output[8]) & (~ (fsm_output[10])) & (fsm_output[9]) & (~ (fsm_output[4])));
  assign or_3556_nl = (~ (fsm_output[1])) | (~ COMP_LOOP_nor_11_itm) | (fsm_output[8])
      | (fsm_output[10]) | (fsm_output[9]) | (~ (fsm_output[4]));
  assign mux_3928_nl = MUX_s_1_2_2(mux_tmp_3902, mux_tmp_3906, fsm_output[1]);
  assign mux_3929_nl = MUX_s_1_2_2(or_3556_nl, mux_3928_nl, fsm_output[6]);
  assign mux_3930_nl = MUX_s_1_2_2(nand_465_nl, mux_3929_nl, fsm_output[3]);
  assign mux_3933_nl = MUX_s_1_2_2(mux_3932_nl, mux_3930_nl, fsm_output[5]);
  assign mux_3937_nl = MUX_s_1_2_2(mux_3936_nl, mux_3933_nl, fsm_output[2]);
  assign mux_3948_nl = MUX_s_1_2_2(mux_3947_nl, mux_3937_nl, fsm_output[7]);
  assign or_3554_nl = (fsm_output[8]) | (fsm_output[10]) | (fsm_output[9]) | (fsm_output[4]);
  assign mux_3922_nl = MUX_s_1_2_2(or_3554_nl, or_tmp_3332, fsm_output[1]);
  assign nand_471_nl = ~((fsm_output[1]) & (fsm_output[8]) & (fsm_output[10]) & (~
      (fsm_output[9])) & (fsm_output[4]));
  assign mux_3923_nl = MUX_s_1_2_2(mux_3922_nl, nand_471_nl, fsm_output[6]);
  assign or_3551_nl = (fsm_output[1]) | (fsm_output[8]) | (fsm_output[10]) | (fsm_output[9])
      | (fsm_output[4]);
  assign or_3550_nl = (~ (fsm_output[1])) | (~ COMP_LOOP_nor_11_itm) | (fsm_output[8])
      | (~ (fsm_output[10])) | (fsm_output[9]) | (fsm_output[4]);
  assign mux_3921_nl = MUX_s_1_2_2(or_3551_nl, or_3550_nl, fsm_output[6]);
  assign mux_3924_nl = MUX_s_1_2_2(mux_3923_nl, mux_3921_nl, fsm_output[3]);
  assign mux_3918_nl = MUX_s_1_2_2(or_tmp_195, or_tmp_182, fsm_output[8]);
  assign nand_460_nl = ~((fsm_output[1]) & COMP_LOOP_nor_11_itm & (~ mux_3918_nl));
  assign or_3548_nl = (~ COMP_LOOP_nor_11_itm) | (~ (fsm_output[8])) | (fsm_output[10])
      | (fsm_output[9]) | (fsm_output[4]);
  assign mux_3917_nl = MUX_s_1_2_2(mux_tmp_3915, or_3548_nl, fsm_output[1]);
  assign mux_3919_nl = MUX_s_1_2_2(nand_460_nl, mux_3917_nl, fsm_output[6]);
  assign or_3546_nl = (~ (fsm_output[8])) | (fsm_output[10]) | (fsm_output[9]) |
      (~ (fsm_output[4]));
  assign or_3544_nl = (fsm_output[10]) | (~ (fsm_output[9])) | (fsm_output[4]);
  assign mux_3914_nl = MUX_s_1_2_2(or_3544_nl, or_2415_cse, fsm_output[8]);
  assign mux_3915_nl = MUX_s_1_2_2(or_3546_nl, mux_3914_nl, fsm_output[1]);
  assign or_3547_nl = (fsm_output[6]) | mux_3915_nl;
  assign mux_3920_nl = MUX_s_1_2_2(mux_3919_nl, or_3547_nl, fsm_output[3]);
  assign mux_3925_nl = MUX_s_1_2_2(mux_3924_nl, mux_3920_nl, fsm_output[5]);
  assign or_3542_nl = (fsm_output[1]) | (~ COMP_LOOP_nor_11_itm) | (~ (fsm_output[8]))
      | (~ (fsm_output[10])) | (fsm_output[9]) | (~ (fsm_output[4]));
  assign or_3540_nl = (fsm_output[6]) | nor_1450_cse | (fsm_output[8]) | nand_201_cse;
  assign mux_3912_nl = MUX_s_1_2_2(or_3542_nl, or_3540_nl, fsm_output[3]);
  assign or_3536_nl = (fsm_output[1]) | (~ COMP_LOOP_nor_11_itm) | (fsm_output[8])
      | (fsm_output[10]) | (~ (fsm_output[9])) | (fsm_output[4]);
  assign mux_3911_nl = MUX_s_1_2_2(or_3536_nl, or_tmp_3343, fsm_output[6]);
  assign nand_459_nl = ~((fsm_output[3]) & (~ mux_3911_nl));
  assign mux_3913_nl = MUX_s_1_2_2(mux_3912_nl, nand_459_nl, fsm_output[5]);
  assign mux_3926_nl = MUX_s_1_2_2(mux_3925_nl, mux_3913_nl, fsm_output[2]);
  assign or_3533_nl = (fsm_output[1]) | (~ COMP_LOOP_nor_11_itm) | (~ (fsm_output[8]))
      | (fsm_output[10]) | (~ (fsm_output[9])) | (fsm_output[4]);
  assign or_3527_nl = (~ COMP_LOOP_nor_11_itm) | (fsm_output[8]) | (~ (fsm_output[10]))
      | (fsm_output[9]) | (fsm_output[4]);
  assign mux_3908_nl = MUX_s_1_2_2(mux_tmp_3906, or_3527_nl, fsm_output[1]);
  assign or_3532_nl = (fsm_output[6]) | mux_3908_nl;
  assign mux_3909_nl = MUX_s_1_2_2(or_3533_nl, or_3532_nl, fsm_output[3]);
  assign or_3534_nl = (fsm_output[5]) | mux_3909_nl;
  assign or_3589_nl = (fsm_output[6]) | (~ (fsm_output[1])) | mux_tmp_3902;
  assign mux_3904_nl = MUX_s_1_2_2(or_3589_nl, nand_tmp, fsm_output[3]);
  assign or_3521_nl = (~ (fsm_output[1])) | (~ COMP_LOOP_nor_11_itm) | (fsm_output[8])
      | (fsm_output[10]) | not_tmp_1034;
  assign mux_3900_nl = MUX_s_1_2_2(or_3521_nl, mux_tmp_3898, fsm_output[6]);
  assign or_3514_nl = (~ (fsm_output[1])) | (~ (fsm_output[8])) | (fsm_output[10])
      | not_tmp_1034;
  assign mux_3897_nl = MUX_s_1_2_2(or_3514_nl, or_tmp_3320, fsm_output[6]);
  assign mux_3901_nl = MUX_s_1_2_2(mux_3900_nl, mux_3897_nl, fsm_output[3]);
  assign mux_3905_nl = MUX_s_1_2_2(mux_3904_nl, mux_3901_nl, fsm_output[5]);
  assign mux_3910_nl = MUX_s_1_2_2(or_3534_nl, mux_3905_nl, fsm_output[2]);
  assign mux_3927_nl = MUX_s_1_2_2(mux_3926_nl, mux_3910_nl, fsm_output[7]);
  assign mux_3949_nl = MUX_s_1_2_2(mux_3948_nl, mux_3927_nl, fsm_output[0]);
  assign or_2515_nl = (fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[0])) | (fsm_output[1])
      | (~ (fsm_output[3])) | (fsm_output[10]);
  assign or_2514_nl = (~ (fsm_output[5])) | (fsm_output[7]) | (fsm_output[0]) | (fsm_output[1])
      | (fsm_output[3]) | (fsm_output[10]);
  assign mux_2648_nl = MUX_s_1_2_2(or_2515_nl, or_2514_nl, fsm_output[4]);
  assign or_2513_nl = (fsm_output[4]) | (fsm_output[5]) | (~ (fsm_output[7])) | (fsm_output[0])
      | (~ (fsm_output[1])) | (fsm_output[3]) | (~ (fsm_output[10]));
  assign mux_2649_nl = MUX_s_1_2_2(mux_2648_nl, or_2513_nl, fsm_output[9]);
  assign or_3477_nl = mux_2649_nl | (fsm_output[6]) | (fsm_output[2]) | (fsm_output[8]);
  assign or_3584_nl = (fsm_output[5:3]!=3'b110);
  assign or_3583_nl = (fsm_output[5:3]!=3'b001);
  assign mux_3950_nl = MUX_s_1_2_2(or_3584_nl, or_3583_nl, fsm_output[0]);
  assign or_3585_nl = (fsm_output[1]) | (fsm_output[9]) | (fsm_output[10]) | mux_3950_nl;
  assign or_3581_nl = (~ (fsm_output[1])) | (~ (fsm_output[9])) | (~ (fsm_output[10]))
      | (fsm_output[0]) | (fsm_output[3]) | (fsm_output[4]) | (fsm_output[5]);
  assign mux_3951_nl = MUX_s_1_2_2(or_3585_nl, or_3581_nl, fsm_output[7]);
  assign or_3587_nl = (fsm_output[6]) | mux_3951_nl;
  assign or_3588_nl = (~ (fsm_output[6])) | (fsm_output[7]) | (fsm_output[1]) | (~
      (fsm_output[9])) | (~ (fsm_output[10])) | (~ (fsm_output[0])) | (fsm_output[3])
      | (fsm_output[4]) | (fsm_output[5]);
  assign mux_3952_nl = MUX_s_1_2_2(or_3587_nl, or_3588_nl, fsm_output[2]);
  assign nor_725_nl = ~((fsm_output[7]) | (fsm_output[9]) | (fsm_output[10]));
  assign mux_2670_nl = MUX_s_1_2_2(nor_725_nl, mux_tmp_2650, and_573_cse);
  assign mux_2669_nl = MUX_s_1_2_2(mux_tmp_2650, and_815_cse, fsm_output[1]);
  assign mux_2671_nl = MUX_s_1_2_2(mux_2670_nl, mux_2669_nl, fsm_output[3]);
  assign mux_2668_nl = MUX_s_1_2_2(mux_tmp_2650, and_815_cse, fsm_output[3]);
  assign mux_2672_nl = MUX_s_1_2_2(mux_2671_nl, mux_2668_nl, fsm_output[2]);
  assign nand_244_nl = ~((fsm_output[3:0]==4'b1101));
  assign mux_2667_nl = MUX_s_1_2_2(mux_tmp_2650, and_815_cse, nand_244_nl);
  assign mux_2673_nl = MUX_s_1_2_2(mux_2672_nl, mux_2667_nl, fsm_output[4]);
  assign or_4_nl = (fsm_output[6:5]!=2'b00);
  assign mux_2674_nl = MUX_s_1_2_2(mux_2673_nl, and_815_cse, or_4_nl);
  assign mux_2675_nl = MUX_s_1_2_2(mux_2674_nl, and_816_cse, fsm_output[8]);
  assign COMP_LOOP_or_8_nl = (COMP_LOOP_COMP_LOOP_nor_itm & and_dcpl_283) | (COMP_LOOP_COMP_LOOP_and_14_itm
      & and_305_m1c) | (COMP_LOOP_COMP_LOOP_and_13_itm & and_307_m1c) | (COMP_LOOP_COMP_LOOP_and_12_itm
      & and_309_m1c) | (COMP_LOOP_COMP_LOOP_and_11_itm & and_312_m1c) | (COMP_LOOP_COMP_LOOP_and_10_itm
      & and_315_m1c) | (COMP_LOOP_COMP_LOOP_and_9_itm & and_317_m1c) | (COMP_LOOP_COMP_LOOP_and_8_itm
      & and_320_m1c) | (COMP_LOOP_COMP_LOOP_and_68_itm & and_322_m1c) | (COMP_LOOP_COMP_LOOP_and_6_itm
      & and_324_m1c) | (COMP_LOOP_COMP_LOOP_and_5_itm & and_327_m1c) | (COMP_LOOP_COMP_LOOP_and_4_itm
      & and_329_m1c) | (COMP_LOOP_COMP_LOOP_and_64_itm & and_331_m1c) | (COMP_LOOP_COMP_LOOP_and_2_itm
      & and_334_m1c) | (COMP_LOOP_COMP_LOOP_and_62_itm & and_336_m1c) | (COMP_LOOP_COMP_LOOP_and_305_itm
      & and_339_m1c);
  assign COMP_LOOP_or_9_nl = (COMP_LOOP_COMP_LOOP_and_305_itm & and_dcpl_283) | (COMP_LOOP_COMP_LOOP_nor_itm
      & and_305_m1c) | (COMP_LOOP_COMP_LOOP_and_14_itm & and_307_m1c) | (COMP_LOOP_COMP_LOOP_and_13_itm
      & and_309_m1c) | (COMP_LOOP_COMP_LOOP_and_12_itm & and_312_m1c) | (COMP_LOOP_COMP_LOOP_and_11_itm
      & and_315_m1c) | (COMP_LOOP_COMP_LOOP_and_10_itm & and_317_m1c) | (COMP_LOOP_COMP_LOOP_and_9_itm
      & and_320_m1c) | (COMP_LOOP_COMP_LOOP_and_8_itm & and_322_m1c) | (COMP_LOOP_COMP_LOOP_and_68_itm
      & and_324_m1c) | (COMP_LOOP_COMP_LOOP_and_6_itm & and_327_m1c) | (COMP_LOOP_COMP_LOOP_and_5_itm
      & and_329_m1c) | (COMP_LOOP_COMP_LOOP_and_4_itm & and_331_m1c) | (COMP_LOOP_COMP_LOOP_and_64_itm
      & and_334_m1c) | (COMP_LOOP_COMP_LOOP_and_2_itm & and_336_m1c) | (COMP_LOOP_COMP_LOOP_and_62_itm
      & and_339_m1c);
  assign COMP_LOOP_or_10_nl = (COMP_LOOP_COMP_LOOP_and_62_itm & and_dcpl_283) | (COMP_LOOP_COMP_LOOP_and_305_itm
      & and_305_m1c) | (COMP_LOOP_COMP_LOOP_nor_itm & and_307_m1c) | (COMP_LOOP_COMP_LOOP_and_14_itm
      & and_309_m1c) | (COMP_LOOP_COMP_LOOP_and_13_itm & and_312_m1c) | (COMP_LOOP_COMP_LOOP_and_12_itm
      & and_315_m1c) | (COMP_LOOP_COMP_LOOP_and_11_itm & and_317_m1c) | (COMP_LOOP_COMP_LOOP_and_10_itm
      & and_320_m1c) | (COMP_LOOP_COMP_LOOP_and_9_itm & and_322_m1c) | (COMP_LOOP_COMP_LOOP_and_8_itm
      & and_324_m1c) | (COMP_LOOP_COMP_LOOP_and_68_itm & and_327_m1c) | (COMP_LOOP_COMP_LOOP_and_6_itm
      & and_329_m1c) | (COMP_LOOP_COMP_LOOP_and_5_itm & and_331_m1c) | (COMP_LOOP_COMP_LOOP_and_4_itm
      & and_334_m1c) | (COMP_LOOP_COMP_LOOP_and_64_itm & and_336_m1c) | (COMP_LOOP_COMP_LOOP_and_2_itm
      & and_339_m1c);
  assign COMP_LOOP_or_11_nl = (COMP_LOOP_COMP_LOOP_and_2_itm & and_dcpl_283) | (COMP_LOOP_COMP_LOOP_and_62_itm
      & and_305_m1c) | (COMP_LOOP_COMP_LOOP_and_305_itm & and_307_m1c) | (COMP_LOOP_COMP_LOOP_nor_itm
      & and_309_m1c) | (COMP_LOOP_COMP_LOOP_and_14_itm & and_312_m1c) | (COMP_LOOP_COMP_LOOP_and_13_itm
      & and_315_m1c) | (COMP_LOOP_COMP_LOOP_and_12_itm & and_317_m1c) | (COMP_LOOP_COMP_LOOP_and_11_itm
      & and_320_m1c) | (COMP_LOOP_COMP_LOOP_and_10_itm & and_322_m1c) | (COMP_LOOP_COMP_LOOP_and_9_itm
      & and_324_m1c) | (COMP_LOOP_COMP_LOOP_and_8_itm & and_327_m1c) | (COMP_LOOP_COMP_LOOP_and_68_itm
      & and_329_m1c) | (COMP_LOOP_COMP_LOOP_and_6_itm & and_331_m1c) | (COMP_LOOP_COMP_LOOP_and_5_itm
      & and_334_m1c) | (COMP_LOOP_COMP_LOOP_and_4_itm & and_336_m1c) | (COMP_LOOP_COMP_LOOP_and_64_itm
      & and_339_m1c);
  assign COMP_LOOP_or_12_nl = (COMP_LOOP_COMP_LOOP_and_64_itm & and_dcpl_283) | (COMP_LOOP_COMP_LOOP_and_2_itm
      & and_305_m1c) | (COMP_LOOP_COMP_LOOP_and_62_itm & and_307_m1c) | (COMP_LOOP_COMP_LOOP_and_305_itm
      & and_309_m1c) | (COMP_LOOP_COMP_LOOP_nor_itm & and_312_m1c) | (COMP_LOOP_COMP_LOOP_and_14_itm
      & and_315_m1c) | (COMP_LOOP_COMP_LOOP_and_13_itm & and_317_m1c) | (COMP_LOOP_COMP_LOOP_and_12_itm
      & and_320_m1c) | (COMP_LOOP_COMP_LOOP_and_11_itm & and_322_m1c) | (COMP_LOOP_COMP_LOOP_and_10_itm
      & and_324_m1c) | (COMP_LOOP_COMP_LOOP_and_9_itm & and_327_m1c) | (COMP_LOOP_COMP_LOOP_and_8_itm
      & and_329_m1c) | (COMP_LOOP_COMP_LOOP_and_68_itm & and_331_m1c) | (COMP_LOOP_COMP_LOOP_and_6_itm
      & and_334_m1c) | (COMP_LOOP_COMP_LOOP_and_5_itm & and_336_m1c) | (COMP_LOOP_COMP_LOOP_and_4_itm
      & and_339_m1c);
  assign COMP_LOOP_or_13_nl = (COMP_LOOP_COMP_LOOP_and_4_itm & and_dcpl_283) | (COMP_LOOP_COMP_LOOP_and_64_itm
      & and_305_m1c) | (COMP_LOOP_COMP_LOOP_and_2_itm & and_307_m1c) | (COMP_LOOP_COMP_LOOP_and_62_itm
      & and_309_m1c) | (COMP_LOOP_COMP_LOOP_and_305_itm & and_312_m1c) | (COMP_LOOP_COMP_LOOP_nor_itm
      & and_315_m1c) | (COMP_LOOP_COMP_LOOP_and_14_itm & and_317_m1c) | (COMP_LOOP_COMP_LOOP_and_13_itm
      & and_320_m1c) | (COMP_LOOP_COMP_LOOP_and_12_itm & and_322_m1c) | (COMP_LOOP_COMP_LOOP_and_11_itm
      & and_324_m1c) | (COMP_LOOP_COMP_LOOP_and_10_itm & and_327_m1c) | (COMP_LOOP_COMP_LOOP_and_9_itm
      & and_329_m1c) | (COMP_LOOP_COMP_LOOP_and_8_itm & and_331_m1c) | (COMP_LOOP_COMP_LOOP_and_68_itm
      & and_334_m1c) | (COMP_LOOP_COMP_LOOP_and_6_itm & and_336_m1c) | (COMP_LOOP_COMP_LOOP_and_5_itm
      & and_339_m1c);
  assign COMP_LOOP_or_14_nl = (COMP_LOOP_COMP_LOOP_and_5_itm & and_dcpl_283) | (COMP_LOOP_COMP_LOOP_and_4_itm
      & and_305_m1c) | (COMP_LOOP_COMP_LOOP_and_64_itm & and_307_m1c) | (COMP_LOOP_COMP_LOOP_and_2_itm
      & and_309_m1c) | (COMP_LOOP_COMP_LOOP_and_62_itm & and_312_m1c) | (COMP_LOOP_COMP_LOOP_and_305_itm
      & and_315_m1c) | (COMP_LOOP_COMP_LOOP_nor_itm & and_317_m1c) | (COMP_LOOP_COMP_LOOP_and_14_itm
      & and_320_m1c) | (COMP_LOOP_COMP_LOOP_and_13_itm & and_322_m1c) | (COMP_LOOP_COMP_LOOP_and_12_itm
      & and_324_m1c) | (COMP_LOOP_COMP_LOOP_and_11_itm & and_327_m1c) | (COMP_LOOP_COMP_LOOP_and_10_itm
      & and_329_m1c) | (COMP_LOOP_COMP_LOOP_and_9_itm & and_331_m1c) | (COMP_LOOP_COMP_LOOP_and_8_itm
      & and_334_m1c) | (COMP_LOOP_COMP_LOOP_and_68_itm & and_336_m1c) | (COMP_LOOP_COMP_LOOP_and_6_itm
      & and_339_m1c);
  assign COMP_LOOP_or_15_nl = (COMP_LOOP_COMP_LOOP_and_6_itm & and_dcpl_283) | (COMP_LOOP_COMP_LOOP_and_5_itm
      & and_305_m1c) | (COMP_LOOP_COMP_LOOP_and_4_itm & and_307_m1c) | (COMP_LOOP_COMP_LOOP_and_64_itm
      & and_309_m1c) | (COMP_LOOP_COMP_LOOP_and_2_itm & and_312_m1c) | (COMP_LOOP_COMP_LOOP_and_62_itm
      & and_315_m1c) | (COMP_LOOP_COMP_LOOP_and_305_itm & and_317_m1c) | (COMP_LOOP_COMP_LOOP_nor_itm
      & and_320_m1c) | (COMP_LOOP_COMP_LOOP_and_14_itm & and_322_m1c) | (COMP_LOOP_COMP_LOOP_and_13_itm
      & and_324_m1c) | (COMP_LOOP_COMP_LOOP_and_12_itm & and_327_m1c) | (COMP_LOOP_COMP_LOOP_and_11_itm
      & and_329_m1c) | (COMP_LOOP_COMP_LOOP_and_10_itm & and_331_m1c) | (COMP_LOOP_COMP_LOOP_and_9_itm
      & and_334_m1c) | (COMP_LOOP_COMP_LOOP_and_8_itm & and_336_m1c) | (COMP_LOOP_COMP_LOOP_and_68_itm
      & and_339_m1c);
  assign COMP_LOOP_or_16_nl = (COMP_LOOP_COMP_LOOP_and_68_itm & and_dcpl_283) | (COMP_LOOP_COMP_LOOP_and_6_itm
      & and_305_m1c) | (COMP_LOOP_COMP_LOOP_and_5_itm & and_307_m1c) | (COMP_LOOP_COMP_LOOP_and_4_itm
      & and_309_m1c) | (COMP_LOOP_COMP_LOOP_and_64_itm & and_312_m1c) | (COMP_LOOP_COMP_LOOP_and_2_itm
      & and_315_m1c) | (COMP_LOOP_COMP_LOOP_and_62_itm & and_317_m1c) | (COMP_LOOP_COMP_LOOP_and_305_itm
      & and_320_m1c) | (COMP_LOOP_COMP_LOOP_nor_itm & and_322_m1c) | (COMP_LOOP_COMP_LOOP_and_14_itm
      & and_324_m1c) | (COMP_LOOP_COMP_LOOP_and_13_itm & and_327_m1c) | (COMP_LOOP_COMP_LOOP_and_12_itm
      & and_329_m1c) | (COMP_LOOP_COMP_LOOP_and_11_itm & and_331_m1c) | (COMP_LOOP_COMP_LOOP_and_10_itm
      & and_334_m1c) | (COMP_LOOP_COMP_LOOP_and_9_itm & and_336_m1c) | (COMP_LOOP_COMP_LOOP_and_8_itm
      & and_339_m1c);
  assign COMP_LOOP_or_17_nl = (COMP_LOOP_COMP_LOOP_and_8_itm & and_dcpl_283) | (COMP_LOOP_COMP_LOOP_and_68_itm
      & and_305_m1c) | (COMP_LOOP_COMP_LOOP_and_6_itm & and_307_m1c) | (COMP_LOOP_COMP_LOOP_and_5_itm
      & and_309_m1c) | (COMP_LOOP_COMP_LOOP_and_4_itm & and_312_m1c) | (COMP_LOOP_COMP_LOOP_and_64_itm
      & and_315_m1c) | (COMP_LOOP_COMP_LOOP_and_2_itm & and_317_m1c) | (COMP_LOOP_COMP_LOOP_and_62_itm
      & and_320_m1c) | (COMP_LOOP_COMP_LOOP_and_305_itm & and_322_m1c) | (COMP_LOOP_COMP_LOOP_nor_itm
      & and_324_m1c) | (COMP_LOOP_COMP_LOOP_and_14_itm & and_327_m1c) | (COMP_LOOP_COMP_LOOP_and_13_itm
      & and_329_m1c) | (COMP_LOOP_COMP_LOOP_and_12_itm & and_331_m1c) | (COMP_LOOP_COMP_LOOP_and_11_itm
      & and_334_m1c) | (COMP_LOOP_COMP_LOOP_and_10_itm & and_336_m1c) | (COMP_LOOP_COMP_LOOP_and_9_itm
      & and_339_m1c);
  assign COMP_LOOP_or_18_nl = (COMP_LOOP_COMP_LOOP_and_9_itm & and_dcpl_283) | (COMP_LOOP_COMP_LOOP_and_8_itm
      & and_305_m1c) | (COMP_LOOP_COMP_LOOP_and_68_itm & and_307_m1c) | (COMP_LOOP_COMP_LOOP_and_6_itm
      & and_309_m1c) | (COMP_LOOP_COMP_LOOP_and_5_itm & and_312_m1c) | (COMP_LOOP_COMP_LOOP_and_4_itm
      & and_315_m1c) | (COMP_LOOP_COMP_LOOP_and_64_itm & and_317_m1c) | (COMP_LOOP_COMP_LOOP_and_2_itm
      & and_320_m1c) | (COMP_LOOP_COMP_LOOP_and_62_itm & and_322_m1c) | (COMP_LOOP_COMP_LOOP_and_305_itm
      & and_324_m1c) | (COMP_LOOP_COMP_LOOP_nor_itm & and_327_m1c) | (COMP_LOOP_COMP_LOOP_and_14_itm
      & and_329_m1c) | (COMP_LOOP_COMP_LOOP_and_13_itm & and_331_m1c) | (COMP_LOOP_COMP_LOOP_and_12_itm
      & and_334_m1c) | (COMP_LOOP_COMP_LOOP_and_11_itm & and_336_m1c) | (COMP_LOOP_COMP_LOOP_and_10_itm
      & and_339_m1c);
  assign COMP_LOOP_or_19_nl = (COMP_LOOP_COMP_LOOP_and_10_itm & and_dcpl_283) | (COMP_LOOP_COMP_LOOP_and_9_itm
      & and_305_m1c) | (COMP_LOOP_COMP_LOOP_and_8_itm & and_307_m1c) | (COMP_LOOP_COMP_LOOP_and_68_itm
      & and_309_m1c) | (COMP_LOOP_COMP_LOOP_and_6_itm & and_312_m1c) | (COMP_LOOP_COMP_LOOP_and_5_itm
      & and_315_m1c) | (COMP_LOOP_COMP_LOOP_and_4_itm & and_317_m1c) | (COMP_LOOP_COMP_LOOP_and_64_itm
      & and_320_m1c) | (COMP_LOOP_COMP_LOOP_and_2_itm & and_322_m1c) | (COMP_LOOP_COMP_LOOP_and_62_itm
      & and_324_m1c) | (COMP_LOOP_COMP_LOOP_and_305_itm & and_327_m1c) | (COMP_LOOP_COMP_LOOP_nor_itm
      & and_329_m1c) | (COMP_LOOP_COMP_LOOP_and_14_itm & and_331_m1c) | (COMP_LOOP_COMP_LOOP_and_13_itm
      & and_334_m1c) | (COMP_LOOP_COMP_LOOP_and_12_itm & and_336_m1c) | (COMP_LOOP_COMP_LOOP_and_11_itm
      & and_339_m1c);
  assign COMP_LOOP_or_20_nl = (COMP_LOOP_COMP_LOOP_and_11_itm & and_dcpl_283) | (COMP_LOOP_COMP_LOOP_and_10_itm
      & and_305_m1c) | (COMP_LOOP_COMP_LOOP_and_9_itm & and_307_m1c) | (COMP_LOOP_COMP_LOOP_and_8_itm
      & and_309_m1c) | (COMP_LOOP_COMP_LOOP_and_68_itm & and_312_m1c) | (COMP_LOOP_COMP_LOOP_and_6_itm
      & and_315_m1c) | (COMP_LOOP_COMP_LOOP_and_5_itm & and_317_m1c) | (COMP_LOOP_COMP_LOOP_and_4_itm
      & and_320_m1c) | (COMP_LOOP_COMP_LOOP_and_64_itm & and_322_m1c) | (COMP_LOOP_COMP_LOOP_and_2_itm
      & and_324_m1c) | (COMP_LOOP_COMP_LOOP_and_62_itm & and_327_m1c) | (COMP_LOOP_COMP_LOOP_and_305_itm
      & and_329_m1c) | (COMP_LOOP_COMP_LOOP_nor_itm & and_331_m1c) | (COMP_LOOP_COMP_LOOP_and_14_itm
      & and_334_m1c) | (COMP_LOOP_COMP_LOOP_and_13_itm & and_336_m1c) | (COMP_LOOP_COMP_LOOP_and_12_itm
      & and_339_m1c);
  assign COMP_LOOP_or_21_nl = (COMP_LOOP_COMP_LOOP_and_12_itm & and_dcpl_283) | (COMP_LOOP_COMP_LOOP_and_11_itm
      & and_305_m1c) | (COMP_LOOP_COMP_LOOP_and_10_itm & and_307_m1c) | (COMP_LOOP_COMP_LOOP_and_9_itm
      & and_309_m1c) | (COMP_LOOP_COMP_LOOP_and_8_itm & and_312_m1c) | (COMP_LOOP_COMP_LOOP_and_68_itm
      & and_315_m1c) | (COMP_LOOP_COMP_LOOP_and_6_itm & and_317_m1c) | (COMP_LOOP_COMP_LOOP_and_5_itm
      & and_320_m1c) | (COMP_LOOP_COMP_LOOP_and_4_itm & and_322_m1c) | (COMP_LOOP_COMP_LOOP_and_64_itm
      & and_324_m1c) | (COMP_LOOP_COMP_LOOP_and_2_itm & and_327_m1c) | (COMP_LOOP_COMP_LOOP_and_62_itm
      & and_329_m1c) | (COMP_LOOP_COMP_LOOP_and_305_itm & and_331_m1c) | (COMP_LOOP_COMP_LOOP_nor_itm
      & and_334_m1c) | (COMP_LOOP_COMP_LOOP_and_14_itm & and_336_m1c) | (COMP_LOOP_COMP_LOOP_and_13_itm
      & and_339_m1c);
  assign COMP_LOOP_or_22_nl = (COMP_LOOP_COMP_LOOP_and_13_itm & and_dcpl_283) | (COMP_LOOP_COMP_LOOP_and_12_itm
      & and_305_m1c) | (COMP_LOOP_COMP_LOOP_and_11_itm & and_307_m1c) | (COMP_LOOP_COMP_LOOP_and_10_itm
      & and_309_m1c) | (COMP_LOOP_COMP_LOOP_and_9_itm & and_312_m1c) | (COMP_LOOP_COMP_LOOP_and_8_itm
      & and_315_m1c) | (COMP_LOOP_COMP_LOOP_and_68_itm & and_317_m1c) | (COMP_LOOP_COMP_LOOP_and_6_itm
      & and_320_m1c) | (COMP_LOOP_COMP_LOOP_and_5_itm & and_322_m1c) | (COMP_LOOP_COMP_LOOP_and_4_itm
      & and_324_m1c) | (COMP_LOOP_COMP_LOOP_and_64_itm & and_327_m1c) | (COMP_LOOP_COMP_LOOP_and_2_itm
      & and_329_m1c) | (COMP_LOOP_COMP_LOOP_and_62_itm & and_331_m1c) | (COMP_LOOP_COMP_LOOP_and_305_itm
      & and_334_m1c) | (COMP_LOOP_COMP_LOOP_nor_itm & and_336_m1c) | (COMP_LOOP_COMP_LOOP_and_14_itm
      & and_339_m1c);
  assign COMP_LOOP_or_23_nl = (COMP_LOOP_COMP_LOOP_and_14_itm & and_dcpl_283) | (COMP_LOOP_COMP_LOOP_and_13_itm
      & and_305_m1c) | (COMP_LOOP_COMP_LOOP_and_12_itm & and_307_m1c) | (COMP_LOOP_COMP_LOOP_and_11_itm
      & and_309_m1c) | (COMP_LOOP_COMP_LOOP_and_10_itm & and_312_m1c) | (COMP_LOOP_COMP_LOOP_and_9_itm
      & and_315_m1c) | (COMP_LOOP_COMP_LOOP_and_8_itm & and_317_m1c) | (COMP_LOOP_COMP_LOOP_and_68_itm
      & and_320_m1c) | (COMP_LOOP_COMP_LOOP_and_6_itm & and_322_m1c) | (COMP_LOOP_COMP_LOOP_and_5_itm
      & and_324_m1c) | (COMP_LOOP_COMP_LOOP_and_4_itm & and_327_m1c) | (COMP_LOOP_COMP_LOOP_and_64_itm
      & and_329_m1c) | (COMP_LOOP_COMP_LOOP_and_2_itm & and_331_m1c) | (COMP_LOOP_COMP_LOOP_and_62_itm
      & and_334_m1c) | (COMP_LOOP_COMP_LOOP_and_305_itm & and_336_m1c) | (COMP_LOOP_COMP_LOOP_nor_itm
      & and_339_m1c);
  assign nor_716_nl = ~((fsm_output[6]) | and_dcpl_124);
  assign mux_2736_nl = MUX_s_1_2_2(nor_716_nl, mux_tmp_2687, fsm_output[7]);
  assign mux_2734_nl = MUX_s_1_2_2(and_dcpl_109, nor_tmp_9, fsm_output[6]);
  assign mux_2735_nl = MUX_s_1_2_2(mux_2734_nl, (fsm_output[6]), fsm_output[7]);
  assign mux_2737_nl = MUX_s_1_2_2(mux_2736_nl, mux_2735_nl, fsm_output[5]);
  assign or_3268_nl = (fsm_output[6]) | and_dcpl_123;
  assign mux_2731_nl = MUX_s_1_2_2(nor_tmp_6, (~ nor_tmp_288), fsm_output[6]);
  assign mux_2732_nl = MUX_s_1_2_2(or_3268_nl, mux_2731_nl, fsm_output[7]);
  assign mux_2729_nl = MUX_s_1_2_2(or_tmp_2483, (~ or_tmp_2233), fsm_output[6]);
  assign mux_2730_nl = MUX_s_1_2_2(mux_2729_nl, nand_tmp_119, fsm_output[7]);
  assign mux_2733_nl = MUX_s_1_2_2(mux_2732_nl, mux_2730_nl, fsm_output[5]);
  assign mux_2738_nl = MUX_s_1_2_2((~ mux_2737_nl), mux_2733_nl, fsm_output[2]);
  assign mux_55_nl = MUX_s_1_2_2((~ (fsm_output[6])), or_tmp_3, fsm_output[7]);
  assign mux_2724_nl = MUX_s_1_2_2((~ nor_tmp_300), or_tmp_9, fsm_output[6]);
  assign mux_2725_nl = MUX_s_1_2_2(mux_2724_nl, (fsm_output[6]), fsm_output[7]);
  assign mux_2727_nl = MUX_s_1_2_2(mux_55_nl, mux_2725_nl, fsm_output[5]);
  assign mux_2722_nl = MUX_s_1_2_2((~ (fsm_output[6])), nand_tmp_93, fsm_output[7]);
  assign mux_50_nl = MUX_s_1_2_2(or_36_cse, (fsm_output[6]), fsm_output[7]);
  assign mux_2723_nl = MUX_s_1_2_2(mux_2722_nl, mux_50_nl, fsm_output[5]);
  assign mux_2728_nl = MUX_s_1_2_2(mux_2727_nl, mux_2723_nl, fsm_output[2]);
  assign mux_2739_nl = MUX_s_1_2_2(mux_2738_nl, mux_2728_nl, fsm_output[8]);
  assign mux_2717_nl = MUX_s_1_2_2(and_dcpl_243, mux_tmp_2696, fsm_output[7]);
  assign mux_2718_nl = MUX_s_1_2_2((~ mux_2717_nl), mux_tmp_2701, fsm_output[5]);
  assign mux_2715_nl = MUX_s_1_2_2(and_dcpl_243, or_tmp_2479, fsm_output[7]);
  assign mux_2716_nl = MUX_s_1_2_2((~ mux_2715_nl), mux_tmp_2698, fsm_output[5]);
  assign mux_2719_nl = MUX_s_1_2_2(mux_2718_nl, mux_2716_nl, fsm_output[2]);
  assign nand_118_nl = ~((fsm_output[6]) & (~ nor_tmp_6));
  assign mux_2712_nl = MUX_s_1_2_2(nand_118_nl, or_tmp_434, fsm_output[7]);
  assign or_3269_nl = (fsm_output[6]) | (~ or_tmp_2248);
  assign mux_2710_nl = MUX_s_1_2_2(nor_tmp_291, (~ nor_tmp_6), fsm_output[6]);
  assign mux_2711_nl = MUX_s_1_2_2(or_3269_nl, mux_2710_nl, fsm_output[7]);
  assign mux_2713_nl = MUX_s_1_2_2(mux_2712_nl, mux_2711_nl, fsm_output[5]);
  assign or_2540_nl = (fsm_output[6]) | (~ or_tmp_2253);
  assign mux_2708_nl = MUX_s_1_2_2(or_tmp_4, or_2540_nl, fsm_output[7]);
  assign mux_2706_nl = MUX_s_1_2_2(nor_tmp_6, (~ nor_tmp_9), fsm_output[6]);
  assign mux_2707_nl = MUX_s_1_2_2(or_tmp_2479, mux_2706_nl, fsm_output[7]);
  assign mux_2709_nl = MUX_s_1_2_2(mux_2708_nl, mux_2707_nl, fsm_output[5]);
  assign mux_2714_nl = MUX_s_1_2_2(mux_2713_nl, mux_2709_nl, fsm_output[2]);
  assign mux_2720_nl = MUX_s_1_2_2(mux_2719_nl, mux_2714_nl, fsm_output[8]);
  assign mux_2740_nl = MUX_s_1_2_2(mux_2739_nl, mux_2720_nl, fsm_output[4]);
  assign mux_29_nl = MUX_s_1_2_2(mux_28_cse, or_tmp_14, fsm_output[7]);
  assign mux_2702_nl = MUX_s_1_2_2(mux_tmp_2701, mux_29_nl, fsm_output[5]);
  assign mux_2697_nl = MUX_s_1_2_2(mux_tmp_2696, or_tmp_14, fsm_output[7]);
  assign mux_2699_nl = MUX_s_1_2_2(mux_tmp_2698, mux_2697_nl, fsm_output[5]);
  assign mux_2703_nl = MUX_s_1_2_2(mux_2702_nl, mux_2699_nl, fsm_output[2]);
  assign or_25_nl = (~((fsm_output[7:6]!=2'b01))) | (fsm_output[10]);
  assign or_24_nl = nor_223_cse | (fsm_output[10]);
  assign mux_22_nl = MUX_s_1_2_2(or_25_nl, or_24_nl, fsm_output[5]);
  assign mux_2704_nl = MUX_s_1_2_2(mux_2703_nl, mux_22_nl, fsm_output[8]);
  assign nand_116_nl = ~((fsm_output[6]) & (~ and_dcpl_240));
  assign mux_2691_nl = MUX_s_1_2_2(nand_116_nl, or_tmp_2474, fsm_output[7]);
  assign mux_17_nl = MUX_s_1_2_2((fsm_output[6]), or_tmp_8, fsm_output[7]);
  assign mux_2692_nl = MUX_s_1_2_2(mux_2691_nl, mux_17_nl, fsm_output[5]);
  assign mux_2688_nl = MUX_s_1_2_2(mux_tmp_2687, or_tmp_14, fsm_output[7]);
  assign or_18_nl = (~((~ (fsm_output[6])) | (fsm_output[3]) | (fsm_output[1])))
      | (fsm_output[10]);
  assign mux_13_nl = MUX_s_1_2_2((fsm_output[6]), or_18_nl, fsm_output[7]);
  assign mux_2689_nl = MUX_s_1_2_2(mux_2688_nl, mux_13_nl, fsm_output[5]);
  assign mux_2693_nl = MUX_s_1_2_2(mux_2692_nl, mux_2689_nl, fsm_output[2]);
  assign mux_10_nl = MUX_s_1_2_2(mux_9_cse, or_15_cse, fsm_output[7]);
  assign mux_8_nl = MUX_s_1_2_2(mux_7_cse, or_tmp_4, fsm_output[7]);
  assign mux_11_nl = MUX_s_1_2_2(mux_10_nl, mux_8_nl, fsm_output[5]);
  assign mux_2677_nl = MUX_s_1_2_2(or_tmp_2230, (fsm_output[10]), fsm_output[6]);
  assign mux_2678_nl = MUX_s_1_2_2(or_tmp_8, mux_2677_nl, fsm_output[7]);
  assign mux_2679_nl = MUX_s_1_2_2(mux_2678_nl, mux_3_cse, fsm_output[5]);
  assign mux_2685_nl = MUX_s_1_2_2(mux_11_nl, mux_2679_nl, fsm_output[2]);
  assign mux_2694_nl = MUX_s_1_2_2(mux_2693_nl, mux_2685_nl, fsm_output[8]);
  assign mux_2705_nl = MUX_s_1_2_2(mux_2704_nl, mux_2694_nl, fsm_output[4]);
  assign and_340_nl = and_dcpl_191 & and_dcpl_98;
  assign COMP_LOOP_or_30_nl = ((~ (modulo_result_rem_cmp_z[63])) & and_345_m1c) |
      (not_tmp_634 & (~ (modulo_result_rem_cmp_z[63])));
  assign COMP_LOOP_or_31_nl = ((modulo_result_rem_cmp_z[63]) & and_345_m1c) | (not_tmp_634
      & (modulo_result_rem_cmp_z[63]));
  assign COMP_LOOP_and_277_nl = COMP_LOOP_COMP_LOOP_nor_1_itm & mux_2770_m1c;
  assign COMP_LOOP_COMP_LOOP_and_932_nl = (COMP_LOOP_acc_10_cse_12_1_1_sva[0]) &
      COMP_LOOP_nor_11_itm & mux_2770_m1c;
  assign COMP_LOOP_COMP_LOOP_and_934_nl = (COMP_LOOP_acc_10_cse_12_1_1_sva[1]) &
      COMP_LOOP_nor_12_itm & mux_2770_m1c;
  assign COMP_LOOP_and_1_nl = COMP_LOOP_COMP_LOOP_and_137_itm & mux_2770_m1c;
  assign COMP_LOOP_COMP_LOOP_and_936_nl = (COMP_LOOP_acc_10_cse_12_1_1_sva[2]) &
      COMP_LOOP_nor_134_itm & mux_2770_m1c;
  assign COMP_LOOP_and_2_nl = COMP_LOOP_COMP_LOOP_and_139_itm & mux_2770_m1c;
  assign COMP_LOOP_and_3_nl = COMP_LOOP_COMP_LOOP_and_140_itm & mux_2770_m1c;
  assign COMP_LOOP_and_4_nl = COMP_LOOP_COMP_LOOP_and_141_itm & mux_2770_m1c;
  assign COMP_LOOP_COMP_LOOP_and_930_nl = (COMP_LOOP_acc_10_cse_12_1_1_sva[3]) &
      COMP_LOOP_nor_137_itm & mux_2770_m1c;
  assign COMP_LOOP_and_5_nl = COMP_LOOP_COMP_LOOP_and_143_itm & mux_2770_m1c;
  assign COMP_LOOP_and_6_nl = COMP_LOOP_COMP_LOOP_and_144_itm & mux_2770_m1c;
  assign COMP_LOOP_and_7_nl = COMP_LOOP_COMP_LOOP_and_145_itm & mux_2770_m1c;
  assign COMP_LOOP_and_8_nl = COMP_LOOP_COMP_LOOP_and_146_itm & mux_2770_m1c;
  assign COMP_LOOP_and_9_nl = COMP_LOOP_COMP_LOOP_and_147_itm & mux_2770_m1c;
  assign COMP_LOOP_and_10_nl = COMP_LOOP_COMP_LOOP_and_148_itm & mux_2770_m1c;
  assign COMP_LOOP_and_11_nl = COMP_LOOP_COMP_LOOP_and_149_itm & mux_2770_m1c;
  assign nor_1265_nl = ~((~ (fsm_output[2])) | (~ (fsm_output[8])) | (~ (fsm_output[7]))
      | (fsm_output[0]) | (fsm_output[3]) | (~ (fsm_output[9])) | (fsm_output[5])
      | (fsm_output[10]));
  assign nor_1266_nl = ~((fsm_output[2]) | (~ (fsm_output[8])) | (fsm_output[7])
      | (fsm_output[0]) | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[5])
      | (~ (fsm_output[10])));
  assign mux_112_nl = MUX_s_1_2_2(nor_1265_nl, nor_1266_nl, fsm_output[4]);
  assign or_113_nl = (~ (fsm_output[7])) | (~ (fsm_output[0])) | (fsm_output[3])
      | (fsm_output[9]) | (fsm_output[5]) | (fsm_output[10]);
  assign nand_395_nl = ~((fsm_output[7]) & (fsm_output[0]) & (fsm_output[3]) & (fsm_output[9])
      & (fsm_output[5]) & (~ (fsm_output[10])));
  assign mux_110_nl = MUX_s_1_2_2(or_113_nl, nand_395_nl, fsm_output[8]);
  assign nor_1267_nl = ~((fsm_output[2]) | mux_110_nl);
  assign nor_1268_nl = ~((~ (fsm_output[8])) | (~ (fsm_output[7])) | (fsm_output[0])
      | (fsm_output[3]) | (fsm_output[9]) | (~ (fsm_output[5])) | (fsm_output[10]));
  assign or_109_nl = (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[5]) | (fsm_output[10]);
  assign or_108_nl = (fsm_output[3]) | (~ (fsm_output[9])) | (fsm_output[5]) | (fsm_output[10]);
  assign mux_107_nl = MUX_s_1_2_2(or_109_nl, or_108_nl, fsm_output[0]);
  assign nor_1269_nl = ~((fsm_output[7]) | mux_107_nl);
  assign nor_1270_nl = ~((fsm_output[7]) | (~ (fsm_output[0])) | (~ (fsm_output[3]))
      | (fsm_output[9]) | not_tmp_45);
  assign mux_108_nl = MUX_s_1_2_2(nor_1269_nl, nor_1270_nl, fsm_output[8]);
  assign mux_109_nl = MUX_s_1_2_2(nor_1268_nl, mux_108_nl, fsm_output[2]);
  assign mux_111_nl = MUX_s_1_2_2(nor_1267_nl, mux_109_nl, fsm_output[4]);
  assign mux_113_nl = MUX_s_1_2_2(mux_112_nl, mux_111_nl, fsm_output[6]);
  assign nor_1271_nl = ~((~ (fsm_output[8])) | (~ (fsm_output[7])) | (~ (fsm_output[0]))
      | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[5]) | (fsm_output[10]));
  assign nor_1272_nl = ~((~ (fsm_output[8])) | (fsm_output[7]) | (fsm_output[0])
      | (fsm_output[3]) | (fsm_output[9]) | (~ (fsm_output[5])) | (fsm_output[10]));
  assign mux_104_nl = MUX_s_1_2_2(nor_1271_nl, nor_1272_nl, fsm_output[2]);
  assign and_795_nl = (fsm_output[3]) & (fsm_output[9]) & (fsm_output[5]) & (~ (fsm_output[10]));
  assign nor_1273_nl = ~((fsm_output[3]) | (fsm_output[9]) | not_tmp_45);
  assign mux_102_nl = MUX_s_1_2_2(and_795_nl, nor_1273_nl, fsm_output[0]);
  assign and_794_nl = (~((fsm_output[8:7]!=2'b01))) & mux_102_nl;
  assign nor_1274_nl = ~((~ (fsm_output[8])) | (fsm_output[7]) | (~ (fsm_output[0]))
      | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[5]) | (fsm_output[10]));
  assign mux_103_nl = MUX_s_1_2_2(and_794_nl, nor_1274_nl, fsm_output[2]);
  assign mux_105_nl = MUX_s_1_2_2(mux_104_nl, mux_103_nl, fsm_output[4]);
  assign or_98_nl = (~ (fsm_output[8])) | (~ (fsm_output[7])) | (fsm_output[0]) |
      (fsm_output[3]) | (fsm_output[9]) | not_tmp_45;
  assign or_95_nl = (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[5]) | (~
      (fsm_output[10]));
  assign or_93_nl = (fsm_output[3]) | (~ (fsm_output[9])) | (fsm_output[5]) | (~
      (fsm_output[10]));
  assign mux_100_nl = MUX_s_1_2_2(or_95_nl, or_93_nl, fsm_output[0]);
  assign or_96_nl = (fsm_output[8:7]!=2'b00) | mux_100_nl;
  assign mux_101_nl = MUX_s_1_2_2(or_98_nl, or_96_nl, fsm_output[2]);
  assign nor_1275_nl = ~((fsm_output[4]) | mux_101_nl);
  assign mux_106_nl = MUX_s_1_2_2(mux_105_nl, nor_1275_nl, fsm_output[6]);
  assign mux_114_nl = MUX_s_1_2_2(mux_113_nl, mux_106_nl, fsm_output[1]);
  assign nor_1303_nl = ~((~ (fsm_output[3])) | (fsm_output[0]) | (~ (fsm_output[1]))
      | (fsm_output[10]));
  assign mux_2862_nl = MUX_s_1_2_2(nor_1303_nl, (fsm_output[10]), fsm_output[6]);
  assign mux_2863_nl = MUX_s_1_2_2((~ mux_2862_nl), mux_tmp_2796, fsm_output[7]);
  assign mux_2861_nl = MUX_s_1_2_2(or_tmp_4, or_tmp_434, fsm_output[7]);
  assign mux_2864_nl = MUX_s_1_2_2(mux_2863_nl, mux_2861_nl, fsm_output[5]);
  assign mux_2858_nl = MUX_s_1_2_2(and_dcpl_109, (fsm_output[10]), and_573_cse);
  assign and_506_nl = (fsm_output[6]) & mux_2858_nl;
  assign and_508_nl = (fsm_output[6]) & (~ nor_tmp_9);
  assign mux_2859_nl = MUX_s_1_2_2(and_506_nl, and_508_nl, fsm_output[7]);
  assign or_2643_nl = (~ (fsm_output[0])) | (fsm_output[1]) | (fsm_output[3]) | (~
      (fsm_output[10]));
  assign mux_2856_nl = MUX_s_1_2_2(or_2643_nl, or_tmp_2253, fsm_output[6]);
  assign mux_2855_nl = MUX_s_1_2_2(or_tmp_21, nor_tmp_300, fsm_output[6]);
  assign mux_2857_nl = MUX_s_1_2_2((~ mux_2856_nl), mux_2855_nl, fsm_output[7]);
  assign mux_2860_nl = MUX_s_1_2_2(mux_2859_nl, mux_2857_nl, fsm_output[5]);
  assign mux_2865_nl = MUX_s_1_2_2((~ mux_2864_nl), mux_2860_nl, fsm_output[2]);
  assign mux_2852_nl = MUX_s_1_2_2(or_tmp_2293, or_tmp_2280, fsm_output[7]);
  assign mux_2849_nl = MUX_s_1_2_2(nor_tmp_6, mux_tmp_2239, nor_412_cse);
  assign mux_2850_nl = MUX_s_1_2_2((~ and_dcpl_240), mux_2849_nl, fsm_output[6]);
  assign and_346_nl = (fsm_output[6]) & (and_573_cse | (fsm_output[3]) | (~ (fsm_output[10])));
  assign mux_2851_nl = MUX_s_1_2_2(mux_2850_nl, and_346_nl, fsm_output[7]);
  assign mux_2853_nl = MUX_s_1_2_2((~ mux_2852_nl), mux_2851_nl, fsm_output[5]);
  assign mux_2846_nl = MUX_s_1_2_2((~ nor_tmp_300), mux_tmp_2800, fsm_output[6]);
  assign mux_2847_nl = MUX_s_1_2_2(and_dcpl_243, mux_2846_nl, fsm_output[7]);
  assign mux_2844_nl = MUX_s_1_2_2((~ mux_tmp_2362), nor_tmp_6, fsm_output[6]);
  assign mux_2845_nl = MUX_s_1_2_2(mux_2844_nl, and_tmp_16, fsm_output[7]);
  assign mux_2848_nl = MUX_s_1_2_2(mux_2847_nl, mux_2845_nl, fsm_output[5]);
  assign mux_2854_nl = MUX_s_1_2_2(mux_2853_nl, mux_2848_nl, fsm_output[2]);
  assign mux_2866_nl = MUX_s_1_2_2(mux_2865_nl, mux_2854_nl, fsm_output[8]);
  assign mux_2840_nl = MUX_s_1_2_2(not_tmp_378, mux_tmp_2813, fsm_output[7]);
  assign or_2639_nl = (fsm_output[6]) | (~ mux_tmp_2800);
  assign or_2638_nl = (fsm_output[6]) | (~ or_tmp_2289);
  assign mux_2839_nl = MUX_s_1_2_2(or_2639_nl, or_2638_nl, fsm_output[7]);
  assign mux_2841_nl = MUX_s_1_2_2(mux_2840_nl, mux_2839_nl, fsm_output[5]);
  assign or_2637_nl = (fsm_output[6]) | (~ and_dcpl_240);
  assign mux_2837_nl = MUX_s_1_2_2(not_tmp_426, or_2637_nl, fsm_output[7]);
  assign or_2636_nl = (~ (fsm_output[0])) | (fsm_output[1]) | (~ (fsm_output[3]))
      | (fsm_output[10]);
  assign mux_2835_nl = MUX_s_1_2_2((~ nand_402_cse), or_2636_nl, fsm_output[6]);
  assign mux_2836_nl = MUX_s_1_2_2(or_36_cse, mux_2835_nl, fsm_output[7]);
  assign mux_2838_nl = MUX_s_1_2_2(mux_2837_nl, mux_2836_nl, fsm_output[5]);
  assign mux_2842_nl = MUX_s_1_2_2(mux_2841_nl, mux_2838_nl, fsm_output[2]);
  assign or_3347_nl = (fsm_output[6]) | (~((fsm_output[1:0]!=2'b00) | (~ mux_tmp_2239)));
  assign mux_2831_nl = MUX_s_1_2_2((fsm_output[10]), (~ or_tmp_2233), fsm_output[6]);
  assign mux_2832_nl = MUX_s_1_2_2(or_3347_nl, mux_2831_nl, fsm_output[7]);
  assign mux_2829_nl = MUX_s_1_2_2(or_tmp_21, mux_tmp_2254, fsm_output[6]);
  assign or_2632_nl = (fsm_output[1:0]!=2'b01) | (~ nor_tmp_6);
  assign mux_2828_nl = MUX_s_1_2_2(or_2632_nl, mux_tmp_2250, fsm_output[6]);
  assign mux_2830_nl = MUX_s_1_2_2(mux_2829_nl, mux_2828_nl, fsm_output[7]);
  assign mux_2833_nl = MUX_s_1_2_2(mux_2832_nl, mux_2830_nl, fsm_output[5]);
  assign mux_2825_nl = MUX_s_1_2_2(and_dcpl_110, or_tmp_2483, fsm_output[6]);
  assign mux_2826_nl = MUX_s_1_2_2(mux_2825_nl, (~ mux_tmp_2349), fsm_output[7]);
  assign mux_2823_nl = MUX_s_1_2_2(and_dcpl_101, or_tmp_2266, fsm_output[6]);
  assign mux_2824_nl = MUX_s_1_2_2((~ mux_2823_nl), or_tmp_4, fsm_output[7]);
  assign mux_2827_nl = MUX_s_1_2_2(mux_2826_nl, mux_2824_nl, fsm_output[5]);
  assign mux_2834_nl = MUX_s_1_2_2(mux_2833_nl, mux_2827_nl, fsm_output[2]);
  assign mux_2843_nl = MUX_s_1_2_2(mux_2842_nl, mux_2834_nl, fsm_output[8]);
  assign mux_2867_nl = MUX_s_1_2_2((~ mux_2866_nl), mux_2843_nl, fsm_output[4]);
  assign nor_680_nl = ~((fsm_output[6]) | and_dcpl_102);
  assign mux_2818_nl = MUX_s_1_2_2(nor_680_nl, or_tmp_4, fsm_output[7]);
  assign mux_2817_nl = MUX_s_1_2_2(or_tmp_3, or_tmp_2246, fsm_output[7]);
  assign mux_2819_nl = MUX_s_1_2_2(mux_2818_nl, mux_2817_nl, fsm_output[5]);
  assign mux_2815_nl = MUX_s_1_2_2(not_tmp_463, or_tmp_3, fsm_output[7]);
  assign mux_2814_nl = MUX_s_1_2_2(mux_tmp_2813, or_tmp_2474, fsm_output[7]);
  assign mux_2816_nl = MUX_s_1_2_2(mux_2815_nl, mux_2814_nl, fsm_output[5]);
  assign mux_2820_nl = MUX_s_1_2_2(mux_2819_nl, mux_2816_nl, fsm_output[2]);
  assign or_2629_nl = (~((fsm_output[3]) | (~ (fsm_output[1])))) | (fsm_output[10]);
  assign mux_2809_nl = MUX_s_1_2_2(or_2629_nl, or_tmp_2238, fsm_output[6]);
  assign mux_2810_nl = MUX_s_1_2_2(or_tmp_2276, mux_2809_nl, fsm_output[7]);
  assign nand_128_nl = ~((fsm_output[6]) & (~((~((fsm_output[1]) | (~ (fsm_output[3]))))
      | (fsm_output[10]))));
  assign mux_2808_nl = MUX_s_1_2_2(or_tmp_14, nand_128_nl, fsm_output[7]);
  assign mux_2811_nl = MUX_s_1_2_2(mux_2810_nl, mux_2808_nl, fsm_output[5]);
  assign mux_2806_nl = MUX_s_1_2_2(or_tmp_2246, or_tmp_2474, fsm_output[7]);
  assign mux_2805_nl = MUX_s_1_2_2(mux_9_cse, nand_tmp_95, fsm_output[7]);
  assign mux_2807_nl = MUX_s_1_2_2(mux_2806_nl, mux_2805_nl, fsm_output[5]);
  assign mux_2812_nl = MUX_s_1_2_2(mux_2811_nl, mux_2807_nl, fsm_output[2]);
  assign mux_2821_nl = MUX_s_1_2_2(mux_2820_nl, mux_2812_nl, fsm_output[8]);
  assign nand_127_nl = ~((fsm_output[6]) & (~ mux_tmp_2800));
  assign or_2626_nl = (fsm_output[6]) | (~ (fsm_output[0])) | (fsm_output[1]) | (fsm_output[3])
      | (fsm_output[10]);
  assign mux_2801_nl = MUX_s_1_2_2(nand_127_nl, or_2626_nl, fsm_output[7]);
  assign or_2625_nl = (fsm_output[6]) | (~ nor_tmp_288);
  assign or_2624_nl = (fsm_output[6]) | (nand_237_cse & (fsm_output[3])) | (fsm_output[10]);
  assign mux_2798_nl = MUX_s_1_2_2(or_2625_nl, or_2624_nl, fsm_output[7]);
  assign mux_2802_nl = MUX_s_1_2_2(mux_2801_nl, mux_2798_nl, fsm_output[5]);
  assign or_2622_nl = (fsm_output[7]) | mux_tmp_2796;
  assign or_2620_nl = (fsm_output[0]) | (~ (fsm_output[1])) | (fsm_output[3]) | (fsm_output[10]);
  assign mux_2794_nl = MUX_s_1_2_2((fsm_output[10]), or_2620_nl, fsm_output[6]);
  assign mux_2795_nl = MUX_s_1_2_2(or_tmp_434, mux_2794_nl, fsm_output[7]);
  assign mux_2797_nl = MUX_s_1_2_2(or_2622_nl, mux_2795_nl, fsm_output[5]);
  assign mux_2803_nl = MUX_s_1_2_2(mux_2802_nl, mux_2797_nl, fsm_output[2]);
  assign mux_2791_nl = MUX_s_1_2_2(mux_9_cse, mux_tmp_2790, fsm_output[7]);
  assign nand_126_nl = ~((fsm_output[6]) & (~ or_tmp_2233));
  assign mux_2789_nl = MUX_s_1_2_2(mux_tmp_2788, nand_126_nl, fsm_output[7]);
  assign mux_2792_nl = MUX_s_1_2_2(mux_2791_nl, mux_2789_nl, fsm_output[5]);
  assign mux_2786_nl = MUX_s_1_2_2(or_tmp_2257, mux_7_cse, fsm_output[7]);
  assign mux_2787_nl = MUX_s_1_2_2(mux_2786_nl, mux_3_cse, fsm_output[5]);
  assign mux_2793_nl = MUX_s_1_2_2(mux_2792_nl, mux_2787_nl, fsm_output[2]);
  assign mux_2804_nl = MUX_s_1_2_2(mux_2803_nl, mux_2793_nl, fsm_output[8]);
  assign mux_2822_nl = MUX_s_1_2_2(mux_2821_nl, mux_2804_nl, fsm_output[4]);
  assign COMP_LOOP_COMP_LOOP_and_17_nl = (z_out_7[4:1]==4'b0011);
  assign nl_COMP_LOOP_1_acc_8_nl = tmp_10_lpi_4_dfm - modulo_result_mux_1_cse;
  assign COMP_LOOP_1_acc_8_nl = nl_COMP_LOOP_1_acc_8_nl[63:0];
  assign or_2838_nl = (fsm_output[3]) | (fsm_output[1]) | (~ (fsm_output[9])) | (~
      (fsm_output[4])) | (fsm_output[10]);
  assign mux_3178_nl = MUX_s_1_2_2(nand_tmp_148, or_2838_nl, fsm_output[0]);
  assign mux_3179_nl = MUX_s_1_2_2(or_2839_cse, mux_3178_nl, fsm_output[7]);
  assign nor_620_nl = ~((fsm_output[6:5]!=2'b00) | mux_3179_nl);
  assign nor_621_nl = ~((~ (fsm_output[5])) | (~ (fsm_output[7])) | (~ (fsm_output[0]))
      | (~ (fsm_output[3])) | (fsm_output[1]) | (fsm_output[9]) | nand_398_cse);
  assign nor_622_nl = ~((fsm_output[0]) | (fsm_output[3]) | (fsm_output[1]) | (~
      (fsm_output[9])) | (fsm_output[4]) | (fsm_output[10]));
  assign mux_3175_nl = MUX_s_1_2_2(and_464_cse, nor_622_nl, fsm_output[7]);
  assign nor_623_nl = ~((fsm_output[7]) | (fsm_output[0]) | (fsm_output[3]) | (~
      (fsm_output[1])) | (fsm_output[9]) | (fsm_output[4]) | (fsm_output[10]));
  assign mux_3176_nl = MUX_s_1_2_2(mux_3175_nl, nor_623_nl, fsm_output[5]);
  assign mux_3177_nl = MUX_s_1_2_2(nor_621_nl, mux_3176_nl, fsm_output[6]);
  assign mux_3180_nl = MUX_s_1_2_2(nor_620_nl, mux_3177_nl, fsm_output[8]);
  assign nor_624_nl = ~((fsm_output[7]) | (fsm_output[0]) | nand_226_cse);
  assign or_2828_nl = (fsm_output[1]) | (fsm_output[9]) | (~ (fsm_output[4])) | (fsm_output[10]);
  assign or_2827_nl = (fsm_output[1]) | (~ (fsm_output[9])) | (fsm_output[4]) | (fsm_output[10]);
  assign mux_3170_nl = MUX_s_1_2_2(or_2828_nl, or_2827_nl, fsm_output[3]);
  assign mux_3171_nl = MUX_s_1_2_2(mux_3170_nl, or_2826_cse, fsm_output[0]);
  assign nor_625_nl = ~((fsm_output[7]) | mux_3171_nl);
  assign mux_3172_nl = MUX_s_1_2_2(nor_624_nl, nor_625_nl, fsm_output[5]);
  assign mux_3169_nl = MUX_s_1_2_2(or_2824_cse, nand_tmp_148, fsm_output[0]);
  assign and_465_nl = (fsm_output[5]) & (fsm_output[7]) & (~ mux_3169_nl);
  assign mux_3173_nl = MUX_s_1_2_2(mux_3172_nl, and_465_nl, fsm_output[6]);
  assign or_2817_nl = (~ (fsm_output[0])) | (fsm_output[3]) | (~ (fsm_output[1]))
      | (fsm_output[9]) | (fsm_output[4]) | (fsm_output[10]);
  assign mux_3167_nl = MUX_s_1_2_2(or_2819_cse, or_2817_nl, fsm_output[7]);
  assign nor_626_nl = ~((fsm_output[6:5]!=2'b10) | mux_3167_nl);
  assign mux_3174_nl = MUX_s_1_2_2(mux_3173_nl, nor_626_nl, fsm_output[8]);
  assign mux_3181_nl = MUX_s_1_2_2(mux_3180_nl, mux_3174_nl, fsm_output[2]);
  assign COMP_LOOP_COMP_LOOP_and_10_nl = (VEC_LOOP_j_sva_11_0[3:0]==4'b1011);
  assign nl_COMP_LOOP_1_acc_nl = ({COMP_LOOP_k_9_4_sva_2 , 4'b0000}) + ({1'b1 , (~
      (STAGE_LOOP_lshift_psp_sva[9:1]))}) + 10'b0000000001;
  assign COMP_LOOP_1_acc_nl = nl_COMP_LOOP_1_acc_nl[9:0];
  assign nor_nl = ~((fsm_output[10]) | (fsm_output[8]) | (fsm_output[7]) | (fsm_output[6])
      | and_359_cse);
  assign mux_3215_nl = MUX_s_1_2_2(and_458_cse, and_459_cse, fsm_output[0]);
  assign or_3259_nl = (fsm_output[5]) | ((fsm_output[4]) & mux_3215_nl);
  assign nor_617_nl = ~((fsm_output[5:3]!=3'b000) | and_563_cse);
  assign mux_3216_nl = MUX_s_1_2_2(or_3259_nl, nor_617_nl, fsm_output[6]);
  assign or_2888_nl = (fsm_output[6:0]!=7'b0000000);
  assign mux_3217_nl = MUX_s_1_2_2(mux_3216_nl, or_2888_nl, fsm_output[7]);
  assign and_1253_nl = (fsm_output[10]) & ((fsm_output[8]) | mux_3217_nl);
  assign mux_3223_nl = MUX_s_1_2_2(mux_tmp_3219, nor_tmp_445, fsm_output[6]);
  assign mux_3220_nl = MUX_s_1_2_2(mux_tmp_3219, nor_tmp_445, or_2898_cse);
  assign and_452_nl = (and_517_cse | (fsm_output[8:7]!=2'b00)) & (fsm_output[9]);
  assign mux_3221_nl = MUX_s_1_2_2(mux_3220_nl, and_452_nl, fsm_output[1]);
  assign and_454_nl = (and_528_cse | (fsm_output[8:7]!=2'b00)) & (fsm_output[9]);
  assign mux_3222_nl = MUX_s_1_2_2(mux_3221_nl, and_454_nl, fsm_output[2]);
  assign mux_3224_nl = MUX_s_1_2_2(mux_3223_nl, mux_3222_nl, and_456_cse);
  assign mux_3231_nl = MUX_s_1_2_2((~ (fsm_output[6])), and_528_cse, fsm_output[7]);
  assign mux_3232_nl = MUX_s_1_2_2(and_dcpl_268, mux_3231_nl, fsm_output[5]);
  assign and_363_nl = (fsm_output[6]) & or_2902_cse;
  assign mux_3229_nl = MUX_s_1_2_2((~ (fsm_output[6])), and_363_nl, fsm_output[7]);
  assign mux_3230_nl = MUX_s_1_2_2(and_dcpl_268, mux_3229_nl, fsm_output[5]);
  assign mux_3233_nl = MUX_s_1_2_2(mux_3232_nl, mux_3230_nl, fsm_output[2]);
  assign nor_729_nl = ~((fsm_output[6]) | (fsm_output[1]) | (fsm_output[3]));
  assign mux_3226_nl = MUX_s_1_2_2(nor_729_nl, (fsm_output[6]), fsm_output[7]);
  assign mux_3227_nl = MUX_s_1_2_2(and_dcpl_268, mux_3226_nl, fsm_output[5]);
  assign mux_3225_nl = MUX_s_1_2_2(and_dcpl_268, and_450_cse, fsm_output[5]);
  assign mux_3228_nl = MUX_s_1_2_2(mux_3227_nl, mux_3225_nl, fsm_output[2]);
  assign mux_3234_nl = MUX_s_1_2_2(mux_3233_nl, mux_3228_nl, fsm_output[4]);
  assign nl_COMP_LOOP_acc_11_psp_sva  = (VEC_LOOP_j_sva_11_0[11:1]) + conv_u2u_8_11({COMP_LOOP_k_9_4_sva_4_0
      , 3'b001});
  assign mux_3239_nl = MUX_s_1_2_2((fsm_output[7]), or_2520_cse, fsm_output[5]);
  assign or_2906_nl = (fsm_output[7]) | and_528_cse;
  assign mux_3238_nl = MUX_s_1_2_2(or_2906_nl, or_2520_cse, fsm_output[5]);
  assign mux_3240_nl = MUX_s_1_2_2(mux_3239_nl, mux_3238_nl, fsm_output[2]);
  assign mux_3241_nl = MUX_s_1_2_2(and_dcpl_268, mux_3240_nl, fsm_output[8]);
  assign mux_3237_nl = MUX_s_1_2_2((~ mux_tmp_3236), or_2520_cse, fsm_output[8]);
  assign mux_3242_nl = MUX_s_1_2_2(mux_3241_nl, mux_3237_nl, fsm_output[4]);
  assign or_3252_nl = (fsm_output[8]) | and_359_cse | (fsm_output[6]);
  assign nand_218_nl = ~((fsm_output[8]) & ((((fsm_output[3:0]!=4'b0000)) & (fsm_output[5:4]==2'b11))
      | (fsm_output[6])));
  assign mux_3243_nl = MUX_s_1_2_2(or_3252_nl, nand_218_nl, fsm_output[7]);
  assign mux_3248_nl = MUX_s_1_2_2(mux_tmp_3244, or_tmp_2849, fsm_output[5]);
  assign mux_3245_nl = MUX_s_1_2_2(mux_tmp_3244, or_tmp_2849, and_563_cse);
  assign or_2915_nl = (~((fsm_output[1]) | (fsm_output[2]) | (fsm_output[6]) | (fsm_output[7])
      | (fsm_output[8]))) | (fsm_output[9]);
  assign mux_3246_nl = MUX_s_1_2_2(mux_3245_nl, or_2915_nl, fsm_output[5]);
  assign or_2913_nl = (~((fsm_output[8:5]!=4'b0000))) | (fsm_output[9]);
  assign mux_3247_nl = MUX_s_1_2_2(mux_3246_nl, or_2913_nl, fsm_output[3]);
  assign mux_3249_nl = MUX_s_1_2_2(mux_3248_nl, mux_3247_nl, fsm_output[4]);
  assign nl_COMP_LOOP_acc_14_psp_sva  = (VEC_LOOP_j_sva_11_0[11:1]) + conv_u2u_8_11({COMP_LOOP_k_9_4_sva_4_0
      , 3'b011});
  assign nor_1317_nl = ~((fsm_output[8]) | mux_tmp_3236);
  assign mux_3250_nl = MUX_s_1_2_2(nor_1316_cse, nor_1317_nl, fsm_output[4]);
  assign or_3346_nl = (fsm_output[8]) | ((fsm_output[7:5]==3'b111));
  assign mux_3251_nl = MUX_s_1_2_2(mux_3250_nl, or_3346_nl, fsm_output[9]);
  assign nl_COMP_LOOP_acc_1_cse_8_sva  = VEC_LOOP_j_sva_11_0 + conv_u2u_9_12({COMP_LOOP_k_9_4_sva_4_0
      , 4'b0111});
  assign nor_611_nl = ~((fsm_output[3]) | (fsm_output[2]) | (fsm_output[1]) | (fsm_output[8])
      | (fsm_output[9]));
  assign mux_3253_nl = MUX_s_1_2_2(nor_610_cse, nor_611_nl, and_456_cse);
  assign and_371_nl = (fsm_output[2]) & or_2348_cse & (fsm_output[9:8]==2'b11);
  assign or_2922_nl = (fsm_output[5:3]!=3'b000);
  assign mux_3252_nl = MUX_s_1_2_2(and_371_nl, nor_tmp_116, or_2922_nl);
  assign mux_3254_nl = MUX_s_1_2_2(mux_3253_nl, mux_3252_nl, fsm_output[6]);
  assign mux_3255_nl = MUX_s_1_2_2(mux_3254_nl, nor_tmp_116, fsm_output[7]);
  assign mux_3259_nl = MUX_s_1_2_2(mux_tmp_3256, nor_tmp_456, fsm_output[3]);
  assign mux_3260_nl = MUX_s_1_2_2(not_tmp_728, mux_3259_nl, fsm_output[4]);
  assign mux_3257_nl = MUX_s_1_2_2(not_tmp_728, mux_tmp_3256, fsm_output[3]);
  assign mux_3258_nl = MUX_s_1_2_2(mux_3257_nl, nor_tmp_456, fsm_output[4]);
  assign mux_3261_nl = MUX_s_1_2_2(mux_3260_nl, mux_3258_nl, or_2385_cse);
  assign mux_3262_nl = MUX_s_1_2_2(not_tmp_728, mux_3261_nl, fsm_output[5]);
  assign mux_3263_nl = MUX_s_1_2_2(mux_3262_nl, nor_tmp_456, fsm_output[6]);
  assign nl_COMP_LOOP_acc_1_cse_10_sva  = VEC_LOOP_j_sva_11_0 + conv_u2u_9_12({COMP_LOOP_k_9_4_sva_4_0
      , 4'b1001});
  assign or_2933_nl = (fsm_output[9:6]!=4'b0000);
  assign mux_3265_nl = MUX_s_1_2_2((~ (fsm_output[10])), (fsm_output[10]), or_2933_nl);
  assign mux_3266_nl = MUX_s_1_2_2(mux_3265_nl, or_tmp_2864, and_440_cse);
  assign mux_3267_nl = MUX_s_1_2_2(mux_3266_nl, or_tmp_2864, fsm_output[5]);
  assign or_2930_nl = (~((fsm_output[1]) | (fsm_output[2]) | (fsm_output[3]) | (fsm_output[6])
      | (fsm_output[7]) | (fsm_output[8]) | (fsm_output[9]))) | (fsm_output[10]);
  assign mux_3264_nl = MUX_s_1_2_2(or_tmp_2864, or_2930_nl, fsm_output[5]);
  assign nl_COMP_LOOP_acc_17_psp_sva  = (VEC_LOOP_j_sva_11_0[11:1]) + conv_u2u_8_11({COMP_LOOP_k_9_4_sva_4_0
      , 3'b101});
  assign mux_3275_nl = MUX_s_1_2_2(and_dcpl_264, (fsm_output[10]), or_2935_cse);
  assign mux_3271_nl = MUX_s_1_2_2(mux_tmp_2220, (fsm_output[10]), fsm_output[7]);
  assign mux_3272_nl = MUX_s_1_2_2(mux_tmp_3269, mux_3271_nl, fsm_output[5]);
  assign and_439_nl = or_2520_cse & (fsm_output[10]);
  assign mux_3270_nl = MUX_s_1_2_2(mux_tmp_3269, and_439_nl, fsm_output[5]);
  assign mux_3273_nl = MUX_s_1_2_2(mux_3272_nl, mux_3270_nl, fsm_output[2]);
  assign mux_3274_nl = MUX_s_1_2_2(mux_3273_nl, (fsm_output[10]), fsm_output[8]);
  assign mux_3276_nl = MUX_s_1_2_2(mux_3275_nl, mux_3274_nl, fsm_output[4]);
  assign nl_COMP_LOOP_acc_1_cse_12_sva  = VEC_LOOP_j_sva_11_0 + conv_u2u_9_12({COMP_LOOP_k_9_4_sva_4_0
      , 4'b1011});
  assign mux_3288_nl = MUX_s_1_2_2(mux_tmp_3281, mux_tmp_3280, fsm_output[5]);
  assign and_434_nl = (fsm_output[0]) & (fsm_output[3]);
  assign mux_3285_nl = MUX_s_1_2_2(mux_tmp_3281, mux_tmp_3280, and_434_nl);
  assign mux_3284_nl = MUX_s_1_2_2(mux_tmp_3280, nor_tmp_461, fsm_output[3]);
  assign mux_3286_nl = MUX_s_1_2_2(mux_3285_nl, mux_3284_nl, fsm_output[5]);
  assign mux_3282_nl = MUX_s_1_2_2(mux_tmp_3281, mux_tmp_3280, fsm_output[3]);
  assign mux_3283_nl = MUX_s_1_2_2(mux_3282_nl, nor_tmp_461, fsm_output[5]);
  assign mux_3287_nl = MUX_s_1_2_2(mux_3286_nl, mux_3283_nl, or_2385_cse);
  assign nor_604_nl = ~((fsm_output[8]) | (fsm_output[10]));
  assign nor_605_nl = ~((fsm_output[2]) | (fsm_output[3]) | (fsm_output[8]) | (fsm_output[10]));
  assign and_431_nl = (fsm_output[2]) & (fsm_output[3]) & (fsm_output[8]) & (fsm_output[10]);
  assign mux_3290_nl = MUX_s_1_2_2(nor_605_nl, and_431_nl, fsm_output[1]);
  assign mux_3291_nl = MUX_s_1_2_2(nor_604_nl, mux_3290_nl, and_456_cse);
  assign and_433_nl = (fsm_output[8]) & (fsm_output[10]);
  assign mux_3292_nl = MUX_s_1_2_2(mux_3291_nl, and_433_nl, or_2520_cse);
  assign nl_COMP_LOOP_acc_1_cse_14_sva  = VEC_LOOP_j_sva_11_0 + conv_u2u_9_12({COMP_LOOP_k_9_4_sva_4_0
      , 4'b1101});
  assign or_2947_nl = (fsm_output[2]) | (fsm_output[3]) | (fsm_output[1]) | (fsm_output[10]);
  assign mux_3296_nl = MUX_s_1_2_2((fsm_output[10]), or_2947_nl, and_456_cse);
  assign nor_603_nl = ~((fsm_output[8]) | (fsm_output[6]) | mux_3296_nl);
  assign and_430_nl = (fsm_output[0]) & (fsm_output[1]) & (fsm_output[10]);
  assign or_2945_nl = (fsm_output[4:2]!=3'b000);
  assign mux_3294_nl = MUX_s_1_2_2(and_430_nl, (fsm_output[10]), or_2945_nl);
  assign and_374_nl = (fsm_output[5]) & mux_3294_nl;
  assign mux_3295_nl = MUX_s_1_2_2(and_374_nl, (fsm_output[10]), fsm_output[6]);
  assign and_375_nl = (fsm_output[8]) & mux_3295_nl;
  assign mux_3297_nl = MUX_s_1_2_2(nor_603_nl, and_375_nl, fsm_output[7]);
  assign nl_COMP_LOOP_acc_20_psp_sva  = (VEC_LOOP_j_sva_11_0[11:1]) + conv_u2u_8_11({COMP_LOOP_k_9_4_sva_4_0
      , 3'b111});
  assign or_2950_nl = (fsm_output[1]) | (fsm_output[2]) | (fsm_output[3]) | (fsm_output[6])
      | (fsm_output[7]) | (fsm_output[8]);
  assign mux_3299_nl = MUX_s_1_2_2(or_2951_cse, or_2950_nl, and_456_cse);
  assign nor_1420_nl = ~((fsm_output[10]) | mux_3299_nl);
  assign and_1254_nl = (fsm_output[10]) & ((fsm_output[8:3]!=6'b000000));
  assign nl_COMP_LOOP_acc_1_cse_sva  = VEC_LOOP_j_sva_11_0 + conv_u2u_9_12({COMP_LOOP_k_9_4_sva_4_0
      , 4'b1111});
  assign nor_1201_nl = ~((fsm_output[6]) | (fsm_output[9]) | (fsm_output[10]));
  assign mux_3302_nl = MUX_s_1_2_2(nor_601_cse, nor_1203_cse, fsm_output[4]);
  assign and_29_nl = (fsm_output[2]) & or_2348_cse & (fsm_output[3]) & (fsm_output[9])
      & (fsm_output[10]);
  assign mux_3301_nl = MUX_s_1_2_2(and_29_nl, and_816_cse, fsm_output[4]);
  assign mux_3303_nl = MUX_s_1_2_2(mux_3302_nl, mux_3301_nl, fsm_output[6]);
  assign mux_3304_nl = MUX_s_1_2_2(nor_1201_nl, mux_3303_nl, fsm_output[5]);
  assign COMP_LOOP_COMP_LOOP_or_15_nl = (VEC_LOOP_j_sva_11_0[11]) | and_850_cse |
      and_857_cse | and_dcpl_378 | and_869_cse | and_875_cse | and_dcpl_394 | and_886_cse
      | and_dcpl_404 | and_dcpl_408 | and_dcpl_411 | and_dcpl_415;
  assign COMP_LOOP_COMP_LOOP_mux_18_nl = MUX_v_9_2_2((VEC_LOOP_j_sva_11_0[10:2]),
      (~ (STAGE_LOOP_lshift_psp_sva[9:1])), COMP_LOOP_or_60_itm);
  assign COMP_LOOP_or_77_nl = (~ and_dcpl_356) | and_850_cse | and_857_cse | and_dcpl_378
      | and_869_cse | and_875_cse | and_dcpl_394 | and_886_cse | and_dcpl_404 | and_dcpl_408
      | and_dcpl_411 | and_dcpl_415;
  assign COMP_LOOP_COMP_LOOP_mux_19_nl = MUX_v_5_2_2(({2'b00 , (COMP_LOOP_k_9_4_sva_4_0[4:2])}),
      COMP_LOOP_k_9_4_sva_4_0, COMP_LOOP_or_60_itm);
  assign COMP_LOOP_COMP_LOOP_or_16_nl = ((COMP_LOOP_k_9_4_sva_4_0[1]) & (~(and_850_cse
      | and_857_cse | and_dcpl_378 | and_869_cse | and_875_cse))) | and_dcpl_394
      | and_886_cse | and_dcpl_404 | and_dcpl_408 | and_dcpl_411 | and_dcpl_415;
  assign COMP_LOOP_COMP_LOOP_or_17_nl = ((COMP_LOOP_k_9_4_sva_4_0[0]) & (~(and_850_cse
      | and_857_cse | and_dcpl_394 | and_886_cse | and_dcpl_404))) | and_dcpl_378
      | and_869_cse | and_875_cse | and_dcpl_408 | and_dcpl_411 | and_dcpl_415;
  assign COMP_LOOP_COMP_LOOP_or_18_nl = (~(and_dcpl_356 | and_850_cse | and_dcpl_378
      | and_869_cse | and_dcpl_394 | and_886_cse | and_dcpl_408 | and_dcpl_411))
      | and_857_cse | and_875_cse | and_dcpl_404 | and_dcpl_415;
  assign COMP_LOOP_COMP_LOOP_or_19_nl = (~(and_857_cse | and_dcpl_378 | and_875_cse
      | and_dcpl_394 | and_dcpl_404 | and_dcpl_408 | and_dcpl_415)) | and_dcpl_356
      | and_850_cse | and_869_cse | and_886_cse | and_dcpl_411;
  assign nl_acc_nl = ({COMP_LOOP_COMP_LOOP_or_15_nl , COMP_LOOP_COMP_LOOP_mux_18_nl
      , COMP_LOOP_or_77_nl}) + conv_u2u_10_11({COMP_LOOP_COMP_LOOP_mux_19_nl , COMP_LOOP_COMP_LOOP_or_16_nl
      , COMP_LOOP_COMP_LOOP_or_17_nl , COMP_LOOP_COMP_LOOP_or_18_nl , COMP_LOOP_COMP_LOOP_or_19_nl
      , 1'b1});
  assign acc_nl = nl_acc_nl[10:0];
  assign z_out = readslicef_11_10_1(acc_nl);
  assign COMP_LOOP_mux_84_nl = MUX_v_10_2_2((VEC_LOOP_j_sva_11_0[11:2]), STAGE_LOOP_lshift_psp_sva,
      COMP_LOOP_or_24_itm);
  assign COMP_LOOP_COMP_LOOP_mux_20_nl = MUX_v_5_2_2(({2'b00 , (COMP_LOOP_k_9_4_sva_4_0[4:2])}),
      COMP_LOOP_k_9_4_sva_4_0, COMP_LOOP_or_24_itm);
  assign COMP_LOOP_mux_85_nl = MUX_v_2_2_2((COMP_LOOP_k_9_4_sva_4_0[1:0]), 2'b01,
      and_dcpl_433);
  assign COMP_LOOP_COMP_LOOP_or_20_nl = MUX_v_2_2_2(COMP_LOOP_mux_85_nl, 2'b11, and_dcpl_441);
  assign nl_z_out_1 = COMP_LOOP_mux_84_nl + conv_u2u_9_10({COMP_LOOP_COMP_LOOP_mux_20_nl
      , COMP_LOOP_COMP_LOOP_or_20_nl , COMP_LOOP_COMP_LOOP_or_6_cse , COMP_LOOP_COMP_LOOP_or_6_cse});
  assign z_out_1 = nl_z_out_1[9:0];
  assign and_1278_nl = and_dcpl_353 & (~ (fsm_output[9])) & (~ (fsm_output[8])) &
      (fsm_output[7]) & (fsm_output[5]) & (fsm_output[3]) & (fsm_output[2]) & (fsm_output[1])
      & and_dcpl_107;
  assign and_1279_nl = (~ (fsm_output[4])) & (~ (fsm_output[10])) & (~ (fsm_output[9]))
      & and_dcpl_373 & (~ (fsm_output[5])) & (fsm_output[3]) & (~ (fsm_output[2]))
      & (~ (fsm_output[1])) & and_dcpl_107;
  assign and_1280_nl = (~ (fsm_output[4])) & (fsm_output[10]) & (~ (fsm_output[9]))
      & and_dcpl_373 & (fsm_output[5]) & and_dcpl_348 & (~ (fsm_output[1])) & (fsm_output[6])
      & (~ (fsm_output[0]));
  assign COMP_LOOP_mux1h_585_nl = MUX1HOT_v_4_4_2(4'b0001, 4'b0011, 4'b0101, 4'b1110,
      {and_1278_nl , and_1279_nl , (fsm_output[9]) , and_1280_nl});
  assign nl_z_out_2 = STAGE_LOOP_lshift_psp_sva + conv_u2u_9_10({COMP_LOOP_k_9_4_sva_4_0
      , COMP_LOOP_mux1h_585_nl});
  assign z_out_2 = nl_z_out_2[9:0];
  assign and_1281_nl = and_dcpl_503 & (~ (fsm_output[9])) & and_dcpl_502 & (fsm_output[3])
      & (fsm_output[2]) & (~ (fsm_output[1])) & (fsm_output[6]) & (~ (fsm_output[0]));
  assign COMP_LOOP_mux_86_nl = MUX_v_2_2_2(2'b10, 2'b01, and_1281_nl);
  assign and_1282_nl = (~ (fsm_output[10])) & (~ (fsm_output[4])) & (~ (fsm_output[9]))
      & (fsm_output[8]) & (~ (fsm_output[7])) & (fsm_output[5]) & and_dcpl_480 &
      and_dcpl_99;
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_53_nl = ~(MUX_v_2_2_2(COMP_LOOP_mux_86_nl,
      2'b11, and_1282_nl));
  assign COMP_LOOP_or_78_nl = MUX_v_2_2_2(COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_53_nl,
      2'b11, and_dcpl_511);
  assign nl_z_out_3 = STAGE_LOOP_lshift_psp_sva + conv_u2u_9_10({COMP_LOOP_k_9_4_sva_4_0
      , COMP_LOOP_or_78_nl , 1'b1 , and_dcpl_511});
  assign z_out_3 = nl_z_out_3[9:0];
  assign and_1283_nl = and_dcpl_375 & (~ (fsm_output[9])) & and_dcpl_517 & (fsm_output[3])
      & (fsm_output[2]) & (fsm_output[1]) & (fsm_output[6]) & (~ (fsm_output[0]));
  assign and_1284_nl = and_dcpl_375 & (fsm_output[9]) & and_dcpl_517 & (fsm_output[3:1]==3'b011)
      & nor_tmp_217;
  assign and_1285_nl = and_dcpl_406 & (fsm_output[8]) & (~ (fsm_output[7])) & (fsm_output[5])
      & (fsm_output[3]) & (~ (fsm_output[2])) & (fsm_output[1]) & nor_tmp_217;
  assign COMP_LOOP_mux1h_586_nl = MUX1HOT_v_4_4_2(4'b0100, 4'b1001, 4'b1011, 4'b1101,
      {and_1283_nl , and_1284_nl , (~ (fsm_output[1])) , and_1285_nl});
  assign nl_z_out_4 = STAGE_LOOP_lshift_psp_sva + conv_u2u_9_10({COMP_LOOP_k_9_4_sva_4_0
      , COMP_LOOP_mux1h_586_nl});
  assign z_out_4 = nl_z_out_4[9:0];
  assign COMP_LOOP_mux1h_587_nl = MUX1HOT_v_64_3_2(({52'b0000000000000000000000000000000000000000000000000000
      , VEC_LOOP_j_sva_11_0}), tmp_10_lpi_4_dfm, ({1'b1 , (~ (operator_64_false_acc_mut_63_0[62:0]))}),
      {and_dcpl_555 , (~ mux_3724_itm) , and_dcpl_564});
  assign COMP_LOOP_mux1h_588_nl = MUX1HOT_v_64_3_2(({55'b0000000000000000000000000000000000000000000000000000000
      , COMP_LOOP_k_9_4_sva_4_0 , 4'b0011}), modulo_result_mux_1_cse, 64'b0000000000000000000000000000000000000000000000000000000000000001,
      {and_dcpl_555 , (~ mux_3724_itm) , and_dcpl_564});
  assign nl_z_out_5 = COMP_LOOP_mux1h_587_nl + COMP_LOOP_mux1h_588_nl;
  assign z_out_5 = nl_z_out_5[63:0];
  assign operator_64_false_1_mux1h_2_nl = MUX1HOT_v_64_4_2(({59'b00000000000000000000000000000000000000000000000000000000001
      , (~ COMP_LOOP_k_9_4_sva_4_0)}), modulo_result_rem_cmp_z, p_sva, ({52'b0000000000000000000000000000000000000000000000000000
      , VEC_LOOP_j_sva_11_0}), {and_dcpl_574 , (~ mux_3788_itm) , and_dcpl_579 ,
      and_dcpl_588});
  assign operator_64_false_1_mux1h_3_nl = MUX1HOT_v_64_3_2(64'b0000000000000000000000000000000000000000000000000000000000000001,
      p_sva, ({54'b000000000000000000000000000000000000000000000000000000 , STAGE_LOOP_lshift_psp_sva}),
      {and_dcpl_574 , (~ mux_3788_itm) , and_dcpl_588});
  assign operator_64_false_1_or_1_nl = MUX_v_64_2_2(operator_64_false_1_mux1h_3_nl,
      64'b1111111111111111111111111111111111111111111111111111111111111111, and_dcpl_579);
  assign nl_z_out_6 = conv_u2u_64_65(operator_64_false_1_mux1h_2_nl) + conv_s2u_64_65(operator_64_false_1_or_1_nl);
  assign z_out_6 = nl_z_out_6[64:0];
  assign COMP_LOOP_COMP_LOOP_or_21_nl = (~(and_dcpl_598 | and_850_cse | and_857_cse
      | and_dcpl_622 | and_dcpl_628 | and_869_cse | and_875_cse | and_dcpl_641 |
      and_dcpl_646 | and_886_cse | and_dcpl_654 | and_dcpl_659 | and_dcpl_663 | and_dcpl_666
      | and_dcpl_669 | and_dcpl_672 | and_dcpl_676)) | and_dcpl_678;
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_54_nl = ~((operator_66_true_div_cmp_z[63])
      | and_dcpl_598 | and_850_cse | and_857_cse | and_dcpl_622 | and_dcpl_628 |
      and_869_cse | and_875_cse | and_dcpl_641 | and_dcpl_646 | and_886_cse | and_dcpl_654
      | and_dcpl_659 | and_dcpl_663 | and_dcpl_666 | and_dcpl_669 | and_dcpl_672
      | and_dcpl_676);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_55_nl = ~((operator_66_true_div_cmp_z[62])
      | and_dcpl_598 | and_850_cse | and_857_cse | and_dcpl_622 | and_dcpl_628 |
      and_869_cse | and_875_cse | and_dcpl_641 | and_dcpl_646 | and_886_cse | and_dcpl_654
      | and_dcpl_659 | and_dcpl_663 | and_dcpl_666 | and_dcpl_669 | and_dcpl_672
      | and_dcpl_676);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_56_nl = ~((operator_66_true_div_cmp_z[61])
      | and_dcpl_598 | and_850_cse | and_857_cse | and_dcpl_622 | and_dcpl_628 |
      and_869_cse | and_875_cse | and_dcpl_641 | and_dcpl_646 | and_886_cse | and_dcpl_654
      | and_dcpl_659 | and_dcpl_663 | and_dcpl_666 | and_dcpl_669 | and_dcpl_672
      | and_dcpl_676);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_57_nl = ~((operator_66_true_div_cmp_z[60])
      | and_dcpl_598 | and_850_cse | and_857_cse | and_dcpl_622 | and_dcpl_628 |
      and_869_cse | and_875_cse | and_dcpl_641 | and_dcpl_646 | and_886_cse | and_dcpl_654
      | and_dcpl_659 | and_dcpl_663 | and_dcpl_666 | and_dcpl_669 | and_dcpl_672
      | and_dcpl_676);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_58_nl = ~((operator_66_true_div_cmp_z[59])
      | and_dcpl_598 | and_850_cse | and_857_cse | and_dcpl_622 | and_dcpl_628 |
      and_869_cse | and_875_cse | and_dcpl_641 | and_dcpl_646 | and_886_cse | and_dcpl_654
      | and_dcpl_659 | and_dcpl_663 | and_dcpl_666 | and_dcpl_669 | and_dcpl_672
      | and_dcpl_676);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_59_nl = ~((operator_66_true_div_cmp_z[58])
      | and_dcpl_598 | and_850_cse | and_857_cse | and_dcpl_622 | and_dcpl_628 |
      and_869_cse | and_875_cse | and_dcpl_641 | and_dcpl_646 | and_886_cse | and_dcpl_654
      | and_dcpl_659 | and_dcpl_663 | and_dcpl_666 | and_dcpl_669 | and_dcpl_672
      | and_dcpl_676);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_60_nl = ~((operator_66_true_div_cmp_z[57])
      | and_dcpl_598 | and_850_cse | and_857_cse | and_dcpl_622 | and_dcpl_628 |
      and_869_cse | and_875_cse | and_dcpl_641 | and_dcpl_646 | and_886_cse | and_dcpl_654
      | and_dcpl_659 | and_dcpl_663 | and_dcpl_666 | and_dcpl_669 | and_dcpl_672
      | and_dcpl_676);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_61_nl = ~((operator_66_true_div_cmp_z[56])
      | and_dcpl_598 | and_850_cse | and_857_cse | and_dcpl_622 | and_dcpl_628 |
      and_869_cse | and_875_cse | and_dcpl_641 | and_dcpl_646 | and_886_cse | and_dcpl_654
      | and_dcpl_659 | and_dcpl_663 | and_dcpl_666 | and_dcpl_669 | and_dcpl_672
      | and_dcpl_676);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_62_nl = ~((operator_66_true_div_cmp_z[55])
      | and_dcpl_598 | and_850_cse | and_857_cse | and_dcpl_622 | and_dcpl_628 |
      and_869_cse | and_875_cse | and_dcpl_641 | and_dcpl_646 | and_886_cse | and_dcpl_654
      | and_dcpl_659 | and_dcpl_663 | and_dcpl_666 | and_dcpl_669 | and_dcpl_672
      | and_dcpl_676);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_63_nl = ~((operator_66_true_div_cmp_z[54])
      | and_dcpl_598 | and_850_cse | and_857_cse | and_dcpl_622 | and_dcpl_628 |
      and_869_cse | and_875_cse | and_dcpl_641 | and_dcpl_646 | and_886_cse | and_dcpl_654
      | and_dcpl_659 | and_dcpl_663 | and_dcpl_666 | and_dcpl_669 | and_dcpl_672
      | and_dcpl_676);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_64_nl = ~((operator_66_true_div_cmp_z[53])
      | and_dcpl_598 | and_850_cse | and_857_cse | and_dcpl_622 | and_dcpl_628 |
      and_869_cse | and_875_cse | and_dcpl_641 | and_dcpl_646 | and_886_cse | and_dcpl_654
      | and_dcpl_659 | and_dcpl_663 | and_dcpl_666 | and_dcpl_669 | and_dcpl_672
      | and_dcpl_676);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_65_nl = ~((operator_66_true_div_cmp_z[52])
      | and_dcpl_598 | and_850_cse | and_857_cse | and_dcpl_622 | and_dcpl_628 |
      and_869_cse | and_875_cse | and_dcpl_641 | and_dcpl_646 | and_886_cse | and_dcpl_654
      | and_dcpl_659 | and_dcpl_663 | and_dcpl_666 | and_dcpl_669 | and_dcpl_672
      | and_dcpl_676);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_66_nl = ~((operator_66_true_div_cmp_z[51])
      | and_dcpl_598 | and_850_cse | and_857_cse | and_dcpl_622 | and_dcpl_628 |
      and_869_cse | and_875_cse | and_dcpl_641 | and_dcpl_646 | and_886_cse | and_dcpl_654
      | and_dcpl_659 | and_dcpl_663 | and_dcpl_666 | and_dcpl_669 | and_dcpl_672
      | and_dcpl_676);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_67_nl = ~((operator_66_true_div_cmp_z[50])
      | and_dcpl_598 | and_850_cse | and_857_cse | and_dcpl_622 | and_dcpl_628 |
      and_869_cse | and_875_cse | and_dcpl_641 | and_dcpl_646 | and_886_cse | and_dcpl_654
      | and_dcpl_659 | and_dcpl_663 | and_dcpl_666 | and_dcpl_669 | and_dcpl_672
      | and_dcpl_676);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_68_nl = ~((operator_66_true_div_cmp_z[49])
      | and_dcpl_598 | and_850_cse | and_857_cse | and_dcpl_622 | and_dcpl_628 |
      and_869_cse | and_875_cse | and_dcpl_641 | and_dcpl_646 | and_886_cse | and_dcpl_654
      | and_dcpl_659 | and_dcpl_663 | and_dcpl_666 | and_dcpl_669 | and_dcpl_672
      | and_dcpl_676);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_69_nl = ~((operator_66_true_div_cmp_z[48])
      | and_dcpl_598 | and_850_cse | and_857_cse | and_dcpl_622 | and_dcpl_628 |
      and_869_cse | and_875_cse | and_dcpl_641 | and_dcpl_646 | and_886_cse | and_dcpl_654
      | and_dcpl_659 | and_dcpl_663 | and_dcpl_666 | and_dcpl_669 | and_dcpl_672
      | and_dcpl_676);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_70_nl = ~((operator_66_true_div_cmp_z[47])
      | and_dcpl_598 | and_850_cse | and_857_cse | and_dcpl_622 | and_dcpl_628 |
      and_869_cse | and_875_cse | and_dcpl_641 | and_dcpl_646 | and_886_cse | and_dcpl_654
      | and_dcpl_659 | and_dcpl_663 | and_dcpl_666 | and_dcpl_669 | and_dcpl_672
      | and_dcpl_676);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_71_nl = ~((operator_66_true_div_cmp_z[46])
      | and_dcpl_598 | and_850_cse | and_857_cse | and_dcpl_622 | and_dcpl_628 |
      and_869_cse | and_875_cse | and_dcpl_641 | and_dcpl_646 | and_886_cse | and_dcpl_654
      | and_dcpl_659 | and_dcpl_663 | and_dcpl_666 | and_dcpl_669 | and_dcpl_672
      | and_dcpl_676);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_72_nl = ~((operator_66_true_div_cmp_z[45])
      | and_dcpl_598 | and_850_cse | and_857_cse | and_dcpl_622 | and_dcpl_628 |
      and_869_cse | and_875_cse | and_dcpl_641 | and_dcpl_646 | and_886_cse | and_dcpl_654
      | and_dcpl_659 | and_dcpl_663 | and_dcpl_666 | and_dcpl_669 | and_dcpl_672
      | and_dcpl_676);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_73_nl = ~((operator_66_true_div_cmp_z[44])
      | and_dcpl_598 | and_850_cse | and_857_cse | and_dcpl_622 | and_dcpl_628 |
      and_869_cse | and_875_cse | and_dcpl_641 | and_dcpl_646 | and_886_cse | and_dcpl_654
      | and_dcpl_659 | and_dcpl_663 | and_dcpl_666 | and_dcpl_669 | and_dcpl_672
      | and_dcpl_676);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_74_nl = ~((operator_66_true_div_cmp_z[43])
      | and_dcpl_598 | and_850_cse | and_857_cse | and_dcpl_622 | and_dcpl_628 |
      and_869_cse | and_875_cse | and_dcpl_641 | and_dcpl_646 | and_886_cse | and_dcpl_654
      | and_dcpl_659 | and_dcpl_663 | and_dcpl_666 | and_dcpl_669 | and_dcpl_672
      | and_dcpl_676);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_75_nl = ~((operator_66_true_div_cmp_z[42])
      | and_dcpl_598 | and_850_cse | and_857_cse | and_dcpl_622 | and_dcpl_628 |
      and_869_cse | and_875_cse | and_dcpl_641 | and_dcpl_646 | and_886_cse | and_dcpl_654
      | and_dcpl_659 | and_dcpl_663 | and_dcpl_666 | and_dcpl_669 | and_dcpl_672
      | and_dcpl_676);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_76_nl = ~((operator_66_true_div_cmp_z[41])
      | and_dcpl_598 | and_850_cse | and_857_cse | and_dcpl_622 | and_dcpl_628 |
      and_869_cse | and_875_cse | and_dcpl_641 | and_dcpl_646 | and_886_cse | and_dcpl_654
      | and_dcpl_659 | and_dcpl_663 | and_dcpl_666 | and_dcpl_669 | and_dcpl_672
      | and_dcpl_676);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_77_nl = ~((operator_66_true_div_cmp_z[40])
      | and_dcpl_598 | and_850_cse | and_857_cse | and_dcpl_622 | and_dcpl_628 |
      and_869_cse | and_875_cse | and_dcpl_641 | and_dcpl_646 | and_886_cse | and_dcpl_654
      | and_dcpl_659 | and_dcpl_663 | and_dcpl_666 | and_dcpl_669 | and_dcpl_672
      | and_dcpl_676);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_78_nl = ~((operator_66_true_div_cmp_z[39])
      | and_dcpl_598 | and_850_cse | and_857_cse | and_dcpl_622 | and_dcpl_628 |
      and_869_cse | and_875_cse | and_dcpl_641 | and_dcpl_646 | and_886_cse | and_dcpl_654
      | and_dcpl_659 | and_dcpl_663 | and_dcpl_666 | and_dcpl_669 | and_dcpl_672
      | and_dcpl_676);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_79_nl = ~((operator_66_true_div_cmp_z[38])
      | and_dcpl_598 | and_850_cse | and_857_cse | and_dcpl_622 | and_dcpl_628 |
      and_869_cse | and_875_cse | and_dcpl_641 | and_dcpl_646 | and_886_cse | and_dcpl_654
      | and_dcpl_659 | and_dcpl_663 | and_dcpl_666 | and_dcpl_669 | and_dcpl_672
      | and_dcpl_676);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_80_nl = ~((operator_66_true_div_cmp_z[37])
      | and_dcpl_598 | and_850_cse | and_857_cse | and_dcpl_622 | and_dcpl_628 |
      and_869_cse | and_875_cse | and_dcpl_641 | and_dcpl_646 | and_886_cse | and_dcpl_654
      | and_dcpl_659 | and_dcpl_663 | and_dcpl_666 | and_dcpl_669 | and_dcpl_672
      | and_dcpl_676);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_81_nl = ~((operator_66_true_div_cmp_z[36])
      | and_dcpl_598 | and_850_cse | and_857_cse | and_dcpl_622 | and_dcpl_628 |
      and_869_cse | and_875_cse | and_dcpl_641 | and_dcpl_646 | and_886_cse | and_dcpl_654
      | and_dcpl_659 | and_dcpl_663 | and_dcpl_666 | and_dcpl_669 | and_dcpl_672
      | and_dcpl_676);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_82_nl = ~((operator_66_true_div_cmp_z[35])
      | and_dcpl_598 | and_850_cse | and_857_cse | and_dcpl_622 | and_dcpl_628 |
      and_869_cse | and_875_cse | and_dcpl_641 | and_dcpl_646 | and_886_cse | and_dcpl_654
      | and_dcpl_659 | and_dcpl_663 | and_dcpl_666 | and_dcpl_669 | and_dcpl_672
      | and_dcpl_676);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_83_nl = ~((operator_66_true_div_cmp_z[34])
      | and_dcpl_598 | and_850_cse | and_857_cse | and_dcpl_622 | and_dcpl_628 |
      and_869_cse | and_875_cse | and_dcpl_641 | and_dcpl_646 | and_886_cse | and_dcpl_654
      | and_dcpl_659 | and_dcpl_663 | and_dcpl_666 | and_dcpl_669 | and_dcpl_672
      | and_dcpl_676);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_84_nl = ~((operator_66_true_div_cmp_z[33])
      | and_dcpl_598 | and_850_cse | and_857_cse | and_dcpl_622 | and_dcpl_628 |
      and_869_cse | and_875_cse | and_dcpl_641 | and_dcpl_646 | and_886_cse | and_dcpl_654
      | and_dcpl_659 | and_dcpl_663 | and_dcpl_666 | and_dcpl_669 | and_dcpl_672
      | and_dcpl_676);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_85_nl = ~((operator_66_true_div_cmp_z[32])
      | and_dcpl_598 | and_850_cse | and_857_cse | and_dcpl_622 | and_dcpl_628 |
      and_869_cse | and_875_cse | and_dcpl_641 | and_dcpl_646 | and_886_cse | and_dcpl_654
      | and_dcpl_659 | and_dcpl_663 | and_dcpl_666 | and_dcpl_669 | and_dcpl_672
      | and_dcpl_676);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_86_nl = ~((operator_66_true_div_cmp_z[31])
      | and_dcpl_598 | and_850_cse | and_857_cse | and_dcpl_622 | and_dcpl_628 |
      and_869_cse | and_875_cse | and_dcpl_641 | and_dcpl_646 | and_886_cse | and_dcpl_654
      | and_dcpl_659 | and_dcpl_663 | and_dcpl_666 | and_dcpl_669 | and_dcpl_672
      | and_dcpl_676);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_87_nl = ~((operator_66_true_div_cmp_z[30])
      | and_dcpl_598 | and_850_cse | and_857_cse | and_dcpl_622 | and_dcpl_628 |
      and_869_cse | and_875_cse | and_dcpl_641 | and_dcpl_646 | and_886_cse | and_dcpl_654
      | and_dcpl_659 | and_dcpl_663 | and_dcpl_666 | and_dcpl_669 | and_dcpl_672
      | and_dcpl_676);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_88_nl = ~((operator_66_true_div_cmp_z[29])
      | and_dcpl_598 | and_850_cse | and_857_cse | and_dcpl_622 | and_dcpl_628 |
      and_869_cse | and_875_cse | and_dcpl_641 | and_dcpl_646 | and_886_cse | and_dcpl_654
      | and_dcpl_659 | and_dcpl_663 | and_dcpl_666 | and_dcpl_669 | and_dcpl_672
      | and_dcpl_676);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_89_nl = ~((operator_66_true_div_cmp_z[28])
      | and_dcpl_598 | and_850_cse | and_857_cse | and_dcpl_622 | and_dcpl_628 |
      and_869_cse | and_875_cse | and_dcpl_641 | and_dcpl_646 | and_886_cse | and_dcpl_654
      | and_dcpl_659 | and_dcpl_663 | and_dcpl_666 | and_dcpl_669 | and_dcpl_672
      | and_dcpl_676);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_90_nl = ~((operator_66_true_div_cmp_z[27])
      | and_dcpl_598 | and_850_cse | and_857_cse | and_dcpl_622 | and_dcpl_628 |
      and_869_cse | and_875_cse | and_dcpl_641 | and_dcpl_646 | and_886_cse | and_dcpl_654
      | and_dcpl_659 | and_dcpl_663 | and_dcpl_666 | and_dcpl_669 | and_dcpl_672
      | and_dcpl_676);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_91_nl = ~((operator_66_true_div_cmp_z[26])
      | and_dcpl_598 | and_850_cse | and_857_cse | and_dcpl_622 | and_dcpl_628 |
      and_869_cse | and_875_cse | and_dcpl_641 | and_dcpl_646 | and_886_cse | and_dcpl_654
      | and_dcpl_659 | and_dcpl_663 | and_dcpl_666 | and_dcpl_669 | and_dcpl_672
      | and_dcpl_676);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_92_nl = ~((operator_66_true_div_cmp_z[25])
      | and_dcpl_598 | and_850_cse | and_857_cse | and_dcpl_622 | and_dcpl_628 |
      and_869_cse | and_875_cse | and_dcpl_641 | and_dcpl_646 | and_886_cse | and_dcpl_654
      | and_dcpl_659 | and_dcpl_663 | and_dcpl_666 | and_dcpl_669 | and_dcpl_672
      | and_dcpl_676);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_93_nl = ~((operator_66_true_div_cmp_z[24])
      | and_dcpl_598 | and_850_cse | and_857_cse | and_dcpl_622 | and_dcpl_628 |
      and_869_cse | and_875_cse | and_dcpl_641 | and_dcpl_646 | and_886_cse | and_dcpl_654
      | and_dcpl_659 | and_dcpl_663 | and_dcpl_666 | and_dcpl_669 | and_dcpl_672
      | and_dcpl_676);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_94_nl = ~((operator_66_true_div_cmp_z[23])
      | and_dcpl_598 | and_850_cse | and_857_cse | and_dcpl_622 | and_dcpl_628 |
      and_869_cse | and_875_cse | and_dcpl_641 | and_dcpl_646 | and_886_cse | and_dcpl_654
      | and_dcpl_659 | and_dcpl_663 | and_dcpl_666 | and_dcpl_669 | and_dcpl_672
      | and_dcpl_676);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_95_nl = ~((operator_66_true_div_cmp_z[22])
      | and_dcpl_598 | and_850_cse | and_857_cse | and_dcpl_622 | and_dcpl_628 |
      and_869_cse | and_875_cse | and_dcpl_641 | and_dcpl_646 | and_886_cse | and_dcpl_654
      | and_dcpl_659 | and_dcpl_663 | and_dcpl_666 | and_dcpl_669 | and_dcpl_672
      | and_dcpl_676);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_96_nl = ~((operator_66_true_div_cmp_z[21])
      | and_dcpl_598 | and_850_cse | and_857_cse | and_dcpl_622 | and_dcpl_628 |
      and_869_cse | and_875_cse | and_dcpl_641 | and_dcpl_646 | and_886_cse | and_dcpl_654
      | and_dcpl_659 | and_dcpl_663 | and_dcpl_666 | and_dcpl_669 | and_dcpl_672
      | and_dcpl_676);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_97_nl = ~((operator_66_true_div_cmp_z[20])
      | and_dcpl_598 | and_850_cse | and_857_cse | and_dcpl_622 | and_dcpl_628 |
      and_869_cse | and_875_cse | and_dcpl_641 | and_dcpl_646 | and_886_cse | and_dcpl_654
      | and_dcpl_659 | and_dcpl_663 | and_dcpl_666 | and_dcpl_669 | and_dcpl_672
      | and_dcpl_676);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_98_nl = ~((operator_66_true_div_cmp_z[19])
      | and_dcpl_598 | and_850_cse | and_857_cse | and_dcpl_622 | and_dcpl_628 |
      and_869_cse | and_875_cse | and_dcpl_641 | and_dcpl_646 | and_886_cse | and_dcpl_654
      | and_dcpl_659 | and_dcpl_663 | and_dcpl_666 | and_dcpl_669 | and_dcpl_672
      | and_dcpl_676);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_99_nl = ~((operator_66_true_div_cmp_z[18])
      | and_dcpl_598 | and_850_cse | and_857_cse | and_dcpl_622 | and_dcpl_628 |
      and_869_cse | and_875_cse | and_dcpl_641 | and_dcpl_646 | and_886_cse | and_dcpl_654
      | and_dcpl_659 | and_dcpl_663 | and_dcpl_666 | and_dcpl_669 | and_dcpl_672
      | and_dcpl_676);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_100_nl = ~((operator_66_true_div_cmp_z[17])
      | and_dcpl_598 | and_850_cse | and_857_cse | and_dcpl_622 | and_dcpl_628 |
      and_869_cse | and_875_cse | and_dcpl_641 | and_dcpl_646 | and_886_cse | and_dcpl_654
      | and_dcpl_659 | and_dcpl_663 | and_dcpl_666 | and_dcpl_669 | and_dcpl_672
      | and_dcpl_676);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_101_nl = ~((operator_66_true_div_cmp_z[16])
      | and_dcpl_598 | and_850_cse | and_857_cse | and_dcpl_622 | and_dcpl_628 |
      and_869_cse | and_875_cse | and_dcpl_641 | and_dcpl_646 | and_886_cse | and_dcpl_654
      | and_dcpl_659 | and_dcpl_663 | and_dcpl_666 | and_dcpl_669 | and_dcpl_672
      | and_dcpl_676);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_102_nl = ~((operator_66_true_div_cmp_z[15])
      | and_dcpl_598 | and_850_cse | and_857_cse | and_dcpl_622 | and_dcpl_628 |
      and_869_cse | and_875_cse | and_dcpl_641 | and_dcpl_646 | and_886_cse | and_dcpl_654
      | and_dcpl_659 | and_dcpl_663 | and_dcpl_666 | and_dcpl_669 | and_dcpl_672
      | and_dcpl_676);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_103_nl = ~((operator_66_true_div_cmp_z[14])
      | and_dcpl_598 | and_850_cse | and_857_cse | and_dcpl_622 | and_dcpl_628 |
      and_869_cse | and_875_cse | and_dcpl_641 | and_dcpl_646 | and_886_cse | and_dcpl_654
      | and_dcpl_659 | and_dcpl_663 | and_dcpl_666 | and_dcpl_669 | and_dcpl_672
      | and_dcpl_676);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_104_nl = ~((operator_66_true_div_cmp_z[13])
      | and_dcpl_598 | and_850_cse | and_857_cse | and_dcpl_622 | and_dcpl_628 |
      and_869_cse | and_875_cse | and_dcpl_641 | and_dcpl_646 | and_886_cse | and_dcpl_654
      | and_dcpl_659 | and_dcpl_663 | and_dcpl_666 | and_dcpl_669 | and_dcpl_672
      | and_dcpl_676);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_105_nl = ~((operator_66_true_div_cmp_z[12])
      | and_dcpl_598 | and_850_cse | and_857_cse | and_dcpl_622 | and_dcpl_628 |
      and_869_cse | and_875_cse | and_dcpl_641 | and_dcpl_646 | and_886_cse | and_dcpl_654
      | and_dcpl_659 | and_dcpl_663 | and_dcpl_666 | and_dcpl_669 | and_dcpl_672
      | and_dcpl_676);
  assign COMP_LOOP_or_79_nl = and_850_cse | and_857_cse | and_dcpl_622 | and_dcpl_628
      | and_869_cse | and_875_cse | and_dcpl_641 | and_dcpl_646 | and_886_cse | and_dcpl_654
      | and_dcpl_659 | and_dcpl_663 | and_dcpl_666 | and_dcpl_669 | and_dcpl_672
      | and_dcpl_676;
  assign COMP_LOOP_mux1h_589_nl = MUX1HOT_v_12_3_2(({6'b000000 , COMP_LOOP_k_9_4_sva_4_0
      , 1'b1}), VEC_LOOP_j_sva_11_0, (~ (operator_66_true_div_cmp_z[11:0])), {and_dcpl_598
      , COMP_LOOP_or_79_nl , and_dcpl_678});
  assign COMP_LOOP_mux1h_590_nl = MUX1HOT_v_7_7_2(({1'b0 , (VEC_LOOP_j_sva_11_0[11:6])}),
      ({(z_out_9[5:0]) , (STAGE_LOOP_lshift_psp_sva[3])}), (z_out_2[9:3]), (z_out_3[9:3]),
      (z_out_4[9:3]), (z_out_1[9:3]), z_out_9, {and_dcpl_598 , and_850_cse , COMP_LOOP_or_55_ssc
      , COMP_LOOP_or_56_ssc , COMP_LOOP_or_57_ssc , COMP_LOOP_or_58_ssc , and_886_cse});
  assign not_8636_nl = ~ and_dcpl_678;
  assign COMP_LOOP_and_285_nl = MUX_v_7_2_2(7'b0000000, COMP_LOOP_mux1h_590_nl, not_8636_nl);
  assign COMP_LOOP_or_80_nl = and_850_cse | and_886_cse;
  assign COMP_LOOP_mux1h_591_nl = MUX1HOT_v_3_7_2((VEC_LOOP_j_sva_11_0[5:3]), (STAGE_LOOP_lshift_psp_sva[2:0]),
      (z_out_2[2:0]), (z_out_3[2:0]), (z_out_4[2:0]), (z_out_1[2:0]), 3'b001, {and_dcpl_598
      , COMP_LOOP_or_80_nl , COMP_LOOP_or_55_ssc , COMP_LOOP_or_56_ssc , COMP_LOOP_or_57_ssc
      , COMP_LOOP_or_58_ssc , and_dcpl_678});
  assign nl_z_out_7 = ({COMP_LOOP_COMP_LOOP_or_21_nl , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_54_nl
      , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_55_nl , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_56_nl
      , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_57_nl , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_58_nl
      , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_59_nl , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_60_nl
      , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_61_nl , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_62_nl
      , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_63_nl , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_64_nl
      , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_65_nl , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_66_nl
      , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_67_nl , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_68_nl
      , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_69_nl , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_70_nl
      , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_71_nl , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_72_nl
      , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_73_nl , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_74_nl
      , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_75_nl , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_76_nl
      , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_77_nl , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_78_nl
      , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_79_nl , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_80_nl
      , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_81_nl , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_82_nl
      , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_83_nl , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_84_nl
      , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_85_nl , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_86_nl
      , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_87_nl , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_88_nl
      , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_89_nl , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_90_nl
      , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_91_nl , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_92_nl
      , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_93_nl , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_94_nl
      , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_95_nl , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_96_nl
      , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_97_nl , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_98_nl
      , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_99_nl , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_100_nl
      , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_101_nl , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_102_nl
      , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_103_nl , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_104_nl
      , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_105_nl , COMP_LOOP_mux1h_589_nl}) + conv_u2u_10_65({COMP_LOOP_and_285_nl
      , COMP_LOOP_mux1h_591_nl});
  assign z_out_7 = nl_z_out_7[64:0];
  assign COMP_LOOP_mux_87_nl = MUX_s_1_2_2((~ modExp_exp_1_7_1_sva), (~ COMP_LOOP_nor_134_itm),
      and_dcpl_707);
  assign COMP_LOOP_COMP_LOOP_or_22_nl = COMP_LOOP_mux_87_nl | and_dcpl_688 | and_dcpl_698;
  assign COMP_LOOP_mux1h_592_nl = MUX1HOT_s_1_3_2((~ (STAGE_LOOP_lshift_psp_sva[9])),
      (~ modExp_exp_1_6_1_sva), (~ modExp_exp_1_7_1_sva), {COMP_LOOP_or_67_itm ,
      not_tmp_980 , and_dcpl_707});
  assign COMP_LOOP_mux1h_593_nl = MUX1HOT_s_1_3_2((~ (STAGE_LOOP_lshift_psp_sva[8])),
      (~ modExp_exp_1_5_1_sva), (~ modExp_exp_1_6_1_sva), {COMP_LOOP_or_67_itm ,
      not_tmp_980 , and_dcpl_707});
  assign COMP_LOOP_mux1h_594_nl = MUX1HOT_s_1_3_2((~ (STAGE_LOOP_lshift_psp_sva[7])),
      (~ modExp_exp_1_4_1_sva), (~ modExp_exp_1_5_1_sva), {COMP_LOOP_or_67_itm ,
      not_tmp_980 , and_dcpl_707});
  assign COMP_LOOP_mux1h_595_nl = MUX1HOT_s_1_3_2((~ (STAGE_LOOP_lshift_psp_sva[6])),
      (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm), (~ modExp_exp_1_4_1_sva), {COMP_LOOP_or_67_itm
      , not_tmp_980 , and_dcpl_707});
  assign COMP_LOOP_mux1h_596_nl = MUX1HOT_s_1_3_2((~ (STAGE_LOOP_lshift_psp_sva[5])),
      (~ COMP_LOOP_nor_137_itm), (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm), {COMP_LOOP_or_67_itm
      , not_tmp_980 , and_dcpl_707});
  assign COMP_LOOP_mux1h_597_nl = MUX1HOT_s_1_3_2((~ (STAGE_LOOP_lshift_psp_sva[4])),
      (~ COMP_LOOP_nor_134_itm), (~ COMP_LOOP_nor_137_itm), {COMP_LOOP_or_67_itm
      , not_tmp_980 , and_dcpl_707});
  assign COMP_LOOP_or_81_nl = not_tmp_980 | and_dcpl_707;
  assign COMP_LOOP_COMP_LOOP_mux_21_nl = MUX_s_1_2_2((~ (STAGE_LOOP_lshift_psp_sva[3])),
      (~ COMP_LOOP_nor_12_itm), COMP_LOOP_or_81_nl);
  assign COMP_LOOP_or_82_nl = COMP_LOOP_nor_680_itm | and_dcpl_688 | and_dcpl_698;
  assign COMP_LOOP_COMP_LOOP_and_990_nl = MUX_v_5_2_2(5'b00000, COMP_LOOP_k_9_4_sva_4_0,
      COMP_LOOP_nor_680_itm);
  assign COMP_LOOP_COMP_LOOP_or_23_nl = (~(and_dcpl_688 | not_tmp_980 | and_dcpl_707))
      | and_dcpl_698;
  assign nl_acc_8_nl = ({COMP_LOOP_COMP_LOOP_or_9_cse , COMP_LOOP_COMP_LOOP_or_22_nl
      , COMP_LOOP_mux1h_592_nl , COMP_LOOP_mux1h_593_nl , COMP_LOOP_mux1h_594_nl
      , COMP_LOOP_mux1h_595_nl , COMP_LOOP_mux1h_596_nl , COMP_LOOP_mux1h_597_nl
      , COMP_LOOP_COMP_LOOP_mux_21_nl , COMP_LOOP_or_82_nl}) + conv_u2u_8_10({COMP_LOOP_COMP_LOOP_and_990_nl
      , COMP_LOOP_COMP_LOOP_or_23_nl , COMP_LOOP_COMP_LOOP_or_9_cse , 1'b1});
  assign acc_8_nl = nl_acc_8_nl[9:0];
  assign z_out_8_8_7 = readslicef_10_2_8(acc_8_nl);
  assign COMP_LOOP_COMP_LOOP_or_24_nl = ((STAGE_LOOP_lshift_psp_sva[9]) & (~(and_dcpl_727
      | and_dcpl_734))) | and_dcpl_717;
  assign COMP_LOOP_mux1h_598_nl = MUX1HOT_v_6_4_2((~ (STAGE_LOOP_lshift_psp_sva[9:4])),
      ({1'b1 , (~ (STAGE_LOOP_lshift_psp_sva[9:5]))}), (STAGE_LOOP_lshift_psp_sva[9:4]),
      (STAGE_LOOP_lshift_psp_sva[8:3]), {and_dcpl_717 , and_dcpl_727 , and_dcpl_734
      , and_dcpl_741});
  assign COMP_LOOP_or_83_nl = (~(and_dcpl_734 | and_dcpl_741)) | and_dcpl_717 | and_dcpl_727;
  assign COMP_LOOP_or_84_nl = and_dcpl_727 | and_dcpl_734;
  assign COMP_LOOP_COMP_LOOP_mux_22_nl = MUX_v_5_2_2(COMP_LOOP_k_9_4_sva_4_0, ({1'b0
      , (COMP_LOOP_k_9_4_sva_4_0[4:1])}), COMP_LOOP_or_84_nl);
  assign COMP_LOOP_COMP_LOOP_or_25_nl = ((COMP_LOOP_k_9_4_sva_4_0[0]) & (~ and_dcpl_717))
      | and_dcpl_741;
  assign nl_acc_9_nl = ({COMP_LOOP_COMP_LOOP_or_24_nl , COMP_LOOP_mux1h_598_nl ,
      COMP_LOOP_or_83_nl}) + conv_u2u_7_8({COMP_LOOP_COMP_LOOP_mux_22_nl , COMP_LOOP_COMP_LOOP_or_25_nl
      , 1'b1});
  assign acc_9_nl = nl_acc_9_nl[7:0];
  assign z_out_9 = readslicef_8_7_1(acc_9_nl);
  assign nor_1463_nl = ~((~ (fsm_output[5])) | (~ (fsm_output[9])) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (fsm_output[8]) | (fsm_output[6]));
  assign nor_1464_nl = ~((~ (fsm_output[5])) | (fsm_output[9]) | (fsm_output[2])
      | (fsm_output[3]) | nand_257_cse);
  assign mux_3958_nl = MUX_s_1_2_2(nor_1463_nl, nor_1464_nl, fsm_output[1]);
  assign nor_1465_nl = ~((fsm_output[1]) | (~ (fsm_output[5])) | (fsm_output[9])
      | (~ (fsm_output[2])) | (fsm_output[3]) | (fsm_output[8]) | (fsm_output[6]));
  assign mux_3957_nl = MUX_s_1_2_2(mux_3958_nl, nor_1465_nl, fsm_output[4]);
  assign nor_1466_nl = ~((fsm_output[1]) | (fsm_output[5]) | (~ (fsm_output[9]))
      | (fsm_output[2]) | (fsm_output[3]) | nand_257_cse);
  assign nor_1467_nl = ~((fsm_output[5]) | (fsm_output[9]) | (fsm_output[2]) | (~
      (fsm_output[3])) | (fsm_output[8]) | (fsm_output[6]));
  assign nor_1468_nl = ~((~ (fsm_output[5])) | (~ (fsm_output[9])) | (~ (fsm_output[2]))
      | (fsm_output[3]) | (fsm_output[8]) | (~ (fsm_output[6])));
  assign mux_3960_nl = MUX_s_1_2_2(nor_1467_nl, nor_1468_nl, fsm_output[1]);
  assign mux_3959_nl = MUX_s_1_2_2(nor_1466_nl, mux_3960_nl, fsm_output[4]);
  assign mux_3956_nl = MUX_s_1_2_2(mux_3957_nl, mux_3959_nl, fsm_output[7]);
  assign nor_1469_nl = ~((~ (fsm_output[1])) | (fsm_output[5]) | (fsm_output[9])
      | (fsm_output[2]) | (~ (fsm_output[3])) | (fsm_output[8]) | (fsm_output[6]));
  assign nor_1470_nl = ~((~ (fsm_output[1])) | (fsm_output[5]) | (~ (fsm_output[9]))
      | (fsm_output[2]) | (~((fsm_output[3]) & (fsm_output[8]) & (fsm_output[6]))));
  assign mux_3962_nl = MUX_s_1_2_2(nor_1469_nl, nor_1470_nl, fsm_output[4]);
  assign nor_1471_nl = ~((~ (fsm_output[1])) | (fsm_output[5]) | (fsm_output[9])
      | (~ (fsm_output[2])) | (fsm_output[3]) | nand_257_cse);
  assign or_3612_nl = (~ (fsm_output[9])) | (fsm_output[2]) | (fsm_output[3]) | (fsm_output[8])
      | (fsm_output[6]);
  assign or_3613_nl = (fsm_output[9]) | (~ (fsm_output[2])) | (~ (fsm_output[3]))
      | (fsm_output[8]) | (~ (fsm_output[6]));
  assign mux_3964_nl = MUX_s_1_2_2(or_3612_nl, or_3613_nl, fsm_output[5]);
  assign nor_1472_nl = ~((fsm_output[1]) | mux_3964_nl);
  assign mux_3963_nl = MUX_s_1_2_2(nor_1471_nl, nor_1472_nl, fsm_output[4]);
  assign mux_3961_nl = MUX_s_1_2_2(mux_3962_nl, mux_3963_nl, fsm_output[7]);
  assign mux_3955_nl = MUX_s_1_2_2(mux_3956_nl, mux_3961_nl, fsm_output[0]);
  assign nor_1473_nl = ~((fsm_output[5]) | (fsm_output[9]) | (~ (fsm_output[2]))
      | (fsm_output[3]) | nand_257_cse);
  assign nor_1474_nl = ~((fsm_output[5]) | (~ (fsm_output[9])) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (fsm_output[8]) | (fsm_output[6]));
  assign mux_3967_nl = MUX_s_1_2_2(nor_1473_nl, nor_1474_nl, fsm_output[1]);
  assign and_1286_nl = (fsm_output[4]) & mux_3967_nl;
  assign nor_1475_nl = ~((fsm_output[4]) | (~ (fsm_output[1])) | (fsm_output[5])
      | (fsm_output[9]) | (fsm_output[2]) | (~ (fsm_output[3])) | (fsm_output[8])
      | (fsm_output[6]));
  assign mux_3966_nl = MUX_s_1_2_2(and_1286_nl, nor_1475_nl, fsm_output[7]);
  assign nor_1476_nl = ~((fsm_output[4]) | (fsm_output[1]) | (~ (fsm_output[5]))
      | (fsm_output[9]) | (~ (fsm_output[2])) | (fsm_output[3]) | (fsm_output[8])
      | (fsm_output[6]));
  assign and_1287_nl = (fsm_output[1]) & (fsm_output[5]) & (~ (fsm_output[9])) &
      (fsm_output[2]) & (fsm_output[3]) & (~ (fsm_output[8])) & (fsm_output[6]);
  assign nor_1477_nl = ~((fsm_output[1]) | (~ (fsm_output[5])) | (fsm_output[9])
      | (fsm_output[2]) | (~ (fsm_output[3])) | (~ (fsm_output[8])) | (fsm_output[6]));
  assign mux_3969_nl = MUX_s_1_2_2(and_1287_nl, nor_1477_nl, fsm_output[4]);
  assign mux_3968_nl = MUX_s_1_2_2(nor_1476_nl, mux_3969_nl, fsm_output[7]);
  assign mux_3965_nl = MUX_s_1_2_2(mux_3966_nl, mux_3968_nl, fsm_output[0]);
  assign mux_3954_nl = MUX_s_1_2_2(mux_3955_nl, mux_3965_nl, fsm_output[10]);
  assign modExp_while_if_mux_1_nl = MUX_v_64_2_2(modExp_result_sva, COMP_LOOP_10_mul_mut,
      mux_3954_nl);
  assign nl_z_out_10 = $signed(conv_u2s_64_65(modExp_while_if_mux_1_nl)) * $signed(COMP_LOOP_10_mul_mut);
  assign z_out_10 = nl_z_out_10[63:0];

  function automatic [0:0] MUX1HOT_s_1_3_2;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [2:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function automatic [0:0] MUX1HOT_s_1_4_2;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [3:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    MUX1HOT_s_1_4_2 = result;
  end
  endfunction


  function automatic [0:0] MUX1HOT_s_1_6_2;
    input [0:0] input_5;
    input [0:0] input_4;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [5:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    result = result | ( input_4 & {1{sel[4]}});
    result = result | ( input_5 & {1{sel[5]}});
    MUX1HOT_s_1_6_2 = result;
  end
  endfunction


  function automatic [11:0] MUX1HOT_v_12_3_2;
    input [11:0] input_2;
    input [11:0] input_1;
    input [11:0] input_0;
    input [2:0] sel;
    reg [11:0] result;
  begin
    result = input_0 & {12{sel[0]}};
    result = result | ( input_1 & {12{sel[1]}});
    result = result | ( input_2 & {12{sel[2]}});
    MUX1HOT_v_12_3_2 = result;
  end
  endfunction


  function automatic [2:0] MUX1HOT_v_3_7_2;
    input [2:0] input_6;
    input [2:0] input_5;
    input [2:0] input_4;
    input [2:0] input_3;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [6:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | ( input_1 & {3{sel[1]}});
    result = result | ( input_2 & {3{sel[2]}});
    result = result | ( input_3 & {3{sel[3]}});
    result = result | ( input_4 & {3{sel[4]}});
    result = result | ( input_5 & {3{sel[5]}});
    result = result | ( input_6 & {3{sel[6]}});
    MUX1HOT_v_3_7_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_4_2;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [3:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | ( input_1 & {4{sel[1]}});
    result = result | ( input_2 & {4{sel[2]}});
    result = result | ( input_3 & {4{sel[3]}});
    MUX1HOT_v_4_4_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_17_2;
    input [63:0] input_16;
    input [63:0] input_15;
    input [63:0] input_14;
    input [63:0] input_13;
    input [63:0] input_12;
    input [63:0] input_11;
    input [63:0] input_10;
    input [63:0] input_9;
    input [63:0] input_8;
    input [63:0] input_7;
    input [63:0] input_6;
    input [63:0] input_5;
    input [63:0] input_4;
    input [63:0] input_3;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [16:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    result = result | ( input_3 & {64{sel[3]}});
    result = result | ( input_4 & {64{sel[4]}});
    result = result | ( input_5 & {64{sel[5]}});
    result = result | ( input_6 & {64{sel[6]}});
    result = result | ( input_7 & {64{sel[7]}});
    result = result | ( input_8 & {64{sel[8]}});
    result = result | ( input_9 & {64{sel[9]}});
    result = result | ( input_10 & {64{sel[10]}});
    result = result | ( input_11 & {64{sel[11]}});
    result = result | ( input_12 & {64{sel[12]}});
    result = result | ( input_13 & {64{sel[13]}});
    result = result | ( input_14 & {64{sel[14]}});
    result = result | ( input_15 & {64{sel[15]}});
    result = result | ( input_16 & {64{sel[16]}});
    MUX1HOT_v_64_17_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_21_2;
    input [63:0] input_20;
    input [63:0] input_19;
    input [63:0] input_18;
    input [63:0] input_17;
    input [63:0] input_16;
    input [63:0] input_15;
    input [63:0] input_14;
    input [63:0] input_13;
    input [63:0] input_12;
    input [63:0] input_11;
    input [63:0] input_10;
    input [63:0] input_9;
    input [63:0] input_8;
    input [63:0] input_7;
    input [63:0] input_6;
    input [63:0] input_5;
    input [63:0] input_4;
    input [63:0] input_3;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [20:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    result = result | ( input_3 & {64{sel[3]}});
    result = result | ( input_4 & {64{sel[4]}});
    result = result | ( input_5 & {64{sel[5]}});
    result = result | ( input_6 & {64{sel[6]}});
    result = result | ( input_7 & {64{sel[7]}});
    result = result | ( input_8 & {64{sel[8]}});
    result = result | ( input_9 & {64{sel[9]}});
    result = result | ( input_10 & {64{sel[10]}});
    result = result | ( input_11 & {64{sel[11]}});
    result = result | ( input_12 & {64{sel[12]}});
    result = result | ( input_13 & {64{sel[13]}});
    result = result | ( input_14 & {64{sel[14]}});
    result = result | ( input_15 & {64{sel[15]}});
    result = result | ( input_16 & {64{sel[16]}});
    result = result | ( input_17 & {64{sel[17]}});
    result = result | ( input_18 & {64{sel[18]}});
    result = result | ( input_19 & {64{sel[19]}});
    result = result | ( input_20 & {64{sel[20]}});
    MUX1HOT_v_64_21_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_3_2;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [2:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    MUX1HOT_v_64_3_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_4_2;
    input [63:0] input_3;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [3:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    result = result | ( input_3 & {64{sel[3]}});
    MUX1HOT_v_64_4_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_6_2;
    input [63:0] input_5;
    input [63:0] input_4;
    input [63:0] input_3;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [5:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    result = result | ( input_3 & {64{sel[3]}});
    result = result | ( input_4 & {64{sel[4]}});
    result = result | ( input_5 & {64{sel[5]}});
    MUX1HOT_v_64_6_2 = result;
  end
  endfunction


  function automatic [64:0] MUX1HOT_v_65_3_2;
    input [64:0] input_2;
    input [64:0] input_1;
    input [64:0] input_0;
    input [2:0] sel;
    reg [64:0] result;
  begin
    result = input_0 & {65{sel[0]}};
    result = result | ( input_1 & {65{sel[1]}});
    result = result | ( input_2 & {65{sel[2]}});
    MUX1HOT_v_65_3_2 = result;
  end
  endfunction


  function automatic [5:0] MUX1HOT_v_6_4_2;
    input [5:0] input_3;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [3:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | ( input_1 & {6{sel[1]}});
    result = result | ( input_2 & {6{sel[2]}});
    result = result | ( input_3 & {6{sel[3]}});
    MUX1HOT_v_6_4_2 = result;
  end
  endfunction


  function automatic [6:0] MUX1HOT_v_7_7_2;
    input [6:0] input_6;
    input [6:0] input_5;
    input [6:0] input_4;
    input [6:0] input_3;
    input [6:0] input_2;
    input [6:0] input_1;
    input [6:0] input_0;
    input [6:0] sel;
    reg [6:0] result;
  begin
    result = input_0 & {7{sel[0]}};
    result = result | ( input_1 & {7{sel[1]}});
    result = result | ( input_2 & {7{sel[2]}});
    result = result | ( input_3 & {7{sel[3]}});
    result = result | ( input_4 & {7{sel[4]}});
    result = result | ( input_5 & {7{sel[5]}});
    result = result | ( input_6 & {7{sel[6]}});
    MUX1HOT_v_7_7_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_19_2;
    input [7:0] input_18;
    input [7:0] input_17;
    input [7:0] input_16;
    input [7:0] input_15;
    input [7:0] input_14;
    input [7:0] input_13;
    input [7:0] input_12;
    input [7:0] input_11;
    input [7:0] input_10;
    input [7:0] input_9;
    input [7:0] input_8;
    input [7:0] input_7;
    input [7:0] input_6;
    input [7:0] input_5;
    input [7:0] input_4;
    input [7:0] input_3;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [18:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | ( input_1 & {8{sel[1]}});
    result = result | ( input_2 & {8{sel[2]}});
    result = result | ( input_3 & {8{sel[3]}});
    result = result | ( input_4 & {8{sel[4]}});
    result = result | ( input_5 & {8{sel[5]}});
    result = result | ( input_6 & {8{sel[6]}});
    result = result | ( input_7 & {8{sel[7]}});
    result = result | ( input_8 & {8{sel[8]}});
    result = result | ( input_9 & {8{sel[9]}});
    result = result | ( input_10 & {8{sel[10]}});
    result = result | ( input_11 & {8{sel[11]}});
    result = result | ( input_12 & {8{sel[12]}});
    result = result | ( input_13 & {8{sel[13]}});
    result = result | ( input_14 & {8{sel[14]}});
    result = result | ( input_15 & {8{sel[15]}});
    result = result | ( input_16 & {8{sel[16]}});
    result = result | ( input_17 & {8{sel[17]}});
    result = result | ( input_18 & {8{sel[18]}});
    MUX1HOT_v_8_19_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [9:0] MUX_v_10_2_2;
    input [9:0] input_0;
    input [9:0] input_1;
    input [0:0] sel;
    reg [9:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_10_2_2 = result;
  end
  endfunction


  function automatic [11:0] MUX_v_12_2_2;
    input [11:0] input_0;
    input [11:0] input_1;
    input [0:0] sel;
    reg [11:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_12_2_2 = result;
  end
  endfunction


  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input [0:0] sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [0:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [4:0] MUX_v_5_2_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input [0:0] sel;
    reg [4:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_5_2_2 = result;
  end
  endfunction


  function automatic [62:0] MUX_v_63_2_2;
    input [62:0] input_0;
    input [62:0] input_1;
    input [0:0] sel;
    reg [62:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_63_2_2 = result;
  end
  endfunction


  function automatic [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function automatic [64:0] MUX_v_65_2_2;
    input [64:0] input_0;
    input [64:0] input_1;
    input [0:0] sel;
    reg [64:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_65_2_2 = result;
  end
  endfunction


  function automatic [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input [0:0] sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function automatic [8:0] MUX_v_9_2_2;
    input [8:0] input_0;
    input [8:0] input_1;
    input [0:0] sel;
    reg [8:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_9_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_10_1_9;
    input [9:0] vector;
    reg [9:0] tmp;
  begin
    tmp = vector >> 9;
    readslicef_10_1_9 = tmp[0:0];
  end
  endfunction


  function automatic [1:0] readslicef_10_2_8;
    input [9:0] vector;
    reg [9:0] tmp;
  begin
    tmp = vector >> 8;
    readslicef_10_2_8 = tmp[1:0];
  end
  endfunction


  function automatic [9:0] readslicef_11_10_1;
    input [10:0] vector;
    reg [10:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_11_10_1 = tmp[9:0];
  end
  endfunction


  function automatic [0:0] readslicef_3_1_2;
    input [2:0] vector;
    reg [2:0] tmp;
  begin
    tmp = vector >> 2;
    readslicef_3_1_2 = tmp[0:0];
  end
  endfunction


  function automatic [6:0] readslicef_8_7_1;
    input [7:0] vector;
    reg [7:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_8_7_1 = tmp[6:0];
  end
  endfunction


  function automatic [64:0] conv_s2u_64_65 ;
    input [63:0]  vector ;
  begin
    conv_s2u_64_65 = {vector[63], vector};
  end
  endfunction


  function automatic [64:0] conv_u2s_64_65 ;
    input [63:0]  vector ;
  begin
    conv_u2s_64_65 =  {1'b0, vector};
  end
  endfunction


  function automatic [5:0] conv_u2u_5_6 ;
    input [4:0]  vector ;
  begin
    conv_u2u_5_6 = {1'b0, vector};
  end
  endfunction


  function automatic [7:0] conv_u2u_5_8 ;
    input [4:0]  vector ;
  begin
    conv_u2u_5_8 = {{3{1'b0}}, vector};
  end
  endfunction


  function automatic [7:0] conv_u2u_7_8 ;
    input [6:0]  vector ;
  begin
    conv_u2u_7_8 = {1'b0, vector};
  end
  endfunction


  function automatic [9:0] conv_u2u_8_10 ;
    input [7:0]  vector ;
  begin
    conv_u2u_8_10 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [10:0] conv_u2u_8_11 ;
    input [7:0]  vector ;
  begin
    conv_u2u_8_11 = {{3{1'b0}}, vector};
  end
  endfunction


  function automatic [9:0] conv_u2u_9_10 ;
    input [8:0]  vector ;
  begin
    conv_u2u_9_10 = {1'b0, vector};
  end
  endfunction


  function automatic [11:0] conv_u2u_9_12 ;
    input [8:0]  vector ;
  begin
    conv_u2u_9_12 = {{3{1'b0}}, vector};
  end
  endfunction


  function automatic [10:0] conv_u2u_10_11 ;
    input [9:0]  vector ;
  begin
    conv_u2u_10_11 = {1'b0, vector};
  end
  endfunction


  function automatic [64:0] conv_u2u_10_65 ;
    input [9:0]  vector ;
  begin
    conv_u2u_10_65 = {{55{1'b0}}, vector};
  end
  endfunction


  function automatic [64:0] conv_u2u_64_65 ;
    input [63:0]  vector ;
  begin
    conv_u2u_64_65 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT
// ------------------------------------------------------------------


module inPlaceNTT_DIT (
  clk, rst, vec_rsc_0_0_adra, vec_rsc_0_0_da, vec_rsc_0_0_wea, vec_rsc_0_0_qa, vec_rsc_triosy_0_0_lz,
      vec_rsc_0_1_adra, vec_rsc_0_1_da, vec_rsc_0_1_wea, vec_rsc_0_1_qa, vec_rsc_triosy_0_1_lz,
      vec_rsc_0_2_adra, vec_rsc_0_2_da, vec_rsc_0_2_wea, vec_rsc_0_2_qa, vec_rsc_triosy_0_2_lz,
      vec_rsc_0_3_adra, vec_rsc_0_3_da, vec_rsc_0_3_wea, vec_rsc_0_3_qa, vec_rsc_triosy_0_3_lz,
      vec_rsc_0_4_adra, vec_rsc_0_4_da, vec_rsc_0_4_wea, vec_rsc_0_4_qa, vec_rsc_triosy_0_4_lz,
      vec_rsc_0_5_adra, vec_rsc_0_5_da, vec_rsc_0_5_wea, vec_rsc_0_5_qa, vec_rsc_triosy_0_5_lz,
      vec_rsc_0_6_adra, vec_rsc_0_6_da, vec_rsc_0_6_wea, vec_rsc_0_6_qa, vec_rsc_triosy_0_6_lz,
      vec_rsc_0_7_adra, vec_rsc_0_7_da, vec_rsc_0_7_wea, vec_rsc_0_7_qa, vec_rsc_triosy_0_7_lz,
      vec_rsc_0_8_adra, vec_rsc_0_8_da, vec_rsc_0_8_wea, vec_rsc_0_8_qa, vec_rsc_triosy_0_8_lz,
      vec_rsc_0_9_adra, vec_rsc_0_9_da, vec_rsc_0_9_wea, vec_rsc_0_9_qa, vec_rsc_triosy_0_9_lz,
      vec_rsc_0_10_adra, vec_rsc_0_10_da, vec_rsc_0_10_wea, vec_rsc_0_10_qa, vec_rsc_triosy_0_10_lz,
      vec_rsc_0_11_adra, vec_rsc_0_11_da, vec_rsc_0_11_wea, vec_rsc_0_11_qa, vec_rsc_triosy_0_11_lz,
      vec_rsc_0_12_adra, vec_rsc_0_12_da, vec_rsc_0_12_wea, vec_rsc_0_12_qa, vec_rsc_triosy_0_12_lz,
      vec_rsc_0_13_adra, vec_rsc_0_13_da, vec_rsc_0_13_wea, vec_rsc_0_13_qa, vec_rsc_triosy_0_13_lz,
      vec_rsc_0_14_adra, vec_rsc_0_14_da, vec_rsc_0_14_wea, vec_rsc_0_14_qa, vec_rsc_triosy_0_14_lz,
      vec_rsc_0_15_adra, vec_rsc_0_15_da, vec_rsc_0_15_wea, vec_rsc_0_15_qa, vec_rsc_triosy_0_15_lz,
      p_rsc_dat, p_rsc_triosy_lz, r_rsc_dat, r_rsc_triosy_lz
);
  input clk;
  input rst;
  output [7:0] vec_rsc_0_0_adra;
  output [63:0] vec_rsc_0_0_da;
  output vec_rsc_0_0_wea;
  input [63:0] vec_rsc_0_0_qa;
  output vec_rsc_triosy_0_0_lz;
  output [7:0] vec_rsc_0_1_adra;
  output [63:0] vec_rsc_0_1_da;
  output vec_rsc_0_1_wea;
  input [63:0] vec_rsc_0_1_qa;
  output vec_rsc_triosy_0_1_lz;
  output [7:0] vec_rsc_0_2_adra;
  output [63:0] vec_rsc_0_2_da;
  output vec_rsc_0_2_wea;
  input [63:0] vec_rsc_0_2_qa;
  output vec_rsc_triosy_0_2_lz;
  output [7:0] vec_rsc_0_3_adra;
  output [63:0] vec_rsc_0_3_da;
  output vec_rsc_0_3_wea;
  input [63:0] vec_rsc_0_3_qa;
  output vec_rsc_triosy_0_3_lz;
  output [7:0] vec_rsc_0_4_adra;
  output [63:0] vec_rsc_0_4_da;
  output vec_rsc_0_4_wea;
  input [63:0] vec_rsc_0_4_qa;
  output vec_rsc_triosy_0_4_lz;
  output [7:0] vec_rsc_0_5_adra;
  output [63:0] vec_rsc_0_5_da;
  output vec_rsc_0_5_wea;
  input [63:0] vec_rsc_0_5_qa;
  output vec_rsc_triosy_0_5_lz;
  output [7:0] vec_rsc_0_6_adra;
  output [63:0] vec_rsc_0_6_da;
  output vec_rsc_0_6_wea;
  input [63:0] vec_rsc_0_6_qa;
  output vec_rsc_triosy_0_6_lz;
  output [7:0] vec_rsc_0_7_adra;
  output [63:0] vec_rsc_0_7_da;
  output vec_rsc_0_7_wea;
  input [63:0] vec_rsc_0_7_qa;
  output vec_rsc_triosy_0_7_lz;
  output [7:0] vec_rsc_0_8_adra;
  output [63:0] vec_rsc_0_8_da;
  output vec_rsc_0_8_wea;
  input [63:0] vec_rsc_0_8_qa;
  output vec_rsc_triosy_0_8_lz;
  output [7:0] vec_rsc_0_9_adra;
  output [63:0] vec_rsc_0_9_da;
  output vec_rsc_0_9_wea;
  input [63:0] vec_rsc_0_9_qa;
  output vec_rsc_triosy_0_9_lz;
  output [7:0] vec_rsc_0_10_adra;
  output [63:0] vec_rsc_0_10_da;
  output vec_rsc_0_10_wea;
  input [63:0] vec_rsc_0_10_qa;
  output vec_rsc_triosy_0_10_lz;
  output [7:0] vec_rsc_0_11_adra;
  output [63:0] vec_rsc_0_11_da;
  output vec_rsc_0_11_wea;
  input [63:0] vec_rsc_0_11_qa;
  output vec_rsc_triosy_0_11_lz;
  output [7:0] vec_rsc_0_12_adra;
  output [63:0] vec_rsc_0_12_da;
  output vec_rsc_0_12_wea;
  input [63:0] vec_rsc_0_12_qa;
  output vec_rsc_triosy_0_12_lz;
  output [7:0] vec_rsc_0_13_adra;
  output [63:0] vec_rsc_0_13_da;
  output vec_rsc_0_13_wea;
  input [63:0] vec_rsc_0_13_qa;
  output vec_rsc_triosy_0_13_lz;
  output [7:0] vec_rsc_0_14_adra;
  output [63:0] vec_rsc_0_14_da;
  output vec_rsc_0_14_wea;
  input [63:0] vec_rsc_0_14_qa;
  output vec_rsc_triosy_0_14_lz;
  output [7:0] vec_rsc_0_15_adra;
  output [63:0] vec_rsc_0_15_da;
  output vec_rsc_0_15_wea;
  input [63:0] vec_rsc_0_15_qa;
  output vec_rsc_triosy_0_15_lz;
  input [63:0] p_rsc_dat;
  output p_rsc_triosy_lz;
  input [63:0] r_rsc_dat;
  output r_rsc_triosy_lz;


  // Interconnect Declarations
  wire [63:0] vec_rsc_0_0_i_qa_d;
  wire vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_1_i_qa_d;
  wire vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_2_i_qa_d;
  wire vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_3_i_qa_d;
  wire vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_4_i_qa_d;
  wire vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_5_i_qa_d;
  wire vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_6_i_qa_d;
  wire vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_7_i_qa_d;
  wire vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_8_i_qa_d;
  wire vec_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_9_i_qa_d;
  wire vec_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_10_i_qa_d;
  wire vec_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_11_i_qa_d;
  wire vec_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_12_i_qa_d;
  wire vec_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_13_i_qa_d;
  wire vec_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_14_i_qa_d;
  wire vec_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_15_i_qa_d;
  wire vec_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] vec_rsc_0_0_i_adra_d_iff;
  wire [63:0] vec_rsc_0_0_i_da_d_iff;
  wire vec_rsc_0_0_i_wea_d_iff;
  wire vec_rsc_0_1_i_wea_d_iff;
  wire vec_rsc_0_2_i_wea_d_iff;
  wire vec_rsc_0_3_i_wea_d_iff;
  wire vec_rsc_0_4_i_wea_d_iff;
  wire vec_rsc_0_5_i_wea_d_iff;
  wire vec_rsc_0_6_i_wea_d_iff;
  wire vec_rsc_0_7_i_wea_d_iff;
  wire vec_rsc_0_8_i_wea_d_iff;
  wire vec_rsc_0_9_i_wea_d_iff;
  wire vec_rsc_0_10_i_wea_d_iff;
  wire vec_rsc_0_11_i_wea_d_iff;
  wire vec_rsc_0_12_i_wea_d_iff;
  wire vec_rsc_0_13_i_wea_d_iff;
  wire vec_rsc_0_14_i_wea_d_iff;
  wire vec_rsc_0_15_i_wea_d_iff;


  // Interconnect Declarations for Component Instantiations 
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_4_8_64_256_256_64_1_gen vec_rsc_0_0_i
      (
      .qa(vec_rsc_0_0_qa),
      .wea(vec_rsc_0_0_wea),
      .da(vec_rsc_0_0_da),
      .adra(vec_rsc_0_0_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_0_i_qa_d),
      .wea_d(vec_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_0_i_wea_d_iff)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_5_8_64_256_256_64_1_gen vec_rsc_0_1_i
      (
      .qa(vec_rsc_0_1_qa),
      .wea(vec_rsc_0_1_wea),
      .da(vec_rsc_0_1_da),
      .adra(vec_rsc_0_1_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_1_i_qa_d),
      .wea_d(vec_rsc_0_1_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_1_i_wea_d_iff)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_6_8_64_256_256_64_1_gen vec_rsc_0_2_i
      (
      .qa(vec_rsc_0_2_qa),
      .wea(vec_rsc_0_2_wea),
      .da(vec_rsc_0_2_da),
      .adra(vec_rsc_0_2_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_2_i_qa_d),
      .wea_d(vec_rsc_0_2_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_2_i_wea_d_iff)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_7_8_64_256_256_64_1_gen vec_rsc_0_3_i
      (
      .qa(vec_rsc_0_3_qa),
      .wea(vec_rsc_0_3_wea),
      .da(vec_rsc_0_3_da),
      .adra(vec_rsc_0_3_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_3_i_qa_d),
      .wea_d(vec_rsc_0_3_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_3_i_wea_d_iff)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_8_8_64_256_256_64_1_gen vec_rsc_0_4_i
      (
      .qa(vec_rsc_0_4_qa),
      .wea(vec_rsc_0_4_wea),
      .da(vec_rsc_0_4_da),
      .adra(vec_rsc_0_4_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_4_i_qa_d),
      .wea_d(vec_rsc_0_4_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_4_i_wea_d_iff)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_9_8_64_256_256_64_1_gen vec_rsc_0_5_i
      (
      .qa(vec_rsc_0_5_qa),
      .wea(vec_rsc_0_5_wea),
      .da(vec_rsc_0_5_da),
      .adra(vec_rsc_0_5_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_5_i_qa_d),
      .wea_d(vec_rsc_0_5_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_5_i_wea_d_iff)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_10_8_64_256_256_64_1_gen
      vec_rsc_0_6_i (
      .qa(vec_rsc_0_6_qa),
      .wea(vec_rsc_0_6_wea),
      .da(vec_rsc_0_6_da),
      .adra(vec_rsc_0_6_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_6_i_qa_d),
      .wea_d(vec_rsc_0_6_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_6_i_wea_d_iff)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_11_8_64_256_256_64_1_gen
      vec_rsc_0_7_i (
      .qa(vec_rsc_0_7_qa),
      .wea(vec_rsc_0_7_wea),
      .da(vec_rsc_0_7_da),
      .adra(vec_rsc_0_7_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_7_i_qa_d),
      .wea_d(vec_rsc_0_7_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_7_i_wea_d_iff)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_12_8_64_256_256_64_1_gen
      vec_rsc_0_8_i (
      .qa(vec_rsc_0_8_qa),
      .wea(vec_rsc_0_8_wea),
      .da(vec_rsc_0_8_da),
      .adra(vec_rsc_0_8_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_8_i_qa_d),
      .wea_d(vec_rsc_0_8_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_8_i_wea_d_iff)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_13_8_64_256_256_64_1_gen
      vec_rsc_0_9_i (
      .qa(vec_rsc_0_9_qa),
      .wea(vec_rsc_0_9_wea),
      .da(vec_rsc_0_9_da),
      .adra(vec_rsc_0_9_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_9_i_qa_d),
      .wea_d(vec_rsc_0_9_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_9_i_wea_d_iff)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_14_8_64_256_256_64_1_gen
      vec_rsc_0_10_i (
      .qa(vec_rsc_0_10_qa),
      .wea(vec_rsc_0_10_wea),
      .da(vec_rsc_0_10_da),
      .adra(vec_rsc_0_10_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_10_i_qa_d),
      .wea_d(vec_rsc_0_10_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_10_i_wea_d_iff)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_15_8_64_256_256_64_1_gen
      vec_rsc_0_11_i (
      .qa(vec_rsc_0_11_qa),
      .wea(vec_rsc_0_11_wea),
      .da(vec_rsc_0_11_da),
      .adra(vec_rsc_0_11_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_11_i_qa_d),
      .wea_d(vec_rsc_0_11_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_11_i_wea_d_iff)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_16_8_64_256_256_64_1_gen
      vec_rsc_0_12_i (
      .qa(vec_rsc_0_12_qa),
      .wea(vec_rsc_0_12_wea),
      .da(vec_rsc_0_12_da),
      .adra(vec_rsc_0_12_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_12_i_qa_d),
      .wea_d(vec_rsc_0_12_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_12_i_wea_d_iff)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_17_8_64_256_256_64_1_gen
      vec_rsc_0_13_i (
      .qa(vec_rsc_0_13_qa),
      .wea(vec_rsc_0_13_wea),
      .da(vec_rsc_0_13_da),
      .adra(vec_rsc_0_13_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_13_i_qa_d),
      .wea_d(vec_rsc_0_13_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_13_i_wea_d_iff)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_18_8_64_256_256_64_1_gen
      vec_rsc_0_14_i (
      .qa(vec_rsc_0_14_qa),
      .wea(vec_rsc_0_14_wea),
      .da(vec_rsc_0_14_da),
      .adra(vec_rsc_0_14_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_14_i_qa_d),
      .wea_d(vec_rsc_0_14_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_14_i_wea_d_iff)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_19_8_64_256_256_64_1_gen
      vec_rsc_0_15_i (
      .qa(vec_rsc_0_15_qa),
      .wea(vec_rsc_0_15_wea),
      .da(vec_rsc_0_15_da),
      .adra(vec_rsc_0_15_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_15_i_qa_d),
      .wea_d(vec_rsc_0_15_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_15_i_wea_d_iff)
    );
  inPlaceNTT_DIT_core inPlaceNTT_DIT_core_inst (
      .clk(clk),
      .rst(rst),
      .vec_rsc_triosy_0_0_lz(vec_rsc_triosy_0_0_lz),
      .vec_rsc_triosy_0_1_lz(vec_rsc_triosy_0_1_lz),
      .vec_rsc_triosy_0_2_lz(vec_rsc_triosy_0_2_lz),
      .vec_rsc_triosy_0_3_lz(vec_rsc_triosy_0_3_lz),
      .vec_rsc_triosy_0_4_lz(vec_rsc_triosy_0_4_lz),
      .vec_rsc_triosy_0_5_lz(vec_rsc_triosy_0_5_lz),
      .vec_rsc_triosy_0_6_lz(vec_rsc_triosy_0_6_lz),
      .vec_rsc_triosy_0_7_lz(vec_rsc_triosy_0_7_lz),
      .vec_rsc_triosy_0_8_lz(vec_rsc_triosy_0_8_lz),
      .vec_rsc_triosy_0_9_lz(vec_rsc_triosy_0_9_lz),
      .vec_rsc_triosy_0_10_lz(vec_rsc_triosy_0_10_lz),
      .vec_rsc_triosy_0_11_lz(vec_rsc_triosy_0_11_lz),
      .vec_rsc_triosy_0_12_lz(vec_rsc_triosy_0_12_lz),
      .vec_rsc_triosy_0_13_lz(vec_rsc_triosy_0_13_lz),
      .vec_rsc_triosy_0_14_lz(vec_rsc_triosy_0_14_lz),
      .vec_rsc_triosy_0_15_lz(vec_rsc_triosy_0_15_lz),
      .p_rsc_dat(p_rsc_dat),
      .p_rsc_triosy_lz(p_rsc_triosy_lz),
      .r_rsc_dat(r_rsc_dat),
      .r_rsc_triosy_lz(r_rsc_triosy_lz),
      .vec_rsc_0_0_i_qa_d(vec_rsc_0_0_i_qa_d),
      .vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_1_i_qa_d(vec_rsc_0_1_i_qa_d),
      .vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_2_i_qa_d(vec_rsc_0_2_i_qa_d),
      .vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_3_i_qa_d(vec_rsc_0_3_i_qa_d),
      .vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_4_i_qa_d(vec_rsc_0_4_i_qa_d),
      .vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_5_i_qa_d(vec_rsc_0_5_i_qa_d),
      .vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_6_i_qa_d(vec_rsc_0_6_i_qa_d),
      .vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_7_i_qa_d(vec_rsc_0_7_i_qa_d),
      .vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_8_i_qa_d(vec_rsc_0_8_i_qa_d),
      .vec_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_9_i_qa_d(vec_rsc_0_9_i_qa_d),
      .vec_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_10_i_qa_d(vec_rsc_0_10_i_qa_d),
      .vec_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_11_i_qa_d(vec_rsc_0_11_i_qa_d),
      .vec_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_12_i_qa_d(vec_rsc_0_12_i_qa_d),
      .vec_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_13_i_qa_d(vec_rsc_0_13_i_qa_d),
      .vec_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_14_i_qa_d(vec_rsc_0_14_i_qa_d),
      .vec_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_15_i_qa_d(vec_rsc_0_15_i_qa_d),
      .vec_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_0_i_adra_d_pff(vec_rsc_0_0_i_adra_d_iff),
      .vec_rsc_0_0_i_da_d_pff(vec_rsc_0_0_i_da_d_iff),
      .vec_rsc_0_0_i_wea_d_pff(vec_rsc_0_0_i_wea_d_iff),
      .vec_rsc_0_1_i_wea_d_pff(vec_rsc_0_1_i_wea_d_iff),
      .vec_rsc_0_2_i_wea_d_pff(vec_rsc_0_2_i_wea_d_iff),
      .vec_rsc_0_3_i_wea_d_pff(vec_rsc_0_3_i_wea_d_iff),
      .vec_rsc_0_4_i_wea_d_pff(vec_rsc_0_4_i_wea_d_iff),
      .vec_rsc_0_5_i_wea_d_pff(vec_rsc_0_5_i_wea_d_iff),
      .vec_rsc_0_6_i_wea_d_pff(vec_rsc_0_6_i_wea_d_iff),
      .vec_rsc_0_7_i_wea_d_pff(vec_rsc_0_7_i_wea_d_iff),
      .vec_rsc_0_8_i_wea_d_pff(vec_rsc_0_8_i_wea_d_iff),
      .vec_rsc_0_9_i_wea_d_pff(vec_rsc_0_9_i_wea_d_iff),
      .vec_rsc_0_10_i_wea_d_pff(vec_rsc_0_10_i_wea_d_iff),
      .vec_rsc_0_11_i_wea_d_pff(vec_rsc_0_11_i_wea_d_iff),
      .vec_rsc_0_12_i_wea_d_pff(vec_rsc_0_12_i_wea_d_iff),
      .vec_rsc_0_13_i_wea_d_pff(vec_rsc_0_13_i_wea_d_iff),
      .vec_rsc_0_14_i_wea_d_pff(vec_rsc_0_14_i_wea_d_iff),
      .vec_rsc_0_15_i_wea_d_pff(vec_rsc_0_15_i_wea_d_iff)
    );
endmodule



